module fake_ariane_2324_n_9788 (n_83, n_8, n_56, n_60, n_64, n_119, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_52, n_73, n_77, n_15, n_118, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_9788);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_9788;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_9604;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_9297;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_416;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_8438;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_462;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_232;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_2482;
wire n_9665;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_146;
wire n_9241;
wire n_9286;
wire n_4853;
wire n_8744;
wire n_338;
wire n_9592;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_8449;
wire n_9683;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_239;
wire n_3261;
wire n_9358;
wire n_1761;
wire n_9466;
wire n_8953;
wire n_7965;
wire n_7368;
wire n_9787;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_625;
wire n_2322;
wire n_8734;
wire n_1107;
wire n_8720;
wire n_331;
wire n_559;
wire n_2663;
wire n_8097;
wire n_6539;
wire n_5481;
wire n_495;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_7467;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_9714;
wire n_1428;
wire n_1284;
wire n_7526;
wire n_1241;
wire n_4741;
wire n_8664;
wire n_561;
wire n_4143;
wire n_4273;
wire n_507;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_9613;
wire n_9354;
wire n_1519;
wire n_7338;
wire n_5896;
wire n_4567;
wire n_786;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_9516;
wire n_365;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_8939;
wire n_533;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_9202;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_9512;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_579;
wire n_7507;
wire n_844;
wire n_1267;
wire n_8176;
wire n_9677;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_8327;
wire n_8991;
wire n_7438;
wire n_8855;
wire n_4443;
wire n_4119;
wire n_4000;
wire n_9508;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_570;
wire n_5843;
wire n_7874;
wire n_8539;
wire n_8630;
wire n_9308;
wire n_8533;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_9638;
wire n_1121;
wire n_490;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_8435;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_5060;
wire n_9199;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_8958;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5452;
wire n_5391;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_249;
wire n_851;
wire n_123;
wire n_444;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_9265;
wire n_6872;
wire n_6644;
wire n_9143;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_8442;
wire n_1386;
wire n_9304;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_8648;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_9449;
wire n_9149;
wire n_9686;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_203;
wire n_9458;
wire n_4951;
wire n_8585;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_4959;
wire n_9717;
wire n_2745;
wire n_8455;
wire n_2087;
wire n_8444;
wire n_619;
wire n_9128;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_292;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_9715;
wire n_4905;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_1812;
wire n_6659;
wire n_4894;
wire n_9399;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_7583;
wire n_1932;
wire n_6210;
wire n_5680;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_632;
wire n_9094;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_9510;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_382;
wire n_9429;
wire n_489;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_9095;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_9048;
wire n_9003;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_5454;
wire n_307;
wire n_1209;
wire n_4254;
wire n_646;
wire n_8913;
wire n_3438;
wire n_8220;
wire n_404;
wire n_2625;
wire n_9309;
wire n_8355;
wire n_9661;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_299;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_133;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_9063;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_367;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_9110;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_424;
wire n_4857;
wire n_8739;
wire n_8927;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_7963;
wire n_6382;
wire n_8423;
wire n_9028;
wire n_670;
wire n_2677;
wire n_4296;
wire n_379;
wire n_138;
wire n_162;
wire n_9654;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_441;
wire n_7294;
wire n_6192;
wire n_7414;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_207;
wire n_9483;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_194;
wire n_5149;
wire n_9256;
wire n_1163;
wire n_3054;
wire n_5280;
wire n_4970;
wire n_6234;
wire n_4153;
wire n_8992;
wire n_1868;
wire n_5052;
wire n_5137;
wire n_7141;
wire n_3601;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_8510;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_9737;
wire n_8961;
wire n_3323;
wire n_4643;
wire n_9719;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7233;
wire n_7092;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_8402;
wire n_8978;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_9105;
wire n_9699;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_9673;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_1828;
wire n_9240;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_9212;
wire n_5985;
wire n_8595;
wire n_604;
wire n_478;
wire n_9040;
wire n_1349;
wire n_9478;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_9742;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_129;
wire n_126;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_8555;
wire n_9456;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_9146;
wire n_688;
wire n_7176;
wire n_636;
wire n_8565;
wire n_8334;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_442;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_9573;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_887;
wire n_9379;
wire n_9219;
wire n_2125;
wire n_1156;
wire n_5123;
wire n_4974;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_8753;
wire n_1498;
wire n_1188;
wire n_7527;
wire n_9706;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_9206;
wire n_2707;
wire n_8485;
wire n_6482;
wire n_5596;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_9434;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_9082;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_9596;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_9559;
wire n_9709;
wire n_2452;
wire n_8626;
wire n_4182;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_8166;
wire n_9356;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_8602;
wire n_9609;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_5613;
wire n_4662;
wire n_7472;
wire n_9342;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_7989;
wire n_8047;
wire n_744;
wire n_2821;
wire n_3696;
wire n_9233;
wire n_7936;
wire n_215;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_8800;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_9435;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_9557;
wire n_2211;
wire n_8955;
wire n_9551;
wire n_951;
wire n_8039;
wire n_8193;
wire n_9073;
wire n_7546;
wire n_8432;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_6456;
wire n_5108;
wire n_722;
wire n_7407;
wire n_9388;
wire n_3277;
wire n_9721;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_6484;
wire n_5435;
wire n_4429;
wire n_3340;
wire n_7182;
wire n_5053;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_9539;
wire n_8617;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_1243;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_3486;
wire n_6639;
wire n_358;
wire n_608;
wire n_9672;
wire n_9187;
wire n_2457;
wire n_9572;
wire n_2992;
wire n_6124;
wire n_9527;
wire n_317;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_266;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_8192;
wire n_9251;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_8573;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_480;
wire n_7918;
wire n_642;
wire n_9546;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9181;
wire n_9602;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_9635;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_386;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_197;
wire n_2723;
wire n_1476;
wire n_7346;
wire n_6036;
wire n_9405;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_6102;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_9726;
wire n_8804;
wire n_9577;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_9250;
wire n_1330;
wire n_906;
wire n_6204;
wire n_9540;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_9350;
wire n_374;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_9441;
wire n_7600;
wire n_9124;
wire n_2386;
wire n_5826;
wire n_8697;
wire n_9626;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_9408;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_6179;
wire n_5441;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_8406;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_8480;
wire n_9754;
wire n_4419;
wire n_8849;
wire n_5405;
wire n_9750;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_9529;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_9566;
wire n_6442;
wire n_8241;
wire n_140;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_8261;
wire n_6840;
wire n_142;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_8235;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_8294;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_2506;
wire n_8349;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_9443;
wire n_9607;
wire n_7497;
wire n_7315;
wire n_8429;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_9298;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_9052;
wire n_2070;
wire n_426;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_398;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_8117;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_9535;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_400;
wire n_7972;
wire n_8672;
wire n_7505;
wire n_3921;
wire n_282;
wire n_467;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_8934;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_168;
wire n_9555;
wire n_1517;
wire n_2647;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_9030;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_7573;
wire n_6630;
wire n_5759;
wire n_5629;
wire n_2411;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_9590;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_8225;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_9583;
wire n_9763;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6395;
wire n_3497;
wire n_6403;
wire n_4542;
wire n_6578;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_565;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_9617;
wire n_4060;
wire n_1647;
wire n_9341;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_8689;
wire n_3396;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_452;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_8330;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_9349;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_8163;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_8907;
wire n_409;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_9423;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_2669;
wire n_8698;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6541;
wire n_6248;
wire n_9034;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_7927;
wire n_161;
wire n_8928;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_8650;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_9041;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_9011;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_9135;
wire n_6744;
wire n_3645;
wire n_9776;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_132;
wire n_9413;
wire n_9107;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_494;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_9775;
wire n_1805;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_9288;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_164;
wire n_2843;
wire n_3714;
wire n_9305;
wire n_9093;
wire n_184;
wire n_7671;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_8643;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_9425;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_160;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_4496;
wire n_9347;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_8477;
wire n_1775;
wire n_908;
wire n_1036;
wire n_9344;
wire n_7109;
wire n_8028;
wire n_341;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_9530;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_8530;
wire n_9446;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_8500;
wire n_6716;
wire n_8713;
wire n_3565;
wire n_7885;
wire n_8297;
wire n_6905;
wire n_8926;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_9025;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_9713;
wire n_3804;
wire n_4659;
wire n_8293;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_9314;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_9660;
wire n_5763;
wire n_3633;
wire n_857;
wire n_363;
wire n_6061;
wire n_1235;
wire n_9769;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_8726;
wire n_731;
wire n_8977;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_7297;
wire n_784;
wire n_4339;
wire n_5907;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_9410;
wire n_2651;
wire n_753;
wire n_9588;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_309;
wire n_1344;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_9740;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_9061;
wire n_7995;
wire n_8113;
wire n_9579;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_8724;
wire n_7140;
wire n_614;
wire n_4066;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_8253;
wire n_9258;
wire n_9228;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_9598;
wire n_248;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_228;
wire n_6668;
wire n_9311;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_8232;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_8803;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_9608;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_9433;
wire n_658;
wire n_362;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_9537;
wire n_1777;
wire n_9552;
wire n_9421;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_8567;
wire n_8259;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_9473;
wire n_860;
wire n_6525;
wire n_3555;
wire n_9469;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_450;
wire n_8578;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_8336;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_7788;
wire n_5548;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_8600;
wire n_8229;
wire n_415;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_9369;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_9757;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_8761;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_304;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_9729;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_174;
wire n_6379;
wire n_9647;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_8948;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_9275;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_9520;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_9493;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5966;
wire n_4591;
wire n_5569;
wire n_9102;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_9424;
wire n_7160;
wire n_7324;
wire n_9333;
wire n_8205;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_1808;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_8440;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_359;
wire n_9670;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_9200;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_9417;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_9386;
wire n_8897;
wire n_7676;
wire n_8177;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_9207;
wire n_1916;
wire n_6285;
wire n_610;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_8829;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_9728;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_137;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_9465;
wire n_3938;
wire n_8937;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_5250;
wire n_4842;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_9702;
wire n_6607;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_9000;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_9610;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_8503;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_9139;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_8315;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_8197;
wire n_402;
wire n_1979;
wire n_9407;
wire n_6616;
wire n_6719;
wire n_829;
wire n_8019;
wire n_8801;
wire n_4814;
wire n_339;
wire n_6178;
wire n_8707;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_8962;
wire n_8931;
wire n_8248;
wire n_1283;
wire n_7550;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_9357;
wire n_2442;
wire n_9477;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_6443;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_518;
wire n_8196;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_8822;
wire n_3474;
wire n_5738;
wire n_9514;
wire n_2458;
wire n_7971;
wire n_8885;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_8474;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_9501;
wire n_9043;
wire n_8152;
wire n_8269;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_9481;
wire n_3571;
wire n_238;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_9351;
wire n_9766;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_8058;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_612;
wire n_333;
wire n_5107;
wire n_7165;
wire n_512;
wire n_9777;
wire n_4680;
wire n_5067;
wire n_9522;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_9748;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_9005;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_9666;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_461;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_9605;
wire n_2981;
wire n_225;
wire n_1006;
wire n_546;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_3429;
wire n_2969;
wire n_9768;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_8748;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_1872;
wire n_9656;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_9475;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_9724;
wire n_2426;
wire n_652;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_4850;
wire n_9154;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_8740;
wire n_5574;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_460;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_8296;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_9589;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_8850;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_8993;
wire n_9205;
wire n_9418;
wire n_288;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_8831;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_2202;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_8758;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_9020;
wire n_9260;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_9619;
wire n_1079;
wire n_5200;
wire n_9235;
wire n_3393;
wire n_8652;
wire n_9112;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_9133;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_9752;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_8999;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_9353;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_425;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_8499;
wire n_9397;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_9767;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_3796;
wire n_9384;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_155;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_9310;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_172;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_9322;
wire n_7616;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_9377;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_9224;
wire n_3981;
wire n_7271;
wire n_9055;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_345;
wire n_9624;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_9145;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_776;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_130;
wire n_6387;
wire n_466;
wire n_9373;
wire n_4201;
wire n_346;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_552;
wire n_9770;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_9468;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_9517;
wire n_926;
wire n_9544;
wire n_2296;
wire n_7959;
wire n_5735;
wire n_8234;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_8488;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_9774;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_9586;
wire n_3377;
wire n_6722;
wire n_9780;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_2059;
wire n_8184;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_6981;
wire n_7776;
wire n_4870;
wire n_4818;
wire n_8001;
wire n_8695;
wire n_7436;
wire n_8767;
wire n_8571;
wire n_7020;
wire n_8064;
wire n_5935;
wire n_6696;
wire n_8472;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_529;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_5488;
wire n_9099;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_7694;
wire n_3734;
wire n_6787;
wire n_8771;
wire n_5711;
wire n_9245;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_2523;
wire n_1945;
wire n_9168;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_3222;
wire n_325;
wire n_1740;
wire n_4616;
wire n_6011;
wire n_5016;
wire n_9367;
wire n_9330;
wire n_7465;
wire n_5470;
wire n_8917;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_9300;
wire n_3868;
wire n_729;
wire n_8230;
wire n_6222;
wire n_2218;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_390;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_9496;
wire n_8914;
wire n_8821;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_5362;
wire n_8209;
wire n_388;
wire n_8986;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_1055;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_8514;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_8151;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_9329;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_9627;
wire n_3551;
wire n_417;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_9585;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_148;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_6547;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_9606;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_476;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_8841;
wire n_9084;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_7818;
wire n_509;
wire n_7645;
wire n_7482;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_8618;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_9616;
wire n_9708;
wire n_1400;
wire n_7862;
wire n_9130;
wire n_3735;
wire n_8703;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_8061;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_4891;
wire n_8837;
wire n_2629;
wire n_3369;
wire n_8915;
wire n_1257;
wire n_1954;
wire n_8784;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_9086;
wire n_1897;
wire n_8768;
wire n_6999;
wire n_8086;
wire n_8072;
wire n_9014;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_9010;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_9044;
wire n_2912;
wire n_5936;
wire n_8307;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_9694;
wire n_1757;
wire n_8470;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_9633;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_3408;
wire n_2884;
wire n_1293;
wire n_961;
wire n_469;
wire n_9261;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_9345;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_8603;
wire n_9487;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_9271;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_2022;
wire n_6850;
wire n_4343;
wire n_3879;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_949;
wire n_2454;
wire n_9101;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_198;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_8509;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_4173;
wire n_8354;
wire n_5309;
wire n_6047;
wire n_9432;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_422;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_7939;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_8609;
wire n_1143;
wire n_9144;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_9693;
wire n_1153;
wire n_9273;
wire n_271;
wire n_465;
wire n_9196;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_9029;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_256;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_8819;
wire n_914;
wire n_7870;
wire n_689;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_455;
wire n_588;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_9733;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_9075;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_8906;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_9442;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_9630;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_9582;
wire n_1534;
wire n_8268;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_9636;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_6455;
wire n_673;
wire n_5020;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_9412;
wire n_8874;
wire n_8228;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_9525;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_8172;
wire n_4455;
wire n_3241;
wire n_6554;
wire n_3899;
wire n_9575;
wire n_5631;
wire n_3481;
wire n_280;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_9738;
wire n_6020;
wire n_2236;
wire n_9252;
wire n_6185;
wire n_8344;
wire n_692;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_223;
wire n_2150;
wire n_8738;
wire n_8936;
wire n_9739;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_9727;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_6501;
wire n_5608;
wire n_2204;
wire n_9148;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_9323;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_8088;
wire n_5702;
wire n_9545;
wire n_8930;
wire n_9155;
wire n_8662;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_9046;
wire n_9430;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_9625;
wire n_8783;
wire n_8663;
wire n_1221;
wire n_4217;
wire n_5182;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_9447;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_8364;
wire n_9485;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_8490;
wire n_9129;
wire n_229;
wire n_8981;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_8785;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_9047;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_8982;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_6993;
wire n_9745;
wire n_508;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_8522;
wire n_1361;
wire n_8381;
wire n_9320;
wire n_8835;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_6558;
wire n_1411;
wire n_1359;
wire n_5687;
wire n_6755;
wire n_9108;
wire n_9457;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_9567;
wire n_294;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_8736;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_8918;
wire n_2402;
wire n_1458;
wire n_679;
wire n_220;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_387;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_8838;
wire n_8908;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_9161;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_8607;
wire n_607;
wire n_8213;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_8436;
wire n_7282;
wire n_372;
wire n_8551;
wire n_2770;
wire n_4550;
wire n_9238;
wire n_4347;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_9248;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_311;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_269;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_9071;
wire n_446;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_9519;
wire n_1629;
wire n_9027;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_3002;
wire n_8984;
wire n_9786;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_8613;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_9404;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_8387;
wire n_9352;
wire n_8105;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_9681;
wire n_8353;
wire n_505;
wire n_9051;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3775;
wire n_3148;
wire n_5682;
wire n_684;
wire n_5461;
wire n_9098;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_6164;
wire n_8711;
wire n_3616;
wire n_4753;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_175;
wire n_3637;
wire n_8534;
wire n_1017;
wire n_8655;
wire n_9210;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_8302;
wire n_4258;
wire n_5756;
wire n_310;
wire n_8496;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_662;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_9756;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_572;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_4767;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_948;
wire n_448;
wire n_6528;
wire n_9700;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_8335;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_9363;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_9532;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_9307;
wire n_3910;
wire n_3947;
wire n_492;
wire n_252;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_3228;
wire n_8834;
wire n_8286;
wire n_8417;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_8964;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_2205;
wire n_2183;
wire n_389;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_9406;
wire n_4520;
wire n_895;
wire n_8639;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_9160;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_7712;
wire n_4444;
wire n_6885;
wire n_7681;
wire n_8566;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_8727;
wire n_5039;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_265;
wire n_1583;
wire n_8599;
wire n_4612;
wire n_5997;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6602;
wire n_6530;
wire n_7915;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_6135;
wire n_246;
wire n_8839;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_8365;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_289;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_9705;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_8367;
wire n_9113;
wire n_3484;
wire n_6001;
wire n_411;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_2095;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_5823;
wire n_8658;
wire n_8898;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_8905;
wire n_9222;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_9394;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_9723;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_8946;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_245;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_9069;
wire n_525;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_3742;
wire n_7601;
wire n_8998;
wire n_4965;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_189;
wire n_8157;
wire n_2006;
wire n_9284;
wire n_4953;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_9556;
wire n_5294;
wire n_8161;
wire n_5570;
wire n_6411;
wire n_9337;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_9211;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_9243;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_9773;
wire n_4674;
wire n_8812;
wire n_568;
wire n_8682;
wire n_8290;
wire n_4796;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_377;
wire n_2750;
wire n_8890;
wire n_2547;
wire n_8747;
wire n_7617;
wire n_279;
wire n_945;
wire n_4575;
wire n_9784;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_9192;
wire n_6008;
wire n_500;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_9134;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_9765;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_7876;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_143;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_6517;
wire n_5665;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_9564;
wire n_9127;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_9306;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_222;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_9332;
wire n_3756;
wire n_8043;
wire n_8223;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_4608;
wire n_9294;
wire n_6691;
wire n_432;
wire n_293;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_9132;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_206;
wire n_2332;
wire n_9547;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6536;
wire n_6029;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_3049;
wire n_8434;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_9762;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_9183;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_6877;
wire n_7308;
wire n_5639;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_209;
wire n_5503;
wire n_5718;
wire n_1461;
wire n_7208;
wire n_5240;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_503;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_9001;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_380;
wire n_3119;
wire n_6671;
wire n_9335;
wire n_4740;
wire n_1108;
wire n_9488;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_6444;
wire n_6637;
wire n_5544;
wire n_9725;
wire n_8842;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_9526;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_577;
wire n_5610;
wire n_407;
wire n_8576;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_8799;
wire n_762;
wire n_1468;
wire n_1253;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_9716;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_513;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_8227;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_436;
wire n_5770;
wire n_7483;
wire n_8756;
wire n_5710;
wire n_324;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_274;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_8604;
wire n_8809;
wire n_8976;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_8940;
wire n_5008;
wire n_1312;
wire n_9077;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_8844;
wire n_6148;
wire n_8995;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_8693;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_712;
wire n_8769;
wire n_9463;
wire n_909;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_8990;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_8512;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_9710;
wire n_2507;
wire n_1633;
wire n_9087;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_7845;
wire n_2328;
wire n_5285;
wire n_347;
wire n_2434;
wire n_183;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_9782;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_9197;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_9140;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_370;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_286;
wire n_9364;
wire n_9452;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_9362;
wire n_9398;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_9203;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_9712;
wire n_9536;
wire n_8450;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_9460;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_8324;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_9772;
wire n_1496;
wire n_2812;
wire n_9057;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_9068;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_8623;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_9348;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_8651;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_9632;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_9500;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_9747;
wire n_2350;
wire n_9470;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_9591;
wire n_9049;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_8413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_158;
wire n_3882;
wire n_9471;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_405;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_7501;
wire n_320;
wire n_9409;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_481;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_547;
wire n_439;
wire n_677;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_703;
wire n_8400;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_326;
wire n_227;
wire n_3773;
wire n_3494;
wire n_9482;
wire n_1278;
wire n_9033;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_545;
wire n_9247;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_536;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_9299;
wire n_3139;
wire n_8889;
wire n_427;
wire n_5681;
wire n_3801;
wire n_9244;
wire n_9785;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_9195;
wire n_8322;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_3653;
wire n_3823;
wire n_9280;
wire n_3403;
wire n_7621;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_314;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_7985;
wire n_9687;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_233;
wire n_8954;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_321;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_1586;
wire n_8728;
wire n_9580;
wire n_9569;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_9680;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_8407;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_9227;
wire n_5657;
wire n_8475;
wire n_297;
wire n_2379;
wire n_3579;
wire n_9072;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_178;
wire n_551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_8511;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_9584;
wire n_9287;
wire n_534;
wire n_2508;
wire n_3186;
wire n_9459;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_9490;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_560;
wire n_8558;
wire n_890;
wire n_9655;
wire n_3626;
wire n_451;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_9147;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_9678;
wire n_2119;
wire n_8641;
wire n_9658;
wire n_2493;
wire n_9560;
wire n_9578;
wire n_5080;
wire n_535;
wire n_9396;
wire n_4565;
wire n_7032;
wire n_9303;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_9553;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_8046;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_8292;
wire n_5567;
wire n_9138;
wire n_5406;
wire n_8647;
wire n_6362;
wire n_9213;
wire n_4328;
wire n_8543;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_9374;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_5867;
wire n_456;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_9179;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_342;
wire n_5602;
wire n_2035;
wire n_7196;
wire n_4928;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8174;
wire n_8187;
wire n_8929;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_8846;
wire n_5817;
wire n_9277;
wire n_4160;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_1668;
wire n_9744;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_9504;
wire n_5417;
wire n_4545;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_9285;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_9190;
wire n_8586;
wire n_8524;
wire n_618;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_9639;
wire n_4385;
wire n_7779;
wire n_9664;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_9109;
wire n_211;
wire n_1804;
wire n_408;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_9741;
wire n_2272;
wire n_5989;
wire n_4766;
wire n_5571;
wire n_592;
wire n_4558;
wire n_1318;
wire n_8764;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_8502;
wire n_4319;
wire n_9360;
wire n_6585;
wire n_7786;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_4358;
wire n_9122;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_2857;
wire n_8564;
wire n_8343;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_9013;
wire n_5431;
wire n_9427;
wire n_8379;
wire n_643;
wire n_8034;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_9126;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_8441;
wire n_9474;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_9538;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_8569;
wire n_9574;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_8592;
wire n_8865;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_8362;
wire n_3336;
wire n_8632;
wire n_7739;
wire n_396;
wire n_7945;
wire n_9372;
wire n_9045;
wire n_8361;
wire n_9657;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_725;
wire n_8611;
wire n_9326;
wire n_8410;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_9476;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_272;
wire n_8492;
wire n_9301;
wire n_7213;
wire n_5313;
wire n_4301;
wire n_2133;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_9382;
wire n_8095;
wire n_7369;
wire n_1472;
wire n_9325;
wire n_1050;
wire n_9643;
wire n_7548;
wire n_2578;
wire n_152;
wire n_1201;
wire n_8735;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_335;
wire n_2665;
wire n_4879;
wire n_344;
wire n_8794;
wire n_5044;
wire n_210;
wire n_1090;
wire n_4536;
wire n_3755;
wire n_9274;
wire n_8549;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_224;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_8593;
wire n_276;
wire n_9649;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_8195;
wire n_8009;
wire n_8588;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_9346;
wire n_6673;
wire n_9696;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_9383;
wire n_9498;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_305;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_361;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_181;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_1362;
wire n_9509;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_7463;
wire n_9621;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_8627;
wire n_1210;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_9563;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_8858;
wire n_414;
wire n_571;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_8916;
wire n_613;
wire n_1022;
wire n_5465;
wire n_171;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_820;
wire n_8260;
wire n_254;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_8688;
wire n_7969;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_9550;
wire n_532;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_621;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_6879;
wire n_9562;
wire n_9612;
wire n_493;
wire n_1311;
wire n_3106;
wire n_7190;
wire n_6208;
wire n_9698;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_9528;
wire n_4620;
wire n_5397;
wire n_6457;
wire n_6255;
wire n_9272;
wire n_9645;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_2305;
wire n_8737;
wire n_9731;
wire n_5996;
wire n_880;
wire n_5566;
wire n_9697;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7237;
wire n_7082;
wire n_8988;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_9642;
wire n_530;
wire n_8723;
wire n_9050;
wire n_4406;
wire n_2180;
wire n_4271;
wire n_7042;
wire n_8419;
wire n_2809;
wire n_5652;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_9531;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_8826;
wire n_3178;
wire n_268;
wire n_7023;
wire n_2251;
wire n_9732;
wire n_5758;
wire n_5842;
wire n_9685;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_8959;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_191;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_8712;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_9378;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_3576;
wire n_9389;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_332;
wire n_8910;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_541;
wire n_499;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_8892;
wire n_9637;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_9491;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_7180;
wire n_5952;
wire n_2086;
wire n_1926;
wire n_8972;
wire n_8494;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_443;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_8941;
wire n_8891;
wire n_406;
wire n_3897;
wire n_7103;
wire n_139;
wire n_6605;
wire n_1735;
wire n_391;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_6832;
wire n_5980;
wire n_8683;
wire n_956;
wire n_9391;
wire n_765;
wire n_4092;
wire n_122;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_2758;
wire n_385;
wire n_6544;
wire n_8810;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_399;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_2471;
wire n_9695;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_9255;
wire n_8882;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_3598;
wire n_7706;
wire n_7813;
wire n_4917;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_153;
wire n_648;
wire n_6836;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_835;
wire n_9136;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_9436;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_9042;
wire n_839;
wire n_1754;
wire n_7236;
wire n_9239;
wire n_4833;
wire n_3394;
wire n_9570;
wire n_6405;
wire n_8345;
wire n_9644;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_9343;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_9131;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_8636;
wire n_9006;
wire n_9221;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_539;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_459;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_9523;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_6175;
wire n_6445;
wire n_8563;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_9411;
wire n_1982;
wire n_7983;
wire n_641;
wire n_5311;
wire n_8765;
wire n_910;
wire n_290;
wire n_5164;
wire n_4964;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_217;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_8601;
wire n_1043;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_8333;
wire n_9097;
wire n_9571;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_196;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_9511;
wire n_3196;
wire n_231;
wire n_8708;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_8659;
wire n_6732;
wire n_8759;
wire n_2548;
wire n_3488;
wire n_9622;
wire n_2381;
wire n_9761;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_3779;
wire n_599;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_8790;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_583;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_378;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_9640;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_9115;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_9534;
wire n_472;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_208;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_7554;
wire n_275;
wire n_4852;
wire n_3202;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_147;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_9594;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_8347;
wire n_131;
wire n_2255;
wire n_5554;
wire n_9503;
wire n_1252;
wire n_3045;
wire n_250;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_8093;
wire n_8899;
wire n_9385;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_8481;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_9182;
wire n_1582;
wire n_8182;
wire n_9426;
wire n_9293;
wire n_1981;
wire n_2824;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_5900;
wire n_8629;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_9400;
wire n_4013;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_691;
wire n_6819;
wire n_6122;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5851;
wire n_7516;
wire n_5432;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_187;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_8750;
wire n_8183;
wire n_4997;
wire n_5065;
wire n_9104;
wire n_6806;
wire n_924;
wire n_7991;
wire n_781;
wire n_8637;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_9542;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_9302;
wire n_1706;
wire n_2461;
wire n_8258;
wire n_3719;
wire n_7154;
wire n_524;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_8416;
wire n_8390;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_5173;
wire n_4683;
wire n_2873;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_7175;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_6316;
wire n_8619;
wire n_419;
wire n_7068;
wire n_2908;
wire n_8594;
wire n_270;
wire n_4106;
wire n_9541;
wire n_285;
wire n_2156;
wire n_1184;
wire n_202;
wire n_8162;
wire n_9735;
wire n_754;
wire n_9576;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_8318;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_3283;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_9039;
wire n_7384;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_6561;
wire n_5678;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_8389;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_200;
wire n_2539;
wire n_8620;
wire n_5555;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_8202;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_8755;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3230;
wire n_3793;
wire n_859;
wire n_8199;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_8004;
wire n_8383;
wire n_3607;
wire n_1637;
wire n_9688;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_9023;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_438;
wire n_8680;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_440;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_7446;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6620;
wire n_6245;
wire n_6030;
wire n_1544;
wire n_6791;
wire n_4360;
wire n_4540;
wire n_9220;
wire n_6821;
wire n_9317;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_1354;
wire n_8665;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_9561;
wire n_491;
wire n_9444;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_9184;
wire n_7559;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_9505;
wire n_9193;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_4495;
wire n_3958;
wire n_4737;
wire n_1838;
wire n_9218;
wire n_9755;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_8782;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_9162;
wire n_9506;
wire n_135;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_1691;
wire n_8250;
wire n_7264;
wire n_7842;
wire n_2549;
wire n_2499;
wire n_6648;
wire n_9415;
wire n_7492;
wire n_804;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_9015;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_9214;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_8922;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_8498;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_3937;
wire n_4763;
wire n_9339;
wire n_1418;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_8267;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_615;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_517;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_824;
wire n_159;
wire n_8319;
wire n_7997;
wire n_5659;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_144;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_8581;
wire n_4267;
wire n_8214;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_3021;
wire n_8989;
wire n_7746;
wire n_477;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_9650;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_7894;
wire n_9282;
wire n_1147;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_8289;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_356;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_8863;
wire n_9371;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_9237;
wire n_2311;
wire n_6857;
wire n_8705;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_205;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_7665;
wire n_4836;
wire n_3889;
wire n_7677;
wire n_5262;
wire n_5522;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_261;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_9480;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_9597;
wire n_348;
wire n_9173;
wire n_2312;
wire n_7203;
wire n_8947;
wire n_9641;
wire n_7797;
wire n_1826;
wire n_9267;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_8786;
wire n_9414;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_9419;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_8276;
wire n_7284;
wire n_3615;
wire n_5516;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_145;
wire n_2146;
wire n_5583;
wire n_4274;
wire n_3276;
wire n_7064;
wire n_8532;
wire n_9533;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_9618;
wire n_5698;
wire n_5731;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_8433;
wire n_9065;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_9674;
wire n_6617;
wire n_553;
wire n_7725;
wire n_814;
wire n_578;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_8467;
wire n_647;
wire n_2027;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_600;
wire n_3118;
wire n_9157;
wire n_5560;
wire n_9170;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_6777;
wire n_502;
wire n_5455;
wire n_8640;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_247;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_8431;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_9416;
wire n_3974;
wire n_9368;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_8089;
wire n_5022;
wire n_9208;
wire n_6370;
wire n_9223;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_9781;
wire n_3009;
wire n_8633;
wire n_777;
wire n_7095;
wire n_7390;
wire n_9392;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_920;
wire n_8541;
wire n_8762;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_9338;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_9492;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_9328;
wire n_6465;
wire n_221;
wire n_8188;
wire n_5673;
wire n_861;
wire n_8615;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_8923;
wire n_281;
wire n_3326;
wire n_8624;
wire n_262;
wire n_8222;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9513;
wire n_3224;
wire n_9393;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_527;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_343;
wire n_1222;
wire n_7139;
wire n_8935;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_8155;
wire n_9334;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_9684;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_9254;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_9083;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_657;
wire n_7060;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_8873;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_7444;
wire n_6750;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_430;
wire n_3953;
wire n_7502;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_9554;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_9116;
wire n_9315;
wire n_8825;
wire n_852;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_9215;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_8395;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_8164;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_8877;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_134;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_1480;
wire n_3670;
wire n_8366;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_157;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_624;
wire n_5577;
wire n_876;
wire n_9100;
wire n_5872;
wire n_7883;
wire n_6692;
wire n_9707;
wire n_5017;
wire n_8854;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_8256;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_8621;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_8577;
wire n_9019;
wire n_2725;
wire n_2667;
wire n_9361;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_421;
wire n_3702;
wire n_5930;
wire n_8952;
wire n_1984;
wire n_3453;
wire n_9438;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_7458;
wire n_4427;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_3543;
wire n_586;
wire n_1324;
wire n_2945;
wire n_8421;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_9327;
wire n_9313;
wire n_605;
wire n_2936;
wire n_3609;
wire n_6334;
wire n_4330;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_8911;
wire n_5537;
wire n_9518;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_8971;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_9291;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_9722;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_151;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_8949;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_9454;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_8983;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_8942;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_173;
wire n_2796;
wire n_858;
wire n_5393;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_2136;
wire n_433;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_253;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_128;
wire n_7916;
wire n_3055;
wire n_8194;
wire n_420;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_9453;
wire n_748;
wire n_7903;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_9331;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4769;
wire n_4139;
wire n_6130;
wire n_330;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_8285;
wire n_7145;
wire n_8521;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_9178;
wire n_7803;
wire n_9689;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_9355;
wire n_9489;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_576;
wire n_8732;
wire n_511;
wire n_7622;
wire n_9359;
wire n_429;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_8420;
wire n_141;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_9568;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_312;
wire n_728;
wire n_4409;
wire n_4191;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_8746;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_9401;
wire n_8857;
wire n_543;
wire n_6986;
wire n_9495;
wire n_3456;
wire n_4532;
wire n_236;
wire n_601;
wire n_7564;
wire n_628;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_9234;
wire n_7960;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_8281;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_593;
wire n_8766;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_609;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_9340;
wire n_9380;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_519;
wire n_8314;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_9064;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_9746;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_9066;
wire n_763;
wire n_6301;
wire n_2174;
wire n_540;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_7686;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_395;
wire n_6737;
wire n_1587;
wire n_213;
wire n_2340;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_9455;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_8505;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_8606;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_9440;
wire n_4759;
wire n_9059;
wire n_5869;
wire n_6753;
wire n_2114;
wire n_5914;
wire n_9690;
wire n_3329;
wire n_3833;
wire n_2927;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_9002;
wire n_3402;
wire n_9620;
wire n_1621;
wire n_6448;
wire n_9229;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_9464;
wire n_434;
wire n_4687;
wire n_7077;
wire n_394;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_4720;
wire n_2889;
wire n_6268;
wire n_6043;
wire n_9497;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_243;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_8408;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_7214;
wire n_8806;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_9587;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_121;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_8377;
wire n_3989;
wire n_7652;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_558;
wire n_5325;
wire n_4231;
wire n_8960;
wire n_9008;
wire n_8957;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_9549;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_9652;
wire n_7975;
wire n_8451;
wire n_6089;
wire n_591;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_8527;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_9089;
wire n_4578;
wire n_318;
wire n_8840;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_3644;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_9080;
wire n_1922;
wire n_9296;
wire n_940;
wire n_1537;
wire n_4877;
wire n_9312;
wire n_2065;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_8287;
wire n_1904;
wire n_8111;
wire n_8341;
wire n_8830;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_9324;
wire n_9631;
wire n_8308;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_8965;
wire n_9736;
wire n_2258;
wire n_7041;
wire n_9365;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_9600;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_6672;
wire n_5343;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_9402;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_6242;
wire n_5947;
wire n_336;
wire n_6601;
wire n_8570;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_8579;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_9711;
wire n_9759;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_6606;
wire n_4497;
wire n_2583;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_8320;
wire n_8635;
wire n_9703;
wire n_4472;
wire n_9118;
wire n_2699;
wire n_9321;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_2973;
wire n_9428;
wire n_8612;
wire n_8778;
wire n_5893;
wire n_9292;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_9018;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_369;
wire n_240;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_9565;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_7337;
wire n_5726;
wire n_4566;
wire n_3933;
wire n_7439;
wire n_4310;
wire n_4371;
wire n_188;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_8458;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_9603;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_8306;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_8342;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_9012;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_383;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_630;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_8445;
wire n_1781;
wire n_9720;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8464;
wire n_8363;
wire n_8921;
wire n_235;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_9646;
wire n_7480;
wire n_8843;
wire n_371;
wire n_5185;
wire n_8405;
wire n_2964;
wire n_8376;
wire n_308;
wire n_5032;
wire n_6990;
wire n_865;
wire n_7071;
wire n_3312;
wire n_5034;
wire n_1041;
wire n_2451;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_8752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8894;
wire n_7380;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_9671;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_5115;
wire n_7376;
wire n_8411;
wire n_902;
wire n_8817;
wire n_8461;
wire n_1723;
wire n_3918;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_6409;
wire n_8391;
wire n_4095;
wire n_8507;
wire n_1310;
wire n_5927;
wire n_8691;
wire n_9188;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_574;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_9614;
wire n_8967;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_9628;
wire n_1896;
wire n_9231;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_8084;
wire n_8856;
wire n_2485;
wire n_6679;
wire n_8631;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_9730;
wire n_5507;
wire n_195;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_8338;
wire n_1631;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_156;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_1794;
wire n_9462;
wire n_5696;
wire n_7998;
wire n_8666;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_496;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_9515;
wire n_9502;
wire n_263;
wire n_5235;
wire n_4516;
wire n_360;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_165;
wire n_9316;
wire n_3217;
wire n_8938;
wire n_6081;
wire n_1249;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_8523;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_177;
wire n_364;
wire n_258;
wire n_7582;
wire n_5521;
wire n_431;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_8924;
wire n_2965;
wire n_7555;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_9494;
wire n_5018;
wire n_4134;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

BUFx10_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_50),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_19),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_47),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_27),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_43),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_27),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_60),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_24),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_70),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_23),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_48),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_21),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_59),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_32),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_88),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_31),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_55),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_53),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_90),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_66),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_64),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_2),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_11),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_71),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_42),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_29),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_45),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_14),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_57),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_51),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_82),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_86),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_25),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_36),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_13),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_97),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_78),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_18),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_7),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_17),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_26),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_61),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_52),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_17),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_15),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_5),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_76),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_24),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_69),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_72),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_141),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_178),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_195),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_129),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_126),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_149),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_121),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_143),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_169),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_148),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_126),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_140),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_142),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_148),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_265),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_264),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_256),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_272),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_223),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_271),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_242),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_274),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_271),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_274),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_252),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_266),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_276),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_187),
.B1(n_207),
.B2(n_155),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_284),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_291),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_285),
.A2(n_155),
.B1(n_207),
.B2(n_187),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_297),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_296),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_308),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_277),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_280),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_254),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_266),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_267),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_206),
.B1(n_181),
.B2(n_172),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_298),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_282),
.A2(n_198),
.B1(n_163),
.B2(n_145),
.Y(n_360)
);

BUFx8_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_254),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_282),
.B(n_267),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_311),
.B(n_257),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_303),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_296),
.B(n_146),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_292),
.B(n_269),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_283),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_287),
.B(n_269),
.Y(n_373)
);

BUFx8_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_276),
.A2(n_135),
.B1(n_228),
.B2(n_229),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_278),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_283),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_283),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_278),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_275),
.B(n_128),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_275),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_283),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_287),
.B(n_240),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_289),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_276),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_283),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_276),
.A2(n_135),
.B1(n_228),
.B2(n_229),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_288),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_278),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_287),
.B(n_257),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_276),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_287),
.B(n_124),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_289),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_276),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_292),
.B(n_240),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_278),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_288),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_R g405 ( 
.A(n_289),
.B(n_241),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_275),
.B(n_130),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_288),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_289),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_288),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_288),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_278),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_283),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_283),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_287),
.B(n_241),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_283),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_278),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_280),
.B(n_127),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_287),
.B(n_133),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_276),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_278),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_278),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_278),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_283),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_287),
.B(n_244),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_283),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_283),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_287),
.B(n_166),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_292),
.B(n_159),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_276),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_289),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_287),
.B(n_244),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_289),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_362),
.B(n_191),
.Y(n_437)
);

AND3x2_ASAP7_75t_L g438 ( 
.A(n_318),
.B(n_245),
.C(n_164),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_348),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_405),
.A2(n_127),
.B1(n_136),
.B2(n_227),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_314),
.B(n_245),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_323),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_349),
.B(n_136),
.Y(n_447)
);

CKINVDCx6p67_ASAP7_75t_R g448 ( 
.A(n_328),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_345),
.B(n_173),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_349),
.B(n_227),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_343),
.B(n_189),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_328),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_368),
.B(n_230),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_370),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_322),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_341),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_317),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_319),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_369),
.B(n_234),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_351),
.B(n_171),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_321),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_380),
.B(n_406),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_338),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_325),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_355),
.B(n_171),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_326),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_332),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_362),
.B(n_230),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_380),
.B(n_406),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_368),
.B(n_231),
.Y(n_475)
);

INVx3_ASAP7_75t_SL g476 ( 
.A(n_331),
.Y(n_476)
);

AND3x2_ASAP7_75t_L g477 ( 
.A(n_318),
.B(n_165),
.C(n_156),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_316),
.B(n_231),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_335),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_338),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_364),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_363),
.B(n_192),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_367),
.B(n_232),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_369),
.B(n_234),
.Y(n_489)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_423),
.A2(n_186),
.B(n_131),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_334),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_316),
.B(n_232),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_337),
.Y(n_495)
);

NOR3xp33_ASAP7_75t_L g496 ( 
.A(n_375),
.B(n_214),
.C(n_201),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_342),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_315),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_363),
.B(n_134),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_346),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_382),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_347),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_381),
.Y(n_504)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_396),
.A2(n_200),
.B(n_224),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_376),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_363),
.B(n_147),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_402),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_373),
.B(n_193),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_373),
.B(n_212),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_379),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_315),
.Y(n_512)
);

INVx8_ASAP7_75t_L g513 ( 
.A(n_363),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_417),
.B(n_151),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_403),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_417),
.B(n_152),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_336),
.B(n_185),
.C(n_211),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_330),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_385),
.B(n_213),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_330),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_421),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_315),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_390),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_315),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_385),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_324),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_327),
.B(n_222),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_400),
.B(n_408),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_324),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_424),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_432),
.B(n_183),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_324),
.Y(n_542)
);

INVxp33_ASAP7_75t_SL g543 ( 
.A(n_430),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

BUFx6f_ASAP7_75t_SL g545 ( 
.A(n_382),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_324),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_431),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_383),
.B(n_431),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_352),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_352),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_358),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_352),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_365),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_352),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_383),
.B(n_171),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_366),
.B(n_399),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_320),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_353),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_353),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_353),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_405),
.B(n_225),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_353),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_356),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_418),
.B(n_205),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_350),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_428),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_356),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_356),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_356),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_386),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_386),
.Y(n_572)
);

NOR2x1p5_ASAP7_75t_L g573 ( 
.A(n_361),
.B(n_153),
.Y(n_573)
);

NOR2x1p5_ASAP7_75t_L g574 ( 
.A(n_361),
.B(n_176),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_386),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_387),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_329),
.A2(n_220),
.B1(n_176),
.B2(n_146),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_357),
.B(n_121),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_387),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_387),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_387),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_360),
.B(n_121),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_394),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_394),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_394),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_398),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_398),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_398),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_327),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_398),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_404),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_404),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_404),
.B(n_122),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_404),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_407),
.B(n_179),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_407),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_R g599 ( 
.A(n_374),
.B(n_139),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_374),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_339),
.B(n_180),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_336),
.B(n_203),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_407),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_407),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_409),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_409),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_409),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_410),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_410),
.B(n_143),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_410),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_391),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_410),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_393),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_339),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_391),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_397),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_397),
.A2(n_175),
.B1(n_238),
.B2(n_237),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_401),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_333),
.B(n_143),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_401),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_419),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_419),
.B(n_132),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_429),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_429),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_345),
.B(n_132),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_377),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_354),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_345),
.B(n_132),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_354),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_377),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_377),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_377),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_354),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_349),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_377),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_377),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_377),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_377),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_359),
.B(n_143),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_377),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_377),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_354),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_348),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_348),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_377),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_349),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_377),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_362),
.B(n_123),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_377),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_362),
.B(n_138),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_349),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_369),
.B(n_2),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_362),
.B(n_144),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_405),
.B(n_184),
.C(n_226),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_345),
.B(n_203),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_377),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_368),
.B(n_203),
.Y(n_657)
);

NAND3x1_ASAP7_75t_L g658 ( 
.A(n_329),
.B(n_3),
.C(n_4),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_405),
.A2(n_199),
.B1(n_162),
.B2(n_161),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_348),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_359),
.B(n_182),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_354),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_345),
.B(n_204),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_377),
.A2(n_255),
.B(n_218),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_354),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_377),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_359),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_354),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_359),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_359),
.Y(n_670)
);

BUFx16f_ASAP7_75t_R g671 ( 
.A(n_374),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_359),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_359),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_349),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_345),
.B(n_202),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_362),
.B(n_170),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_354),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_345),
.B(n_210),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_377),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_369),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_377),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_354),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_362),
.B(n_168),
.Y(n_683)
);

INVxp33_ASAP7_75t_SL g684 ( 
.A(n_348),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_349),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_369),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_377),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_359),
.B(n_167),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_359),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_354),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_377),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_377),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_349),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_354),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_354),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_345),
.B(n_150),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_348),
.B(n_174),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_369),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_362),
.B(n_188),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_377),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_377),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_362),
.B(n_160),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_354),
.Y(n_703)
);

BUFx6f_ASAP7_75t_SL g704 ( 
.A(n_328),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_354),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_362),
.B(n_197),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_354),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_369),
.B(n_3),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_359),
.B(n_196),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_314),
.B(n_8),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_377),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_377),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_327),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_354),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_377),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_359),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_369),
.B(n_11),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_323),
.Y(n_718)
);

AND2x6_ASAP7_75t_L g719 ( 
.A(n_670),
.B(n_255),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_448),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_657),
.A2(n_194),
.B1(n_158),
.B2(n_157),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_557),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_476),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_495),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_470),
.B(n_154),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_495),
.Y(n_726)
);

BUFx4f_ASAP7_75t_L g727 ( 
.A(n_448),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_433),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_513),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_531),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_621),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_634),
.B(n_12),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_531),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_433),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_557),
.B(n_255),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_12),
.Y(n_737)
);

AND2x6_ASAP7_75t_L g738 ( 
.A(n_670),
.B(n_255),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_548),
.B(n_15),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_470),
.B(n_16),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_497),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_566),
.B(n_465),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_543),
.B(n_657),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_543),
.B(n_16),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_497),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_646),
.B(n_651),
.Y(n_746)
);

NAND3x1_ASAP7_75t_L g747 ( 
.A(n_613),
.B(n_19),
.C(n_20),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_500),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_500),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_513),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_718),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_465),
.B(n_21),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_600),
.B(n_22),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_680),
.B(n_526),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_670),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_503),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_464),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_646),
.B(n_35),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_452),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_670),
.B(n_38),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_503),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_513),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_511),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_667),
.B(n_41),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_511),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_515),
.Y(n_767)
);

AND2x2_ASAP7_75t_SL g768 ( 
.A(n_579),
.B(n_46),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_626),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_667),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_667),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_515),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_548),
.B(n_49),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_680),
.B(n_62),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_516),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_474),
.B(n_65),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_513),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_522),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_465),
.B(n_75),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_556),
.B(n_79),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_525),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_718),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_482),
.B(n_85),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_516),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_518),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_518),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_453),
.B(n_100),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_453),
.B(n_105),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_651),
.B(n_109),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_630),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_674),
.B(n_685),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_667),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_504),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_527),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_630),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_533),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_475),
.B(n_437),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_527),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_631),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_480),
.B(n_486),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_689),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_528),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_475),
.B(n_686),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_533),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_528),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_452),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_458),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_480),
.B(n_486),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_545),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_460),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_616),
.B(n_618),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_545),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_545),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_631),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_462),
.B(n_469),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_689),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_616),
.B(n_618),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_632),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_480),
.B(n_486),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_632),
.B(n_635),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_698),
.B(n_482),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_501),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_689),
.B(n_716),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_463),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_466),
.Y(n_825)
);

AND2x6_ASAP7_75t_L g826 ( 
.A(n_689),
.B(n_716),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_476),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_462),
.B(n_469),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_471),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_704),
.Y(n_830)
);

AND2x6_ASAP7_75t_L g831 ( 
.A(n_716),
.B(n_443),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_716),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_635),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_636),
.B(n_637),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_611),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_439),
.B(n_684),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_636),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_439),
.B(n_684),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_624),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_637),
.B(n_638),
.Y(n_840)
);

AND2x6_ASAP7_75t_L g841 ( 
.A(n_443),
.B(n_669),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_638),
.B(n_640),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_640),
.B(n_641),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_704),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_579),
.B(n_583),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_623),
.B(n_624),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_443),
.B(n_669),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_492),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_674),
.B(n_685),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_693),
.B(n_451),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_619),
.A2(n_561),
.B1(n_540),
.B2(n_613),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_600),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_611),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_619),
.A2(n_561),
.B1(n_540),
.B2(n_613),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_501),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_L g856 ( 
.A(n_615),
.B(n_614),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_693),
.B(n_447),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_704),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_502),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_641),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_506),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_621),
.Y(n_862)
);

XNOR2xp5_ASAP7_75t_L g863 ( 
.A(n_536),
.B(n_591),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_590),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_447),
.B(n_450),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_534),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_599),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_450),
.B(n_625),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_514),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_538),
.B(n_544),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_520),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_446),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_524),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_643),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_713),
.B(n_454),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_621),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_628),
.B(n_655),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_586),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_529),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_669),
.B(n_672),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_547),
.B(n_454),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_508),
.B(n_710),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_645),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_647),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_436),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_498),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_541),
.B(n_583),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_648),
.B(n_650),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_672),
.B(n_673),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_555),
.B(n_508),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_649),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_455),
.Y(n_892)
);

BUFx10_ASAP7_75t_L g893 ( 
.A(n_449),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_649),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_710),
.B(n_442),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_541),
.B(n_473),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_656),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_498),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_656),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_455),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_653),
.B(n_676),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_683),
.B(n_699),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_446),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_702),
.B(n_706),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_659),
.B(n_446),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_498),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_666),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_456),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_590),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_620),
.B(n_461),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_666),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_456),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_457),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_643),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_457),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_479),
.B(n_654),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_459),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_459),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_672),
.B(n_673),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_679),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_681),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_479),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_442),
.B(n_602),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_467),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_602),
.B(n_555),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_479),
.B(n_551),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_467),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_622),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_468),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_614),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_643),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_567),
.B(n_573),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_551),
.B(n_484),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_468),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_687),
.A2(n_701),
.B1(n_715),
.B2(n_712),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_622),
.B(n_440),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_687),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_461),
.B(n_489),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_590),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_472),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_472),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_691),
.Y(n_942)
);

BUFx6f_ASAP7_75t_SL g943 ( 
.A(n_644),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_644),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_481),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_586),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_663),
.A2(n_696),
.B1(n_675),
.B2(n_678),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_481),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_691),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_R g950 ( 
.A(n_614),
.B(n_478),
.Y(n_950)
);

AND2x6_ASAP7_75t_L g951 ( 
.A(n_673),
.B(n_441),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_692),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_441),
.B(n_445),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_578),
.B(n_644),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_660),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_489),
.B(n_537),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_660),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_660),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_652),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_574),
.B(n_601),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_483),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_445),
.B(n_444),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_498),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_692),
.B(n_700),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_483),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_652),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_700),
.B(n_701),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_485),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_711),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_711),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_708),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_708),
.B(n_717),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_537),
.B(n_717),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_438),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_712),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_715),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_485),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_487),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_487),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_586),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_491),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_671),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_496),
.B(n_697),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_491),
.A2(n_494),
.B1(n_564),
.B2(n_553),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_517),
.B(n_519),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_509),
.B(n_510),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_493),
.Y(n_987)
);

INVxp33_ASAP7_75t_L g988 ( 
.A(n_517),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_542),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_477),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_521),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_434),
.B(n_435),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_494),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_494),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_627),
.B(n_629),
.Y(n_995)
);

AO21x2_ASAP7_75t_L g996 ( 
.A1(n_664),
.A2(n_507),
.B(n_499),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_617),
.B(n_633),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_642),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_519),
.B(n_488),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_658),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_662),
.B(n_665),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_488),
.B(n_523),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_697),
.B(n_668),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_677),
.B(n_714),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_682),
.B(n_690),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_694),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_695),
.B(n_705),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_703),
.B(n_707),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_542),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_586),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_570),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_542),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_499),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_507),
.B(n_605),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_512),
.B(n_577),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_661),
.B(n_709),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_586),
.B(n_606),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_490),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_571),
.Y(n_1019)
);

NOR2x1p5_ASAP7_75t_L g1020 ( 
.A(n_512),
.B(n_572),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_512),
.B(n_577),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_530),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_661),
.B(n_709),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_530),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_532),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_575),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_581),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_658),
.A2(n_688),
.B1(n_585),
.B2(n_608),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_542),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_582),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_584),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_598),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_688),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_532),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_606),
.Y(n_1035)
);

AND2x6_ASAP7_75t_L g1036 ( 
.A(n_554),
.B(n_577),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_535),
.B(n_576),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_535),
.B(n_576),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_606),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_603),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_554),
.B(n_588),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_604),
.B(n_572),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_606),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_612),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_539),
.B(n_587),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_612),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_539),
.B(n_587),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_546),
.B(n_569),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_554),
.B(n_588),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_546),
.B(n_589),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_549),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_572),
.B(n_588),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_612),
.B(n_589),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_505),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_549),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_612),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_550),
.B(n_552),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_550),
.B(n_552),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_558),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_558),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_559),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_559),
.B(n_560),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_560),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_562),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_SL g1065 ( 
.A(n_562),
.B(n_563),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_563),
.B(n_568),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_639),
.A2(n_568),
.B1(n_569),
.B2(n_580),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_580),
.Y(n_1068)
);

AND2x2_ASAP7_75t_SL g1069 ( 
.A(n_592),
.B(n_593),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_592),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_593),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_594),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_594),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_596),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_596),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_605),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_607),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_639),
.A2(n_607),
.B1(n_610),
.B2(n_595),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_610),
.B(n_597),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_609),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_728),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_807),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_780),
.B(n_609),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_729),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_845),
.B(n_923),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_877),
.B(n_896),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_L g1087 ( 
.A(n_740),
.B(n_744),
.C(n_947),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_735),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_815),
.B(n_828),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_887),
.B(n_904),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_727),
.Y(n_1091)
);

NOR2x1p5_ASAP7_75t_L g1092 ( 
.A(n_720),
.B(n_730),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_810),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_824),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_936),
.B(n_928),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_780),
.A2(n_901),
.B(n_902),
.C(n_888),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_825),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_829),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_923),
.B(n_928),
.Y(n_1099)
);

AND2x6_ASAP7_75t_SL g1100 ( 
.A(n_836),
.B(n_838),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_776),
.B(n_904),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_868),
.A2(n_768),
.B1(n_776),
.B2(n_956),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_848),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_765),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_859),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_850),
.A2(n_1003),
.B(n_779),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_797),
.B(n_878),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_878),
.B(n_946),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_933),
.A2(n_865),
.B(n_905),
.C(n_793),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_729),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_988),
.B(n_743),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_866),
.B(n_895),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_789),
.B(n_733),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_754),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_861),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_869),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_871),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_866),
.B(n_895),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_873),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_925),
.B(n_793),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_722),
.B(n_821),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_878),
.B(n_946),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1000),
.A2(n_721),
.B1(n_985),
.B2(n_870),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_769),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_925),
.B(n_973),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_879),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_790),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_727),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_867),
.B(n_734),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_721),
.A2(n_985),
.B1(n_870),
.B2(n_1028),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_722),
.B(n_987),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_954),
.A2(n_983),
.B1(n_999),
.B2(n_778),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_987),
.B(n_803),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_795),
.Y(n_1134)
);

NOR2x1p5_ASAP7_75t_L g1135 ( 
.A(n_720),
.B(n_751),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1002),
.A2(n_997),
.B(n_725),
.C(n_742),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_796),
.B(n_804),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_796),
.B(n_804),
.Y(n_1138)
);

AND2x4_ASAP7_75t_SL g1139 ( 
.A(n_809),
.B(n_812),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_799),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_814),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_L g1142 ( 
.A(n_916),
.B(n_1028),
.C(n_857),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_818),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_959),
.A2(n_938),
.B(n_954),
.C(n_971),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_833),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_878),
.B(n_946),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_986),
.B(n_971),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_946),
.B(n_787),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_788),
.B(n_732),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_835),
.B(n_853),
.C(n_959),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_732),
.B(n_755),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_890),
.A2(n_966),
.B1(n_972),
.B2(n_851),
.C(n_854),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_972),
.B(n_739),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_851),
.B(n_854),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_724),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_732),
.B(n_755),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_882),
.B(n_881),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_882),
.B(n_881),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_791),
.B(n_893),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_755),
.B(n_1016),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_782),
.B(n_813),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1023),
.B(n_771),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_726),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_791),
.B(n_893),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_837),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_SL g1166 ( 
.A(n_809),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_741),
.A2(n_748),
.B1(n_749),
.B2(n_745),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_756),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_778),
.B(n_781),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_849),
.B(n_975),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_771),
.B(n_770),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_761),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_860),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_975),
.B(n_976),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_976),
.B(n_773),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_781),
.A2(n_1033),
.B1(n_950),
.B2(n_774),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_763),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_771),
.B(n_770),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_875),
.B(n_910),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_852),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_771),
.B(n_770),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_930),
.B(n_811),
.Y(n_1182)
);

INVx8_ASAP7_75t_L g1183 ( 
.A(n_841),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_750),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_766),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_984),
.B(n_767),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_772),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_883),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_984),
.B(n_775),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_826),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_784),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_792),
.B(n_816),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_817),
.B(n_839),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_785),
.B(n_786),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_884),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_783),
.A2(n_733),
.B1(n_737),
.B2(n_958),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_794),
.A2(n_798),
.B1(n_805),
.B2(n_802),
.Y(n_1197)
);

NOR2x1p5_ASAP7_75t_L g1198 ( 
.A(n_903),
.B(n_982),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_792),
.B(n_816),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_792),
.B(n_816),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_832),
.B(n_886),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_885),
.Y(n_1202)
);

NAND2x1p5_ASAP7_75t_L g1203 ( 
.A(n_750),
.B(n_762),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_846),
.B(n_872),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_852),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1073),
.B(n_1013),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_892),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_832),
.B(n_886),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1013),
.B(n_1046),
.Y(n_1209)
);

OR2x2_ASAP7_75t_SL g1210 ( 
.A(n_863),
.B(n_747),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_832),
.B(n_886),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_759),
.B(n_806),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_974),
.B(n_822),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_900),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_737),
.B(n_1004),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_757),
.A2(n_960),
.B1(n_783),
.B2(n_731),
.C(n_862),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_891),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1004),
.B(n_1008),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_894),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_897),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_908),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_922),
.B(n_855),
.Y(n_1222)
);

AO221x1_ASAP7_75t_L g1223 ( 
.A1(n_898),
.A2(n_1009),
.B1(n_1044),
.B2(n_1039),
.C(n_1012),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_753),
.Y(n_1224)
);

BUFx8_ASAP7_75t_L g1225 ( 
.A(n_943),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_912),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_L g1227 ( 
.A(n_812),
.B(n_830),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_899),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_757),
.A2(n_808),
.B1(n_819),
.B2(n_800),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_913),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_907),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1008),
.B(n_1069),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1064),
.B(n_1006),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_915),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_917),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1064),
.B(n_1025),
.Y(n_1236)
);

NOR3xp33_ASAP7_75t_L g1237 ( 
.A(n_926),
.B(n_876),
.C(n_746),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_911),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_920),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1025),
.B(n_1005),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1007),
.B(n_998),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_856),
.A2(n_789),
.B1(n_723),
.B2(n_827),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_921),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_918),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_937),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_841),
.B(n_847),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_841),
.B(n_847),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_L g1248 ( 
.A(n_1036),
.B(n_826),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_830),
.B(n_858),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_898),
.B(n_906),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_889),
.B(n_992),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_942),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_L g1253 ( 
.A(n_874),
.B(n_957),
.C(n_914),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_889),
.B(n_992),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_898),
.B(n_906),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_924),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_927),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_844),
.Y(n_1258)
);

INVx4_ASAP7_75t_SL g1259 ( 
.A(n_764),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_906),
.B(n_989),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_889),
.B(n_995),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_858),
.B(n_1020),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_989),
.B(n_1009),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_989),
.B(n_1009),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_762),
.B(n_777),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_808),
.A2(n_819),
.B(n_1049),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_826),
.Y(n_1267)
);

INVxp33_ASAP7_75t_L g1268 ( 
.A(n_1056),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_L g1269 ( 
.A(n_1036),
.B(n_826),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_753),
.B(n_960),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1036),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_929),
.A2(n_968),
.B1(n_941),
.B2(n_940),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_995),
.B(n_1001),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1012),
.B(n_1039),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1001),
.B(n_1015),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_949),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1015),
.B(n_1021),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_753),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_952),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1021),
.B(n_1041),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_934),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_777),
.B(n_874),
.Y(n_1282)
);

NAND2xp33_ASAP7_75t_L g1283 ( 
.A(n_1036),
.B(n_831),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_945),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_931),
.B(n_944),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_990),
.Y(n_1286)
);

OAI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_752),
.A2(n_955),
.B(n_1052),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1041),
.B(n_820),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1017),
.A2(n_1042),
.B(n_1079),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_914),
.B(n_957),
.Y(n_1290)
);

BUFx2_ASAP7_75t_SL g1291 ( 
.A(n_943),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_820),
.B(n_834),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_948),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_834),
.B(n_840),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_969),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1029),
.A2(n_1043),
.B(n_1045),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1012),
.B(n_1039),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_932),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_932),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1044),
.B(n_864),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_961),
.A2(n_965),
.B1(n_977),
.B2(n_978),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1044),
.B(n_864),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_970),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_962),
.A2(n_991),
.B1(n_951),
.B2(n_831),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_840),
.B(n_842),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_842),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_909),
.B(n_939),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_843),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_L g1309 ( 
.A(n_831),
.B(n_951),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_843),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_993),
.B(n_994),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_979),
.A2(n_981),
.B1(n_1032),
.B2(n_1030),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_964),
.B(n_967),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_964),
.B(n_967),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1011),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_752),
.A2(n_1031),
.B(n_1040),
.C(n_1027),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1078),
.B(n_1067),
.C(n_1019),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1026),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_909),
.B(n_939),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_801),
.B(n_963),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_831),
.B(n_935),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1022),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_801),
.B(n_963),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_980),
.B(n_1010),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1056),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1055),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_980),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1068),
.B(n_1076),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1024),
.A2(n_1072),
.B1(n_1077),
.B2(n_1051),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1061),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1034),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_880),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_935),
.B(n_1043),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_880),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1035),
.B(n_1010),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1059),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1060),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1063),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1029),
.B(n_1062),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_953),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1065),
.B(n_823),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1071),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_SL g1346 ( 
.A(n_764),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_823),
.B(n_1062),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_919),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_919),
.B(n_1038),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1075),
.A2(n_1074),
.B1(n_1014),
.B2(n_1066),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_736),
.B(n_1014),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_962),
.B(n_951),
.Y(n_1352)
);

INVxp33_ASAP7_75t_L g1353 ( 
.A(n_736),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_962),
.B(n_951),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1038),
.B(n_1047),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_953),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_962),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_L g1360 ( 
.A(n_953),
.B(n_764),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1048),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_953),
.B(n_1050),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1050),
.A2(n_1066),
.B1(n_1080),
.B2(n_1054),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_764),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_L g1365 ( 
.A(n_758),
.B(n_1053),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1018),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1067),
.B(n_1078),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_760),
.B(n_719),
.Y(n_1368)
);

AND2x2_ASAP7_75t_SL g1369 ( 
.A(n_719),
.B(n_738),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_996),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_719),
.B(n_738),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_719),
.B(n_738),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_728),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_780),
.B(n_776),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_845),
.A2(n_657),
.B1(n_768),
.B2(n_333),
.Y(n_1375)
);

AND2x2_ASAP7_75t_SL g1376 ( 
.A(n_768),
.B(n_845),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_727),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_877),
.B(n_896),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_807),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_780),
.B(n_776),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_778),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_807),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_728),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_754),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_723),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_877),
.B(n_896),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_807),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_877),
.B(n_896),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_807),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_780),
.A2(n_904),
.B(n_896),
.C(n_797),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_728),
.Y(n_1391)
);

NOR2xp67_ASAP7_75t_L g1392 ( 
.A(n_720),
.B(n_531),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_728),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_936),
.A2(n_474),
.B1(n_464),
.B2(n_887),
.C(n_613),
.Y(n_1394)
);

AND2x6_ASAP7_75t_L g1395 ( 
.A(n_780),
.B(n_789),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_780),
.B(n_776),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_877),
.B(n_896),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_877),
.B(n_323),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_877),
.B(n_896),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_727),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_780),
.B(n_776),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_877),
.B(n_896),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_877),
.B(n_323),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_778),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_807),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_728),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_877),
.B(n_323),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_878),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_807),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_877),
.B(n_896),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_877),
.B(n_896),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_877),
.B(n_896),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_877),
.B(n_896),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_L g1416 ( 
.A(n_720),
.B(n_531),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_780),
.B(n_776),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_807),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_727),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_877),
.B(n_896),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_877),
.B(n_896),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_877),
.B(n_896),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_793),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_845),
.A2(n_657),
.B1(n_768),
.B2(n_333),
.Y(n_1424)
);

BUFx5_ASAP7_75t_L g1425 ( 
.A(n_1036),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_807),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_780),
.B(n_776),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_729),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_877),
.B(n_896),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_878),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_727),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_877),
.B(n_323),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_877),
.B(n_323),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_780),
.B(n_776),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_728),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_728),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1438)
);

NAND2xp33_ASAP7_75t_L g1439 ( 
.A(n_947),
.B(n_1036),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_720),
.B(n_895),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_L g1441 ( 
.A(n_947),
.B(n_1036),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_877),
.B(n_896),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_877),
.B(n_896),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_947),
.B(n_1036),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_807),
.Y(n_1445)
);

AND2x6_ASAP7_75t_SL g1446 ( 
.A(n_836),
.B(n_838),
.Y(n_1446)
);

AO21x1_ASAP7_75t_L g1447 ( 
.A1(n_776),
.A2(n_780),
.B(n_904),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_877),
.B(n_323),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_754),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_SL g1450 ( 
.A(n_809),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_780),
.B(n_776),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1036),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_720),
.B(n_895),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_877),
.B(n_896),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_812),
.B(n_513),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_754),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_728),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_845),
.B(n_548),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_727),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_877),
.B(n_896),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_877),
.B(n_896),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_780),
.B(n_776),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_L g1463 ( 
.A(n_947),
.B(n_1036),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_878),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_877),
.B(n_896),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_877),
.B(n_947),
.C(n_780),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_780),
.B(n_776),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_877),
.B(n_896),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_877),
.B(n_323),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_780),
.B(n_776),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_877),
.B(n_896),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_728),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_877),
.B(n_323),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1036),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_780),
.B(n_776),
.Y(n_1475)
);

AO22x2_ASAP7_75t_L g1476 ( 
.A1(n_985),
.A2(n_619),
.B1(n_453),
.B2(n_475),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_877),
.B(n_896),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_780),
.B(n_776),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_L g1480 ( 
.A(n_877),
.B(n_744),
.C(n_740),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_877),
.B(n_896),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_877),
.B(n_896),
.Y(n_1482)
);

INVxp33_ASAP7_75t_L g1483 ( 
.A(n_754),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_807),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_727),
.Y(n_1485)
);

NOR3xp33_ASAP7_75t_L g1486 ( 
.A(n_877),
.B(n_744),
.C(n_740),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_877),
.B(n_896),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_728),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_780),
.B(n_776),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_877),
.B(n_947),
.C(n_780),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_845),
.B(n_548),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_728),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_845),
.A2(n_657),
.B1(n_768),
.B2(n_333),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_728),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_SL g1495 ( 
.A(n_809),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_878),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_877),
.B(n_896),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_877),
.B(n_896),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_877),
.B(n_896),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_727),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_877),
.B(n_896),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_SL g1503 ( 
.A(n_730),
.B(n_328),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_877),
.B(n_896),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_728),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_877),
.B(n_896),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_780),
.B(n_776),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_778),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_877),
.B(n_896),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_728),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_877),
.B(n_896),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_877),
.B(n_323),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_727),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_727),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_727),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_877),
.B(n_323),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_728),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_728),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_877),
.B(n_323),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_938),
.B(n_522),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_878),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_877),
.B(n_896),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_728),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_780),
.B(n_776),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_728),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_877),
.B(n_323),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_877),
.B(n_896),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_845),
.B(n_548),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_877),
.B(n_896),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_877),
.B(n_896),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_877),
.B(n_323),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_728),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_730),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_807),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_938),
.B(n_522),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_754),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_878),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_728),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_793),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_728),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_812),
.B(n_513),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_807),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_727),
.Y(n_1544)
);

NOR3xp33_ASAP7_75t_L g1545 ( 
.A(n_877),
.B(n_744),
.C(n_740),
.Y(n_1545)
);

INVx8_ASAP7_75t_L g1546 ( 
.A(n_841),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_780),
.A2(n_904),
.B(n_896),
.C(n_797),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_877),
.B(n_896),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_877),
.B(n_896),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_877),
.B(n_323),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_807),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_904),
.A2(n_901),
.B(n_888),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_768),
.B(n_845),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_754),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_727),
.Y(n_1555)
);

NOR2xp67_ASAP7_75t_L g1556 ( 
.A(n_720),
.B(n_531),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_SL g1557 ( 
.A(n_809),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_877),
.B(n_896),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_877),
.B(n_896),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_877),
.B(n_896),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_780),
.B(n_776),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_723),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_727),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_SL g1564 ( 
.A(n_809),
.Y(n_1564)
);

NAND2xp33_ASAP7_75t_L g1565 ( 
.A(n_947),
.B(n_1036),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_727),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_728),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_807),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_780),
.B(n_776),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_728),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_780),
.B(n_776),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_780),
.B(n_776),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_727),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_877),
.B(n_896),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_877),
.B(n_323),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_728),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_877),
.B(n_323),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_877),
.B(n_323),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_936),
.A2(n_326),
.B1(n_331),
.B2(n_323),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_877),
.B(n_896),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_728),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_807),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_1375),
.B2(n_1493),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1366),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1466),
.B(n_1490),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1113),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1366),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1102),
.B(n_1390),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1190),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1086),
.B(n_1378),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1386),
.B(n_1388),
.Y(n_1592)
);

AO22x1_ASAP7_75t_L g1593 ( 
.A1(n_1395),
.A2(n_1480),
.B1(n_1545),
.B2(n_1486),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_1424),
.B2(n_1087),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1169),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1306),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1598)
);

INVx5_ASAP7_75t_L g1599 ( 
.A(n_1183),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1398),
.B(n_1403),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1308),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1190),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1271),
.B(n_1452),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1308),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1179),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1113),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1310),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1452),
.B(n_1474),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1190),
.Y(n_1611)
);

BUFx4f_ASAP7_75t_L g1612 ( 
.A(n_1183),
.Y(n_1612)
);

AOI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1374),
.A2(n_1396),
.B(n_1380),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1407),
.B(n_1432),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1183),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1370),
.Y(n_1616)
);

AND2x6_ASAP7_75t_L g1617 ( 
.A(n_1357),
.B(n_1346),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1394),
.A2(n_1395),
.B1(n_1380),
.B2(n_1374),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1183),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1434),
.B(n_1469),
.C(n_1448),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1546),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1361),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1473),
.B(n_1512),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1402),
.B(n_1412),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1236),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1396),
.A2(n_1401),
.B1(n_1427),
.B2(n_1417),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1401),
.A2(n_1417),
.B1(n_1435),
.B2(n_1427),
.Y(n_1627)
);

AND2x6_ASAP7_75t_L g1628 ( 
.A(n_1357),
.B(n_1346),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1435),
.A2(n_1462),
.B(n_1451),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1370),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1546),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1517),
.B(n_1520),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1534),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1546),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1395),
.A2(n_1462),
.B1(n_1467),
.B2(n_1451),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1467),
.A2(n_1470),
.B1(n_1479),
.B2(n_1475),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1546),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1415),
.B(n_1420),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1343),
.B(n_1452),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1489),
.A2(n_1525),
.B1(n_1561),
.B2(n_1507),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1081),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1088),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1355),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_SL g1645 ( 
.A(n_1262),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1381),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1355),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1346),
.B(n_1129),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1429),
.B(n_1442),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1443),
.B(n_1454),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1474),
.B(n_1330),
.Y(n_1652)
);

O2A1O1Ixp5_ASAP7_75t_L g1653 ( 
.A1(n_1489),
.A2(n_1507),
.B(n_1561),
.C(n_1525),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1356),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1562),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1385),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1404),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1369),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_L g1659 ( 
.A(n_1474),
.B(n_1364),
.Y(n_1659)
);

BUFx12f_ASAP7_75t_L g1660 ( 
.A(n_1385),
.Y(n_1660)
);

BUFx4f_ASAP7_75t_L g1661 ( 
.A(n_1113),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1104),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1356),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1562),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1359),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1460),
.B(n_1461),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1465),
.B(n_1468),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1104),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1471),
.B(n_1478),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1569),
.A2(n_1572),
.B1(n_1571),
.B2(n_1395),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1571),
.A2(n_1572),
.B1(n_1395),
.B2(n_1101),
.Y(n_1671)
);

XNOR2xp5_ASAP7_75t_L g1672 ( 
.A(n_1210),
.B(n_1408),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1359),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1458),
.B(n_1491),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1194),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1225),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1481),
.B(n_1482),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1101),
.A2(n_1095),
.B1(n_1447),
.B2(n_1527),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1487),
.B(n_1497),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1532),
.B(n_1550),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1124),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1575),
.B(n_1577),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1223),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1127),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1127),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1578),
.B(n_1502),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1134),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1504),
.B(n_1506),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1509),
.B(n_1511),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_SL g1692 ( 
.A(n_1285),
.B(n_1089),
.C(n_1523),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1425),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1531),
.B(n_1548),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1508),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1549),
.B(n_1558),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1529),
.B(n_1125),
.Y(n_1698)
);

INVx6_ASAP7_75t_L g1699 ( 
.A(n_1084),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1134),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1559),
.B(n_1560),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1574),
.B(n_1580),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1193),
.B(n_1131),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1337),
.B(n_1130),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1521),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1536),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1225),
.Y(n_1707)
);

OR2x2_ASAP7_75t_SL g1708 ( 
.A(n_1121),
.B(n_1112),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1133),
.B(n_1114),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1338),
.B(n_1358),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1384),
.B(n_1449),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1140),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1140),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1141),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1141),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1153),
.B(n_1085),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1327),
.B(n_1343),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1456),
.B(n_1537),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1139),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1106),
.A2(n_1441),
.B(n_1439),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1143),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1425),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1136),
.A2(n_1441),
.B(n_1444),
.C(n_1439),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1483),
.B(n_1409),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1143),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1554),
.B(n_1147),
.Y(n_1726)
);

NAND2x1p5_ASAP7_75t_L g1727 ( 
.A(n_1344),
.B(n_1338),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1455),
.B(n_1542),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1145),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1132),
.B(n_1216),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1455),
.B(n_1542),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1213),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1128),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1483),
.B(n_1433),
.Y(n_1734)
);

NAND2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1503),
.B(n_1092),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1145),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1438),
.B(n_1477),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1165),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1165),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1225),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1425),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1139),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1173),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1455),
.B(n_1542),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1501),
.B(n_1516),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1118),
.B(n_1240),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1173),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1188),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1410),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1142),
.B(n_1463),
.C(n_1444),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1579),
.B(n_1423),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1176),
.B(n_1144),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1540),
.B(n_1273),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1113),
.A2(n_1476),
.B1(n_1565),
.B2(n_1463),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1425),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1410),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1188),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1196),
.B(n_1109),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1195),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1195),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1217),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1113),
.A2(n_1152),
.B1(n_1565),
.B2(n_1476),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_SL g1764 ( 
.A(n_1287),
.B(n_1222),
.C(n_1290),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1099),
.B(n_1100),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1182),
.B(n_1204),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1325),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1369),
.B(n_1108),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1446),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1425),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1123),
.B(n_1155),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1425),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1410),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_SL g1774 ( 
.A(n_1242),
.B(n_1150),
.C(n_1096),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1161),
.B(n_1128),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1159),
.B(n_1164),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1175),
.B(n_1304),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1241),
.B(n_1206),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1217),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1219),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1275),
.B(n_1251),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1219),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1224),
.A2(n_1278),
.B1(n_1453),
.B2(n_1440),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_SL g1784 ( 
.A(n_1552),
.B(n_1135),
.C(n_1209),
.Y(n_1784)
);

O2A1O1Ixp5_ASAP7_75t_L g1785 ( 
.A1(n_1083),
.A2(n_1149),
.B(n_1148),
.C(n_1107),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1113),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_R g1787 ( 
.A(n_1419),
.B(n_1485),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1410),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1321),
.B(n_1476),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1218),
.B(n_1170),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1220),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1298),
.A2(n_1220),
.B1(n_1231),
.B2(n_1228),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1228),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1163),
.B(n_1168),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1215),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1231),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1455),
.B(n_1542),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1238),
.A2(n_1243),
.B1(n_1245),
.B2(n_1239),
.Y(n_1799)
);

BUFx12f_ASAP7_75t_L g1800 ( 
.A(n_1198),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1082),
.B(n_1093),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1262),
.B(n_1336),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1262),
.B(n_1336),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1172),
.B(n_1177),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1094),
.B(n_1097),
.Y(n_1805)
);

OR2x6_ASAP7_75t_L g1806 ( 
.A(n_1342),
.B(n_1262),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1098),
.B(n_1103),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1212),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1238),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1430),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1315),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1105),
.B(n_1115),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1239),
.Y(n_1813)
);

NAND2x1p5_ASAP7_75t_L g1814 ( 
.A(n_1108),
.B(n_1122),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1243),
.Y(n_1816)
);

O2A1O1Ixp33_ASAP7_75t_L g1817 ( 
.A1(n_1229),
.A2(n_1237),
.B(n_1107),
.C(n_1316),
.Y(n_1817)
);

OR2x2_ASAP7_75t_SL g1818 ( 
.A(n_1258),
.B(n_1232),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1245),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1252),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1430),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1252),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1119),
.B(n_1126),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1277),
.B(n_1280),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1425),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1336),
.B(n_1282),
.Y(n_1826)
);

BUFx8_ASAP7_75t_L g1827 ( 
.A(n_1166),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1430),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1276),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1379),
.B(n_1382),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1440),
.B(n_1453),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1387),
.B(n_1389),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1440),
.A2(n_1453),
.B1(n_1270),
.B2(n_1162),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1162),
.A2(n_1137),
.B1(n_1138),
.B2(n_1283),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1405),
.B(n_1411),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1248),
.A2(n_1269),
.B(n_1283),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1276),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1279),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_SL g1840 ( 
.A(n_1253),
.B(n_1286),
.C(n_1261),
.Y(n_1840)
);

AND2x2_ASAP7_75t_SL g1841 ( 
.A(n_1360),
.B(n_1269),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1279),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1309),
.A2(n_1360),
.B(n_1149),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1186),
.B(n_1189),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1299),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1254),
.B(n_1288),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1191),
.B(n_1418),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1295),
.A2(n_1488),
.B1(n_1581),
.B2(n_1576),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1426),
.B(n_1445),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1289),
.B(n_1266),
.C(n_1311),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1464),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1484),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1464),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1295),
.Y(n_1854)
);

INVx5_ASAP7_75t_L g1855 ( 
.A(n_1464),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1535),
.B(n_1543),
.Y(n_1856)
);

AND3x1_ASAP7_75t_L g1857 ( 
.A(n_1091),
.B(n_1400),
.C(n_1377),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1303),
.A2(n_1488),
.B1(n_1581),
.B2(n_1576),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1551),
.Y(n_1859)
);

NAND2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1122),
.B(n_1146),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1373),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1496),
.Y(n_1862)
);

AND2x6_ASAP7_75t_SL g1863 ( 
.A(n_1282),
.B(n_1265),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1373),
.Y(n_1864)
);

OR2x2_ASAP7_75t_SL g1865 ( 
.A(n_1202),
.B(n_1318),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1282),
.B(n_1265),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1419),
.B(n_1485),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1265),
.B(n_1496),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1568),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_SL g1870 ( 
.A(n_1160),
.B(n_1416),
.C(n_1392),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1496),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1383),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1582),
.B(n_1233),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1371),
.A2(n_1368),
.B(n_1319),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1180),
.B(n_1205),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1391),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1362),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1879)
);

AND2x6_ASAP7_75t_SL g1880 ( 
.A(n_1265),
.B(n_1328),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1391),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1291),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1522),
.B(n_1538),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1566),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1522),
.B(n_1538),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1522),
.B(n_1538),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1393),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1522),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1309),
.A2(n_1160),
.B1(n_1556),
.B2(n_1317),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1406),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1246),
.B(n_1247),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1166),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1406),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1436),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1084),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1436),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1566),
.B(n_1573),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1437),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1363),
.A2(n_1351),
.B1(n_1148),
.B2(n_1367),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1292),
.A2(n_1294),
.B(n_1314),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1573),
.B(n_1268),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1166),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1431),
.B(n_1459),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1146),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1326),
.A2(n_1331),
.B1(n_1341),
.B2(n_1515),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1450),
.Y(n_1907)
);

AND2x6_ASAP7_75t_SL g1908 ( 
.A(n_1372),
.B(n_1450),
.Y(n_1908)
);

AND2x6_ASAP7_75t_SL g1909 ( 
.A(n_1450),
.B(n_1495),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1457),
.Y(n_1910)
);

NAND3xp33_ASAP7_75t_L g1911 ( 
.A(n_1349),
.B(n_1365),
.C(n_1350),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1514),
.B(n_1544),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1268),
.B(n_1312),
.C(n_1302),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1084),
.B(n_1110),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1110),
.B(n_1184),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1555),
.A2(n_1563),
.B1(n_1353),
.B2(n_1227),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1457),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1207),
.B(n_1214),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1221),
.B(n_1226),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1230),
.B(n_1234),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1110),
.B(n_1184),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1184),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1192),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1192),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1495),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1472),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1334),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1472),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1235),
.B(n_1244),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1428),
.B(n_1333),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1335),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1348),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1256),
.B(n_1257),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1281),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1199),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1492),
.Y(n_1937)
);

OR2x2_ASAP7_75t_SL g1938 ( 
.A(n_1284),
.B(n_1293),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1494),
.A2(n_1570),
.B1(n_1567),
.B2(n_1505),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1494),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1203),
.Y(n_1941)
);

OR2x2_ASAP7_75t_SL g1942 ( 
.A(n_1495),
.B(n_1557),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1296),
.B(n_1368),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1505),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1428),
.B(n_1249),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1510),
.Y(n_1946)
);

NOR2xp67_ASAP7_75t_L g1947 ( 
.A(n_1428),
.B(n_1181),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1305),
.B(n_1313),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1518),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1557),
.Y(n_1950)
);

BUFx4f_ASAP7_75t_L g1951 ( 
.A(n_1322),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1557),
.Y(n_1952)
);

NOR3xp33_ASAP7_75t_L g1953 ( 
.A(n_1320),
.B(n_1323),
.C(n_1300),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1564),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1518),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1347),
.B(n_1178),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1519),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1171),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1519),
.B(n_1570),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1524),
.Y(n_1961)
);

NOR2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1564),
.B(n_1322),
.Y(n_1962)
);

OR2x6_ASAP7_75t_L g1963 ( 
.A(n_1181),
.B(n_1324),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1151),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1526),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1167),
.A2(n_1197),
.B1(n_1564),
.B2(n_1301),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1533),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1199),
.B(n_1263),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1332),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1539),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1272),
.A2(n_1263),
.B1(n_1200),
.B2(n_1201),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1541),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1339),
.B(n_1345),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1200),
.B(n_1264),
.C(n_1201),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1208),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1339),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1208),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1340),
.B(n_1329),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1156),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1211),
.B(n_1250),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1211),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1250),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1255),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1260),
.B(n_1264),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1274),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1297),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1297),
.B(n_1466),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1366),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1398),
.B(n_1403),
.Y(n_1990)
);

INVx4_ASAP7_75t_L g1991 ( 
.A(n_1546),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1366),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1190),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1086),
.B(n_1378),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1376),
.B(n_1553),
.Y(n_1996)
);

O2A1O1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1390),
.A2(n_1547),
.B(n_1480),
.C(n_1545),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1086),
.B(n_1378),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1366),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1190),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1385),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1190),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1366),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1366),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1190),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1259),
.B(n_1267),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1366),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1534),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1466),
.A2(n_1490),
.B1(n_1374),
.B2(n_1396),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1183),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1374),
.A2(n_1396),
.B(n_1380),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1376),
.B(n_439),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1366),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1366),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1366),
.Y(n_2022)
);

AO22x1_ASAP7_75t_L g2023 ( 
.A1(n_1395),
.A2(n_1480),
.B1(n_1545),
.B2(n_1486),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1366),
.Y(n_2025)
);

CKINVDCx8_ASAP7_75t_R g2026 ( 
.A(n_1291),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1374),
.A2(n_1396),
.B(n_1380),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1366),
.Y(n_2028)
);

NOR2x2_ASAP7_75t_L g2029 ( 
.A(n_1262),
.B(n_616),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1366),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1366),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1366),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1546),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1366),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2037)
);

INVxp67_ASAP7_75t_L g2038 ( 
.A(n_1169),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1390),
.A2(n_1547),
.B(n_1480),
.C(n_1545),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1183),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1183),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1366),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_1190),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1366),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2048)
);

BUFx4f_ASAP7_75t_L g2049 ( 
.A(n_1183),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2050)
);

INVxp67_ASAP7_75t_SL g2051 ( 
.A(n_1236),
.Y(n_2051)
);

INVx5_ASAP7_75t_L g2052 ( 
.A(n_1183),
.Y(n_2052)
);

AND2x6_ASAP7_75t_L g2053 ( 
.A(n_1267),
.B(n_1190),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1366),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1183),
.Y(n_2057)
);

BUFx4f_ASAP7_75t_L g2058 ( 
.A(n_1183),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1183),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1534),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2062)
);

INVxp67_ASAP7_75t_SL g2063 ( 
.A(n_1236),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1374),
.A2(n_1396),
.B(n_1380),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1366),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1366),
.Y(n_2070)
);

NOR3xp33_ASAP7_75t_SL g2071 ( 
.A(n_1398),
.B(n_326),
.C(n_323),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_1190),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1183),
.Y(n_2073)
);

INVx2_ASAP7_75t_SL g2074 ( 
.A(n_1190),
.Y(n_2074)
);

BUFx4f_ASAP7_75t_L g2075 ( 
.A(n_1183),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2076)
);

OAI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1466),
.A2(n_1490),
.B(n_1380),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1534),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1366),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1366),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_L g2082 ( 
.A(n_1466),
.B(n_1490),
.C(n_1390),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1534),
.Y(n_2085)
);

AND2x6_ASAP7_75t_SL g2086 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1366),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2090)
);

NOR2x1p5_ASAP7_75t_L g2091 ( 
.A(n_1128),
.B(n_448),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1366),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1190),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1366),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1190),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1190),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1190),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_SL g2100 ( 
.A(n_1480),
.B(n_1545),
.C(n_1486),
.Y(n_2100)
);

INVx4_ASAP7_75t_L g2101 ( 
.A(n_1546),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1190),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1366),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1366),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_1190),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_R g2106 ( 
.A(n_1534),
.B(n_327),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1366),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1366),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1366),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1259),
.B(n_1267),
.Y(n_2111)
);

AND2x4_ASAP7_75t_SL g2112 ( 
.A(n_1190),
.B(n_1452),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_1385),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1113),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_1169),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1534),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1366),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1366),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_1183),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1366),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1366),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1534),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1366),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1183),
.Y(n_2132)
);

AND2x6_ASAP7_75t_SL g2133 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1366),
.Y(n_2134)
);

BUFx12f_ASAP7_75t_L g2135 ( 
.A(n_1385),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1366),
.Y(n_2137)
);

INVx2_ASAP7_75t_SL g2138 ( 
.A(n_1190),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1576),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1366),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2142)
);

AO22x1_ASAP7_75t_L g2143 ( 
.A1(n_1395),
.A2(n_1480),
.B1(n_1545),
.B2(n_1486),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1366),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1366),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1366),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1366),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1534),
.Y(n_2152)
);

AND3x2_ASAP7_75t_SL g2153 ( 
.A(n_1447),
.B(n_1553),
.C(n_1376),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1366),
.Y(n_2154)
);

NOR3xp33_ASAP7_75t_SL g2155 ( 
.A(n_1398),
.B(n_326),
.C(n_323),
.Y(n_2155)
);

NOR2x2_ASAP7_75t_L g2156 ( 
.A(n_1262),
.B(n_616),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1366),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1190),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_1190),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2160)
);

NOR2x1p5_ASAP7_75t_L g2161 ( 
.A(n_1128),
.B(n_448),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1366),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1183),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1366),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2171)
);

INVx5_ASAP7_75t_L g2172 ( 
.A(n_1183),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1366),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_1102),
.A2(n_1490),
.B1(n_1466),
.B2(n_1086),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_1374),
.A2(n_1396),
.B(n_1380),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1534),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1366),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1366),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1366),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_SL g2185 ( 
.A(n_1480),
.B(n_1545),
.C(n_1486),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_1090),
.B(n_1154),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1366),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_1190),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2190)
);

BUFx12f_ASAP7_75t_L g2191 ( 
.A(n_1385),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_1376),
.A2(n_1553),
.B1(n_845),
.B2(n_333),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_1190),
.Y(n_2193)
);

OAI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_1102),
.A2(n_1490),
.B1(n_1466),
.B2(n_1086),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1366),
.Y(n_2198)
);

INVx5_ASAP7_75t_L g2199 ( 
.A(n_1183),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_1190),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1366),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_1099),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1366),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1366),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1366),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1366),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1366),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1366),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1576),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_1099),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2215)
);

CKINVDCx20_ASAP7_75t_R g2216 ( 
.A(n_1385),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1366),
.Y(n_2218)
);

INVx1_ASAP7_75t_SL g2219 ( 
.A(n_1521),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1366),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1366),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_1259),
.B(n_1267),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_1466),
.A2(n_1490),
.B1(n_1374),
.B2(n_1396),
.Y(n_2223)
);

HB1xp67_ASAP7_75t_L g2224 ( 
.A(n_1099),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1259),
.B(n_1267),
.Y(n_2225)
);

BUFx12f_ASAP7_75t_L g2226 ( 
.A(n_1385),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1366),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_1190),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1394),
.A2(n_1087),
.B1(n_1490),
.B2(n_1466),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_1398),
.B(n_1403),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1376),
.B(n_1553),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1366),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1366),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1366),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1099),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1366),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1366),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_1190),
.Y(n_2239)
);

INVxp67_ASAP7_75t_L g2240 ( 
.A(n_1169),
.Y(n_2240)
);

INVx5_ASAP7_75t_L g2241 ( 
.A(n_1183),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1466),
.B(n_1490),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_1546),
.Y(n_2243)
);

INVx2_ASAP7_75t_SL g2244 ( 
.A(n_1190),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_1099),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1086),
.B(n_1378),
.Y(n_2246)
);

HB1xp67_ASAP7_75t_L g2247 ( 
.A(n_1099),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_1521),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1366),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1366),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2251)
);

O2A1O1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2100),
.A2(n_2185),
.B(n_1614),
.C(n_1623),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2253)
);

A2O1A1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_1999),
.A2(n_2018),
.B(n_2044),
.C(n_2042),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1702),
.B(n_1687),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2176),
.B(n_2194),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1591),
.B(n_1592),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_1997),
.A2(n_2039),
.B(n_1723),
.Y(n_2258)
);

OAI321xp33_ASAP7_75t_L g2259 ( 
.A1(n_1999),
.A2(n_2044),
.A3(n_2018),
.B1(n_2171),
.B2(n_2167),
.C(n_2042),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2014),
.A2(n_2223),
.B(n_1901),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1598),
.B(n_1624),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1678),
.B(n_2019),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_1976),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1730),
.A2(n_2167),
.B1(n_2196),
.B2(n_2171),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_1996),
.B(n_2002),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2083),
.A2(n_2108),
.B1(n_2150),
.B2(n_2145),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1836),
.A2(n_1641),
.B(n_2082),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1996),
.B(n_2002),
.Y(n_2268)
);

INVx4_ASAP7_75t_L g2269 ( 
.A(n_1863),
.Y(n_2269)
);

CKINVDCx10_ASAP7_75t_R g2270 ( 
.A(n_1655),
.Y(n_2270)
);

A2O1A1Ixp33_ASAP7_75t_L g2271 ( 
.A1(n_2230),
.A2(n_2196),
.B(n_2201),
.C(n_1678),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1632),
.B(n_1639),
.Y(n_2272)
);

O2A1O1Ixp5_ASAP7_75t_L g2273 ( 
.A1(n_1589),
.A2(n_1593),
.B(n_2143),
.C(n_2023),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_1693),
.Y(n_2274)
);

A2O1A1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2201),
.A2(n_2230),
.B(n_1594),
.C(n_1750),
.Y(n_2275)
);

INVxp67_ASAP7_75t_L g2276 ( 
.A(n_1808),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1648),
.B(n_1650),
.Y(n_2277)
);

NOR2xp67_ASAP7_75t_L g2278 ( 
.A(n_1750),
.B(n_1874),
.Y(n_2278)
);

INVxp67_ASAP7_75t_L g2279 ( 
.A(n_1711),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1666),
.B(n_1667),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_2053),
.Y(n_2281)
);

AOI21x1_ASAP7_75t_L g2282 ( 
.A1(n_1593),
.A2(n_2143),
.B(n_2023),
.Y(n_2282)
);

OAI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2082),
.A2(n_2077),
.B(n_2010),
.Y(n_2283)
);

AO21x1_ASAP7_75t_L g2284 ( 
.A1(n_1759),
.A2(n_1817),
.B(n_1586),
.Y(n_2284)
);

A2O1A1Ixp33_ASAP7_75t_L g2285 ( 
.A1(n_1600),
.A2(n_1633),
.B(n_1683),
.C(n_1680),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_L g2286 ( 
.A(n_1874),
.B(n_1850),
.Y(n_2286)
);

NAND2x1p5_ASAP7_75t_L g2287 ( 
.A(n_1661),
.B(n_1786),
.Y(n_2287)
);

O2A1O1Ixp33_ASAP7_75t_L g2288 ( 
.A1(n_1990),
.A2(n_2089),
.B(n_2127),
.C(n_2087),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_1618),
.A2(n_2179),
.B1(n_2189),
.B2(n_2169),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2037),
.B(n_2067),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1661),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2231),
.B(n_1764),
.Y(n_2292)
);

AOI21x1_ASAP7_75t_L g2293 ( 
.A1(n_1629),
.A2(n_2027),
.B(n_2017),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_1911),
.B(n_1774),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_1927),
.B(n_1605),
.Y(n_2295)
);

O2A1O1Ixp33_ASAP7_75t_L g2296 ( 
.A1(n_2024),
.A2(n_2056),
.B(n_2069),
.C(n_2048),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2084),
.A2(n_2117),
.B(n_2115),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1677),
.B(n_1681),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2066),
.A2(n_2178),
.B(n_2130),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2125),
.A2(n_2142),
.B(n_2139),
.Y(n_2300)
);

AOI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2163),
.A2(n_2165),
.B(n_2164),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_1626),
.A2(n_1627),
.B1(n_1637),
.B2(n_2166),
.Y(n_2302)
);

AOI21x1_ASAP7_75t_L g2303 ( 
.A1(n_2190),
.A2(n_2213),
.B(n_2212),
.Y(n_2303)
);

BUFx3_ASAP7_75t_L g2304 ( 
.A(n_2053),
.Y(n_2304)
);

NOR2x1p5_ASAP7_75t_SL g2305 ( 
.A(n_1644),
.B(n_1647),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2228),
.A2(n_2242),
.B(n_1653),
.Y(n_2306)
);

OA22x2_ASAP7_75t_L g2307 ( 
.A1(n_2037),
.A2(n_2067),
.B1(n_2099),
.B2(n_2090),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1616),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_1948),
.A2(n_1841),
.B(n_1613),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1751),
.B(n_1752),
.Y(n_2311)
);

AOI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_1841),
.A2(n_1843),
.B(n_1636),
.Y(n_2312)
);

OAI321xp33_ASAP7_75t_L g2313 ( 
.A1(n_1626),
.A2(n_1627),
.A3(n_1637),
.B1(n_1584),
.B2(n_2192),
.C(n_2160),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1644),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_1724),
.A2(n_1734),
.B1(n_1607),
.B2(n_1737),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_1763),
.A2(n_1670),
.B(n_1671),
.C(n_1620),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_R g2317 ( 
.A(n_1664),
.B(n_1634),
.Y(n_2317)
);

CKINVDCx10_ASAP7_75t_R g2318 ( 
.A(n_1655),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1690),
.B(n_1695),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2086),
.B(n_2133),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1697),
.B(n_1701),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1995),
.B(n_1998),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2086),
.B(n_2133),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1766),
.B(n_1916),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_1841),
.A2(n_1670),
.B(n_1661),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2005),
.B(n_2007),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2015),
.B(n_2032),
.Y(n_2327)
);

O2A1O1Ixp33_ASAP7_75t_SL g2328 ( 
.A1(n_1745),
.A2(n_1669),
.B(n_1679),
.C(n_1651),
.Y(n_2328)
);

NAND3xp33_ASAP7_75t_L g2329 ( 
.A(n_1671),
.B(n_1692),
.C(n_1988),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_1718),
.Y(n_2330)
);

A2O1A1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_1763),
.A2(n_1753),
.B(n_1900),
.C(n_2186),
.Y(n_2331)
);

INVxp67_ASAP7_75t_L g2332 ( 
.A(n_1811),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2033),
.B(n_2040),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2050),
.B(n_2054),
.Y(n_2334)
);

OAI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2059),
.A2(n_2064),
.B1(n_2065),
.B2(n_2062),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2336)
);

CKINVDCx6p67_ASAP7_75t_R g2337 ( 
.A(n_1660),
.Y(n_2337)
);

AOI21xp33_ASAP7_75t_L g2338 ( 
.A1(n_2186),
.A2(n_1966),
.B(n_1911),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2076),
.B(n_2078),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1647),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2098),
.B(n_2120),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2123),
.B(n_2131),
.Y(n_2342)
);

NOR2x1_ASAP7_75t_L g2343 ( 
.A(n_1975),
.B(n_1840),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_1943),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2136),
.B(n_2148),
.Y(n_2345)
);

BUFx4f_ASAP7_75t_L g2346 ( 
.A(n_1617),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1654),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_1943),
.A2(n_1754),
.B(n_1951),
.Y(n_2349)
);

OAI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2151),
.A2(n_2174),
.B1(n_2177),
.B2(n_2175),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_1951),
.A2(n_1834),
.B(n_1914),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2180),
.B(n_2195),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2197),
.B(n_2215),
.Y(n_2353)
);

O2A1O1Ixp33_ASAP7_75t_L g2354 ( 
.A1(n_2217),
.A2(n_2246),
.B(n_1767),
.C(n_2155),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_1755),
.A2(n_1708),
.B1(n_1865),
.B2(n_1672),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_1916),
.B(n_1649),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2013),
.B(n_2061),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1654),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1693),
.Y(n_2359)
);

AOI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_1951),
.A2(n_1834),
.B(n_1915),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_1921),
.A2(n_1777),
.B(n_1958),
.Y(n_2361)
);

AOI21x1_ASAP7_75t_L g2362 ( 
.A1(n_1891),
.A2(n_1846),
.B(n_1981),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2079),
.B(n_2085),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_1873),
.A2(n_1866),
.B(n_1612),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_1616),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1703),
.B(n_1709),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1663),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_1744),
.B(n_1798),
.Y(n_2368)
);

A2O1A1Ixp33_ASAP7_75t_L g2369 ( 
.A1(n_1900),
.A2(n_1906),
.B(n_2099),
.C(n_2090),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1663),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_1726),
.B(n_1791),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_1735),
.B(n_1765),
.C(n_1769),
.Y(n_2372)
);

AO21x1_ASAP7_75t_L g2373 ( 
.A1(n_1781),
.A2(n_1673),
.B(n_1665),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1665),
.Y(n_2374)
);

AND2x4_ASAP7_75t_L g2375 ( 
.A(n_1744),
.B(n_1798),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_1866),
.A2(n_2049),
.B(n_1612),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1673),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1778),
.B(n_1746),
.Y(n_2378)
);

O2A1O1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2071),
.A2(n_1852),
.B(n_1869),
.C(n_1859),
.Y(n_2379)
);

AND2x2_ASAP7_75t_SL g2380 ( 
.A(n_1658),
.B(n_1786),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1746),
.B(n_1595),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_1866),
.A2(n_2049),
.B(n_1612),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2038),
.B(n_2116),
.Y(n_2383)
);

AOI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_1866),
.A2(n_2058),
.B(n_2049),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2118),
.B(n_2128),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2240),
.B(n_1705),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2219),
.B(n_2248),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2075),
.A2(n_1922),
.B(n_1895),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_1895),
.A2(n_1922),
.B(n_1785),
.Y(n_2389)
);

CKINVDCx6p67_ASAP7_75t_R g2390 ( 
.A(n_1660),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1693),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2152),
.B(n_2181),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2205),
.B(n_2232),
.Y(n_2393)
);

OAI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_1889),
.A2(n_1784),
.B(n_1906),
.Y(n_2394)
);

INVx3_ASAP7_75t_SL g2395 ( 
.A(n_1892),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_1706),
.B(n_1824),
.Y(n_2396)
);

O2A1O1Ixp33_ASAP7_75t_L g2397 ( 
.A1(n_1935),
.A2(n_1775),
.B(n_1657),
.C(n_1696),
.Y(n_2397)
);

O2A1O1Ixp5_ASAP7_75t_L g2398 ( 
.A1(n_1968),
.A2(n_1985),
.B(n_1980),
.C(n_1930),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1616),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1698),
.B(n_1605),
.Y(n_2400)
);

O2A1O1Ixp33_ASAP7_75t_SL g2401 ( 
.A1(n_1945),
.A2(n_1903),
.B(n_1925),
.C(n_1907),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1630),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1857),
.B(n_1889),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1585),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_1818),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1698),
.B(n_1790),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1796),
.B(n_2203),
.Y(n_2407)
);

BUFx2_ASAP7_75t_L g2408 ( 
.A(n_1963),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2205),
.B(n_2232),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_1674),
.B(n_1847),
.Y(n_2410)
);

AOI221xp5_ASAP7_75t_L g2411 ( 
.A1(n_1672),
.A2(n_1856),
.B1(n_1807),
.B2(n_1812),
.C(n_1805),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_1771),
.A2(n_1704),
.B1(n_1789),
.B2(n_1674),
.Y(n_2412)
);

NAND2x1p5_ASAP7_75t_L g2413 ( 
.A(n_1599),
.B(n_2052),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1630),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1989),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1989),
.Y(n_2416)
);

NAND3xp33_ASAP7_75t_L g2417 ( 
.A(n_1953),
.B(n_1934),
.C(n_1972),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1992),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2214),
.B(n_2224),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_1963),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2236),
.B(n_2245),
.Y(n_2421)
);

BUFx12f_ASAP7_75t_L g2422 ( 
.A(n_1656),
.Y(n_2422)
);

AO21x2_ASAP7_75t_L g2423 ( 
.A1(n_1992),
.A2(n_2006),
.B(n_2000),
.Y(n_2423)
);

AND2x6_ASAP7_75t_L g2424 ( 
.A(n_1658),
.B(n_1583),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_1693),
.A2(n_1741),
.B(n_1722),
.Y(n_2425)
);

OAI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_1972),
.A2(n_1684),
.B(n_1986),
.Y(n_2426)
);

INVxp33_ASAP7_75t_L g2427 ( 
.A(n_2106),
.Y(n_2427)
);

AND2x6_ASAP7_75t_L g2428 ( 
.A(n_1658),
.B(n_1583),
.Y(n_2428)
);

INVx4_ASAP7_75t_L g2429 ( 
.A(n_1863),
.Y(n_2429)
);

AOI33xp33_ASAP7_75t_L g2430 ( 
.A1(n_1856),
.A2(n_1716),
.A3(n_1847),
.B1(n_1882),
.B2(n_1884),
.B3(n_1622),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2247),
.B(n_1675),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_1587),
.A2(n_2114),
.B(n_1608),
.Y(n_2432)
);

NOR2xp67_ASAP7_75t_L g2433 ( 
.A(n_1821),
.B(n_1855),
.Y(n_2433)
);

NAND2x1p5_ASAP7_75t_L g2434 ( 
.A(n_1599),
.B(n_2052),
.Y(n_2434)
);

BUFx8_ASAP7_75t_L g2435 ( 
.A(n_2003),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_1684),
.A2(n_1987),
.B(n_1622),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_1857),
.B(n_1833),
.Y(n_2437)
);

OA22x2_ASAP7_75t_L g2438 ( 
.A1(n_1833),
.A2(n_1966),
.B1(n_1783),
.B2(n_2153),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_1716),
.B(n_1776),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_1704),
.A2(n_1771),
.B1(n_1783),
.B2(n_1936),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_1789),
.A2(n_1628),
.B1(n_1617),
.B2(n_1658),
.Y(n_2441)
);

AOI21x1_ASAP7_75t_L g2442 ( 
.A1(n_1717),
.A2(n_1978),
.B(n_1947),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_1818),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_1876),
.B(n_1879),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2114),
.A2(n_1947),
.B(n_1826),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_1826),
.A2(n_1741),
.B(n_1722),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_1795),
.B(n_1804),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2053),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1630),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_1826),
.A2(n_1741),
.B(n_1722),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1675),
.B(n_1795),
.Y(n_2451)
);

AOI21x1_ASAP7_75t_L g2452 ( 
.A1(n_1883),
.A2(n_1898),
.B(n_1980),
.Y(n_2452)
);

BUFx4f_ASAP7_75t_L g2453 ( 
.A(n_1617),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2000),
.Y(n_2454)
);

NAND2xp33_ASAP7_75t_SL g2455 ( 
.A(n_1870),
.B(n_1787),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_1804),
.B(n_1838),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_1838),
.B(n_1732),
.Y(n_2457)
);

A2O1A1Ixp33_ASAP7_75t_L g2458 ( 
.A1(n_2153),
.A2(n_1831),
.B(n_1902),
.C(n_1801),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_1826),
.B(n_1905),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2006),
.Y(n_2460)
);

O2A1O1Ixp33_ASAP7_75t_SL g2461 ( 
.A1(n_1615),
.A2(n_1635),
.B(n_1619),
.C(n_1719),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_2053),
.Y(n_2462)
);

OAI21xp33_ASAP7_75t_L g2463 ( 
.A1(n_2153),
.A2(n_1913),
.B(n_1823),
.Y(n_2463)
);

INVx11_ASAP7_75t_L g2464 ( 
.A(n_1800),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_1789),
.A2(n_1628),
.B1(n_1617),
.B2(n_1658),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1646),
.B(n_1815),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1588),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_1927),
.B(n_1789),
.Y(n_2468)
);

BUFx6f_ASAP7_75t_L g2469 ( 
.A(n_1601),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_1756),
.Y(n_2470)
);

AO21x1_ASAP7_75t_L g2471 ( 
.A1(n_1727),
.A2(n_1984),
.B(n_1983),
.Y(n_2471)
);

AOI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_1802),
.A2(n_1803),
.B1(n_1956),
.B2(n_1652),
.Y(n_2472)
);

INVx11_ASAP7_75t_L g2473 ( 
.A(n_1800),
.Y(n_2473)
);

BUFx3_ASAP7_75t_L g2474 ( 
.A(n_2053),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1830),
.B(n_1832),
.Y(n_2475)
);

OAI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_1983),
.A2(n_1984),
.B(n_1849),
.Y(n_2476)
);

INVxp67_ASAP7_75t_SL g2477 ( 
.A(n_1625),
.Y(n_2477)
);

HB1xp67_ASAP7_75t_L g2478 ( 
.A(n_1835),
.Y(n_2478)
);

AO22x1_ASAP7_75t_L g2479 ( 
.A1(n_1617),
.A2(n_1628),
.B1(n_2053),
.B2(n_1597),
.Y(n_2479)
);

OR2x6_ASAP7_75t_SL g2480 ( 
.A(n_1952),
.B(n_1676),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2020),
.B(n_2021),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2053),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_1897),
.B(n_1867),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2051),
.B(n_2063),
.Y(n_2484)
);

NAND3xp33_ASAP7_75t_L g2485 ( 
.A(n_1964),
.B(n_1982),
.C(n_1963),
.Y(n_2485)
);

OAI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_1708),
.A2(n_1865),
.B1(n_1938),
.B2(n_1699),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2020),
.Y(n_2487)
);

BUFx8_ASAP7_75t_L g2488 ( 
.A(n_2003),
.Y(n_2488)
);

O2A1O1Ixp33_ASAP7_75t_L g2489 ( 
.A1(n_1904),
.A2(n_1912),
.B(n_1875),
.C(n_1950),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1918),
.B(n_1919),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_1905),
.B(n_1802),
.Y(n_2491)
);

O2A1O1Ixp33_ASAP7_75t_L g2492 ( 
.A1(n_1950),
.A2(n_1954),
.B(n_1742),
.C(n_1719),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_1733),
.B(n_2026),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1920),
.B(n_1933),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_1740),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_1770),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1588),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_1601),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_1588),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1929),
.B(n_1844),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1929),
.B(n_1844),
.Y(n_2501)
);

OAI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_1923),
.A2(n_1924),
.B(n_1727),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_1770),
.Y(n_2503)
);

BUFx4f_ASAP7_75t_L g2504 ( 
.A(n_1617),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_1772),
.A2(n_1825),
.B(n_1963),
.Y(n_2505)
);

A2O1A1Ixp33_ASAP7_75t_L g2506 ( 
.A1(n_1601),
.A2(n_1659),
.B(n_1956),
.C(n_1597),
.Y(n_2506)
);

A2O1A1Ixp33_ASAP7_75t_L g2507 ( 
.A1(n_1601),
.A2(n_1659),
.B(n_1956),
.C(n_1597),
.Y(n_2507)
);

A2O1A1Ixp33_ASAP7_75t_L g2508 ( 
.A1(n_1956),
.A2(n_1597),
.B(n_1994),
.C(n_1583),
.Y(n_2508)
);

INVx3_ASAP7_75t_L g2509 ( 
.A(n_1772),
.Y(n_2509)
);

A2O1A1Ixp33_ASAP7_75t_L g2510 ( 
.A1(n_1583),
.A2(n_1994),
.B(n_2111),
.C(n_2011),
.Y(n_2510)
);

OAI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_1727),
.A2(n_1959),
.B(n_1860),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_1733),
.B(n_2026),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_1938),
.A2(n_1699),
.B1(n_1806),
.B2(n_1803),
.Y(n_2513)
);

NOR2x1_ASAP7_75t_L g2514 ( 
.A(n_1950),
.B(n_1954),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_1950),
.B(n_1954),
.C(n_1742),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2022),
.B(n_2025),
.Y(n_2516)
);

A2O1A1Ixp33_ASAP7_75t_L g2517 ( 
.A1(n_1994),
.A2(n_2011),
.B(n_2222),
.C(n_2111),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2008),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_1994),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_1596),
.B(n_1602),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_1596),
.B(n_1602),
.Y(n_2521)
);

O2A1O1Ixp33_ASAP7_75t_SL g2522 ( 
.A1(n_1615),
.A2(n_1635),
.B(n_1619),
.C(n_1941),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_1606),
.B(n_1609),
.Y(n_2523)
);

A2O1A1Ixp33_ASAP7_75t_L g2524 ( 
.A1(n_2011),
.A2(n_2111),
.B(n_2225),
.C(n_2222),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_1802),
.A2(n_1803),
.B1(n_1652),
.B2(n_1806),
.Y(n_2525)
);

BUFx3_ASAP7_75t_L g2526 ( 
.A(n_1628),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_1878),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_R g2528 ( 
.A(n_1707),
.B(n_2113),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_1789),
.B(n_1878),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_1905),
.B(n_1803),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2011),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1845),
.B(n_1733),
.Y(n_2532)
);

A2O1A1Ixp33_ASAP7_75t_L g2533 ( 
.A1(n_2111),
.A2(n_2225),
.B(n_2222),
.C(n_1962),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2222),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_1628),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1931),
.B(n_1932),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_1931),
.B(n_1932),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_SL g2538 ( 
.A(n_1628),
.B(n_1645),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2022),
.B(n_2025),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_1905),
.B(n_1868),
.Y(n_2540)
);

NOR2x1_ASAP7_75t_L g2541 ( 
.A(n_1954),
.B(n_1898),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_1868),
.B(n_1941),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_SL g2543 ( 
.A(n_1628),
.B(n_1645),
.Y(n_2543)
);

INVx4_ASAP7_75t_L g2544 ( 
.A(n_2172),
.Y(n_2544)
);

NOR3xp33_ASAP7_75t_L g2545 ( 
.A(n_1828),
.B(n_1862),
.C(n_1851),
.Y(n_2545)
);

OAI22xp5_ASAP7_75t_L g2546 ( 
.A1(n_1699),
.A2(n_1806),
.B1(n_1744),
.B2(n_1798),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2199),
.A2(n_2241),
.B(n_1806),
.Y(n_2547)
);

CKINVDCx10_ASAP7_75t_R g2548 ( 
.A(n_2135),
.Y(n_2548)
);

AOI21xp5_ASAP7_75t_L g2549 ( 
.A1(n_2199),
.A2(n_2241),
.B(n_1806),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2008),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2216),
.B(n_2135),
.Y(n_2551)
);

AOI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2199),
.A2(n_2241),
.B(n_1710),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_1898),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_1710),
.A2(n_1798),
.B(n_1744),
.Y(n_2554)
);

BUFx8_ASAP7_75t_L g2555 ( 
.A(n_2191),
.Y(n_2555)
);

A2O1A1Ixp33_ASAP7_75t_L g2556 ( 
.A1(n_2225),
.A2(n_1962),
.B(n_1959),
.C(n_1652),
.Y(n_2556)
);

INVxp67_ASAP7_75t_L g2557 ( 
.A(n_1652),
.Y(n_2557)
);

O2A1O1Ixp33_ASAP7_75t_L g2558 ( 
.A1(n_2091),
.A2(n_2161),
.B(n_1621),
.C(n_1638),
.Y(n_2558)
);

AOI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_1710),
.A2(n_1604),
.B(n_1868),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2028),
.B(n_2030),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_1710),
.A2(n_1604),
.B(n_1610),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2191),
.B(n_2226),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2028),
.B(n_2030),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_1604),
.A2(n_1610),
.B(n_1640),
.Y(n_2564)
);

AOI21xp5_ASAP7_75t_L g2565 ( 
.A1(n_1610),
.A2(n_1640),
.B(n_2225),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2008),
.Y(n_2566)
);

O2A1O1Ixp33_ASAP7_75t_L g2567 ( 
.A1(n_2091),
.A2(n_2161),
.B(n_1621),
.C(n_1638),
.Y(n_2567)
);

NOR2x1_ASAP7_75t_L g2568 ( 
.A(n_1828),
.B(n_1851),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2226),
.B(n_1827),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2031),
.B(n_2036),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_1610),
.A2(n_1640),
.B(n_1768),
.Y(n_2571)
);

INVx1_ASAP7_75t_SL g2572 ( 
.A(n_2029),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2031),
.B(n_2036),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2045),
.B(n_2047),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_1827),
.B(n_1942),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_1964),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2045),
.B(n_2047),
.Y(n_2577)
);

AND2x2_ASAP7_75t_SL g2578 ( 
.A(n_1991),
.B(n_2035),
.Y(n_2578)
);

OR2x6_ASAP7_75t_SL g2579 ( 
.A(n_1942),
.B(n_1880),
.Y(n_2579)
);

AOI21xp5_ASAP7_75t_L g2580 ( 
.A1(n_1768),
.A2(n_2112),
.B(n_1855),
.Y(n_2580)
);

NAND3xp33_ASAP7_75t_L g2581 ( 
.A(n_1964),
.B(n_1982),
.C(n_1827),
.Y(n_2581)
);

OR2x6_ASAP7_75t_SL g2582 ( 
.A(n_1880),
.B(n_1908),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2055),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2055),
.B(n_2068),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2068),
.B(n_2070),
.Y(n_2585)
);

OAI21xp33_ASAP7_75t_L g2586 ( 
.A1(n_1793),
.A2(n_1860),
.B(n_1814),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2070),
.B(n_2080),
.Y(n_2587)
);

OAI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_1699),
.A2(n_1768),
.B1(n_2035),
.B2(n_1991),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2088),
.B(n_2092),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_1827),
.B(n_1909),
.Y(n_2590)
);

INVx2_ASAP7_75t_SL g2591 ( 
.A(n_1788),
.Y(n_2591)
);

AO21x1_ASAP7_75t_L g2592 ( 
.A1(n_1688),
.A2(n_1860),
.B(n_1814),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2088),
.B(n_2092),
.Y(n_2593)
);

BUFx2_ASAP7_75t_L g2594 ( 
.A(n_1964),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_1964),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_1909),
.B(n_1862),
.Y(n_2596)
);

BUFx12f_ASAP7_75t_L g2597 ( 
.A(n_1908),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2103),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_1871),
.B(n_1788),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2103),
.B(n_2104),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2104),
.B(n_2107),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2107),
.B(n_2110),
.Y(n_2602)
);

BUFx4f_ASAP7_75t_L g2603 ( 
.A(n_2004),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2110),
.B(n_2119),
.Y(n_2604)
);

O2A1O1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_1631),
.A2(n_2041),
.B(n_2043),
.C(n_2016),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2119),
.A2(n_2121),
.B1(n_2137),
.B2(n_2129),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2121),
.B(n_2250),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_1821),
.A2(n_2041),
.B(n_2016),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2129),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2137),
.B(n_2141),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2141),
.B(n_2144),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2012),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2004),
.B(n_2095),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_1688),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_1871),
.B(n_1788),
.Y(n_2615)
);

AOI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_2041),
.A2(n_2057),
.B(n_2043),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2012),
.Y(n_2617)
);

AO32x1_ASAP7_75t_L g2618 ( 
.A1(n_2144),
.A2(n_2250),
.A3(n_2249),
.B1(n_2238),
.B2(n_2237),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2146),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2146),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_1991),
.A2(n_2035),
.B1(n_2101),
.B2(n_2243),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2095),
.B(n_2158),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_SL g2623 ( 
.A(n_1991),
.B(n_2035),
.Y(n_2623)
);

O2A1O1Ixp33_ASAP7_75t_L g2624 ( 
.A1(n_2043),
.A2(n_2060),
.B(n_2168),
.C(n_2122),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2147),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2149),
.Y(n_2626)
);

O2A1O1Ixp33_ASAP7_75t_L g2627 ( 
.A1(n_2057),
.A2(n_2060),
.B(n_2132),
.C(n_2122),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2149),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2154),
.B(n_2170),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2034),
.Y(n_2630)
);

OAI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2101),
.A2(n_2243),
.B1(n_2057),
.B2(n_2168),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2034),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2154),
.A2(n_2249),
.B1(n_2238),
.B2(n_2237),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_1871),
.B(n_1788),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2173),
.B(n_2183),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2034),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2073),
.A2(n_2132),
.B1(n_2168),
.B2(n_2101),
.Y(n_2637)
);

O2A1O1Ixp5_ASAP7_75t_L g2638 ( 
.A1(n_1885),
.A2(n_1886),
.B(n_2182),
.C(n_2162),
.Y(n_2638)
);

OAI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2173),
.A2(n_2207),
.B1(n_2198),
.B2(n_2234),
.Y(n_2639)
);

CKINVDCx11_ASAP7_75t_R g2640 ( 
.A(n_2095),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2183),
.A2(n_2184),
.B1(n_2187),
.B2(n_2234),
.Y(n_2641)
);

A2O1A1Ixp33_ASAP7_75t_L g2642 ( 
.A1(n_2001),
.A2(n_2200),
.B(n_2102),
.C(n_2096),
.Y(n_2642)
);

OAI321xp33_ASAP7_75t_L g2643 ( 
.A1(n_2198),
.A2(n_2233),
.A3(n_2227),
.B1(n_2221),
.B2(n_2220),
.C(n_2210),
.Y(n_2643)
);

NAND2x1_ASAP7_75t_L g2644 ( 
.A(n_1982),
.B(n_1788),
.Y(n_2644)
);

NAND2xp33_ASAP7_75t_L g2645 ( 
.A(n_1853),
.B(n_1888),
.Y(n_2645)
);

NOR2xp67_ASAP7_75t_L g2646 ( 
.A(n_1749),
.B(n_1757),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2202),
.A2(n_2208),
.B1(n_2233),
.B2(n_2227),
.Y(n_2647)
);

BUFx12f_ASAP7_75t_L g2648 ( 
.A(n_2158),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2001),
.A2(n_2200),
.B1(n_2102),
.B2(n_2096),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2081),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2202),
.B(n_2204),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2204),
.Y(n_2652)
);

INVx1_ASAP7_75t_SL g2653 ( 
.A(n_2156),
.Y(n_2653)
);

BUFx4f_ASAP7_75t_L g2654 ( 
.A(n_2158),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2206),
.B(n_2207),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2206),
.Y(n_2656)
);

OR2x2_ASAP7_75t_L g2657 ( 
.A(n_2208),
.B(n_2209),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2094),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2209),
.B(n_2210),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2220),
.B(n_2221),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2158),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_1970),
.B(n_2109),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2124),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2001),
.B(n_2072),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2126),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2244),
.A2(n_1590),
.B1(n_1603),
.B2(n_1611),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2134),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2157),
.Y(n_2668)
);

NOR2xp67_ASAP7_75t_L g2669 ( 
.A(n_1749),
.B(n_1757),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_1979),
.A2(n_1881),
.B1(n_1965),
.B2(n_1957),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2218),
.A2(n_2235),
.B(n_1810),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_1685),
.B(n_1686),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_1685),
.B(n_1686),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_1689),
.Y(n_2674)
);

O2A1O1Ixp33_ASAP7_75t_SL g2675 ( 
.A1(n_1773),
.A2(n_2244),
.B(n_1603),
.C(n_1611),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_1642),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_1642),
.Y(n_2677)
);

BUFx8_ASAP7_75t_L g2678 ( 
.A(n_2158),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_1689),
.Y(n_2679)
);

O2A1O1Ixp33_ASAP7_75t_SL g2680 ( 
.A1(n_2239),
.A2(n_2229),
.B(n_2193),
.C(n_2188),
.Y(n_2680)
);

OA22x2_ASAP7_75t_L g2681 ( 
.A1(n_1993),
.A2(n_2193),
.B1(n_2009),
.B2(n_2046),
.Y(n_2681)
);

NAND3xp33_ASAP7_75t_L g2682 ( 
.A(n_1853),
.B(n_1888),
.C(n_1848),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2072),
.Y(n_2683)
);

INVx5_ASAP7_75t_L g2684 ( 
.A(n_1853),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_1700),
.Y(n_2685)
);

O2A1O1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2046),
.A2(n_2188),
.B(n_2074),
.C(n_2159),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2074),
.A2(n_2159),
.B1(n_2138),
.B2(n_2105),
.Y(n_2687)
);

INVx3_ASAP7_75t_L g2688 ( 
.A(n_1853),
.Y(n_2688)
);

BUFx6f_ASAP7_75t_L g2689 ( 
.A(n_2072),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_L g2690 ( 
.A(n_1888),
.B(n_2093),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2093),
.Y(n_2691)
);

AOI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_2097),
.A2(n_2138),
.B(n_2105),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_1642),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_1700),
.B(n_1712),
.Y(n_2694)
);

AOI21xp5_ASAP7_75t_L g2695 ( 
.A1(n_1960),
.A2(n_1974),
.B(n_1969),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2093),
.Y(n_2696)
);

BUFx3_ASAP7_75t_L g2697 ( 
.A(n_2096),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2102),
.B(n_2200),
.Y(n_2698)
);

OAI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_1712),
.A2(n_1822),
.B1(n_1955),
.B2(n_1949),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_1714),
.A2(n_1837),
.B1(n_1965),
.B2(n_1971),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_1714),
.B(n_1715),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_1721),
.B(n_1729),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_1643),
.Y(n_2703)
);

INVxp67_ASAP7_75t_L g2704 ( 
.A(n_1721),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_1729),
.B(n_1736),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_SL g2706 ( 
.A(n_1662),
.B(n_1668),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_1799),
.A2(n_1939),
.B1(n_1858),
.B2(n_1854),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_1736),
.A2(n_1864),
.B1(n_1977),
.B2(n_1973),
.Y(n_2708)
);

CKINVDCx20_ASAP7_75t_R g2709 ( 
.A(n_1738),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_1738),
.B(n_1739),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_1739),
.A2(n_1872),
.B1(n_1977),
.B2(n_1973),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_1743),
.B(n_1971),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_1743),
.B(n_1967),
.Y(n_2713)
);

A2O1A1Ixp33_ASAP7_75t_L g2714 ( 
.A1(n_1747),
.A2(n_1854),
.B(n_1949),
.C(n_1946),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_1747),
.B(n_1967),
.Y(n_2715)
);

NOR3xp33_ASAP7_75t_L g2716 ( 
.A(n_1748),
.B(n_1842),
.C(n_1944),
.Y(n_2716)
);

BUFx6f_ASAP7_75t_L g2717 ( 
.A(n_1682),
.Y(n_2717)
);

NOR3xp33_ASAP7_75t_L g2718 ( 
.A(n_1748),
.B(n_1872),
.C(n_1944),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_1758),
.A2(n_1864),
.B(n_1940),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_1758),
.B(n_1877),
.Y(n_2720)
);

INVx4_ASAP7_75t_L g2721 ( 
.A(n_1713),
.Y(n_2721)
);

NOR3xp33_ASAP7_75t_L g2722 ( 
.A(n_1761),
.B(n_1877),
.C(n_1957),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_1761),
.B(n_1861),
.Y(n_2723)
);

O2A1O1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_1779),
.A2(n_1861),
.B(n_1955),
.C(n_1926),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_1779),
.B(n_1946),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_1780),
.A2(n_1829),
.B(n_1940),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_1725),
.Y(n_2727)
);

A2O1A1Ixp33_ASAP7_75t_L g2728 ( 
.A1(n_1780),
.A2(n_1829),
.B(n_1937),
.C(n_1899),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_1792),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_1792),
.B(n_1881),
.Y(n_2730)
);

A2O1A1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_1794),
.A2(n_1937),
.B(n_1910),
.C(n_1899),
.Y(n_2731)
);

INVx3_ASAP7_75t_L g2732 ( 
.A(n_1760),
.Y(n_2732)
);

OAI21xp33_ASAP7_75t_L g2733 ( 
.A1(n_1794),
.A2(n_1822),
.B(n_1896),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_1816),
.B(n_1926),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_1816),
.A2(n_1837),
.B(n_1917),
.C(n_1894),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_1819),
.Y(n_2736)
);

AND2x2_ASAP7_75t_SL g2737 ( 
.A(n_1839),
.B(n_1890),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_1762),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_1762),
.Y(n_2739)
);

O2A1O1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_1839),
.A2(n_1890),
.B(n_1896),
.C(n_1894),
.Y(n_2740)
);

OAI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_1842),
.A2(n_1887),
.B(n_1910),
.Y(n_2741)
);

A2O1A1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_1893),
.A2(n_1917),
.B(n_1928),
.C(n_1762),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_1782),
.Y(n_2743)
);

AOI21x1_ASAP7_75t_L g2744 ( 
.A1(n_1797),
.A2(n_1813),
.B(n_1809),
.Y(n_2744)
);

O2A1O1Ixp33_ASAP7_75t_L g2745 ( 
.A1(n_1820),
.A2(n_2211),
.B(n_1961),
.C(n_2140),
.Y(n_2745)
);

AOI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_1730),
.A2(n_1087),
.B1(n_1394),
.B2(n_1466),
.Y(n_2746)
);

NOR2xp67_ASAP7_75t_L g2747 ( 
.A(n_1750),
.B(n_1874),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_1927),
.B(n_1605),
.Y(n_2750)
);

A2O1A1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2042),
.A2(n_1490),
.B(n_1466),
.C(n_1374),
.Y(n_2751)
);

AOI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2176),
.A2(n_1087),
.B1(n_1480),
.B2(n_1545),
.C(n_1486),
.Y(n_2752)
);

OAI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_1644),
.Y(n_2754)
);

O2A1O1Ixp33_ASAP7_75t_L g2755 ( 
.A1(n_2100),
.A2(n_1486),
.B(n_1545),
.C(n_1480),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_1616),
.Y(n_2756)
);

AOI33xp33_ASAP7_75t_L g2757 ( 
.A1(n_1999),
.A2(n_2167),
.A3(n_2042),
.B1(n_2171),
.B2(n_2044),
.B3(n_2018),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_1661),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_1730),
.A2(n_1087),
.B1(n_1394),
.B2(n_1466),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2766)
);

OAI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2768)
);

AOI21x1_ASAP7_75t_L g2769 ( 
.A1(n_1593),
.A2(n_2143),
.B(n_2023),
.Y(n_2769)
);

OAI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2106),
.Y(n_2771)
);

OR2x6_ASAP7_75t_L g2772 ( 
.A(n_1658),
.B(n_1786),
.Y(n_2772)
);

AOI33xp33_ASAP7_75t_L g2773 ( 
.A1(n_1999),
.A2(n_2167),
.A3(n_2042),
.B1(n_2171),
.B2(n_2044),
.B3(n_2018),
.Y(n_2773)
);

AOI21xp33_ASAP7_75t_L g2774 ( 
.A1(n_2176),
.A2(n_1490),
.B(n_1466),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_1730),
.A2(n_1376),
.B1(n_1553),
.B2(n_845),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2777)
);

A2O1A1Ixp33_ASAP7_75t_SL g2778 ( 
.A1(n_1600),
.A2(n_1480),
.B(n_1545),
.C(n_1486),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1644),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_1996),
.B(n_2002),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_2053),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_1644),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2042),
.A2(n_1490),
.B(n_1466),
.C(n_1374),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2785)
);

A2O1A1Ixp33_ASAP7_75t_L g2786 ( 
.A1(n_2042),
.A2(n_1490),
.B(n_1466),
.C(n_1374),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_1616),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2788)
);

NAND2x1p5_ASAP7_75t_L g2789 ( 
.A(n_1661),
.B(n_1786),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2790)
);

NAND2x1p5_ASAP7_75t_L g2791 ( 
.A(n_1661),
.B(n_1786),
.Y(n_2791)
);

OAI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2792)
);

O2A1O1Ixp33_ASAP7_75t_L g2793 ( 
.A1(n_2100),
.A2(n_1486),
.B(n_1545),
.C(n_1480),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_1644),
.Y(n_2794)
);

OAI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2797)
);

AOI21x1_ASAP7_75t_L g2798 ( 
.A1(n_1593),
.A2(n_2143),
.B(n_2023),
.Y(n_2798)
);

OAI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2799)
);

NAND2xp33_ASAP7_75t_L g2800 ( 
.A(n_1620),
.B(n_1480),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_1996),
.B(n_2002),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_1927),
.B(n_1605),
.Y(n_2802)
);

NAND3xp33_ASAP7_75t_SL g2803 ( 
.A(n_1600),
.B(n_1486),
.C(n_1480),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_1616),
.Y(n_2804)
);

OAI22x1_ASAP7_75t_L g2805 ( 
.A1(n_1678),
.A2(n_1763),
.B1(n_1102),
.B2(n_1999),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2807)
);

NOR3xp33_ASAP7_75t_L g2808 ( 
.A(n_2100),
.B(n_1490),
.C(n_1466),
.Y(n_2808)
);

CKINVDCx11_ASAP7_75t_R g2809 ( 
.A(n_2113),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2810)
);

INVxp67_ASAP7_75t_L g2811 ( 
.A(n_1808),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2815)
);

OR2x2_ASAP7_75t_L g2816 ( 
.A(n_1927),
.B(n_1605),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_1616),
.Y(n_2817)
);

HB1xp67_ASAP7_75t_L g2818 ( 
.A(n_1767),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_1730),
.A2(n_1087),
.B1(n_1394),
.B2(n_1466),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2053),
.Y(n_2821)
);

BUFx3_ASAP7_75t_L g2822 ( 
.A(n_2053),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2824)
);

O2A1O1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2100),
.A2(n_1486),
.B(n_1545),
.C(n_1480),
.Y(n_2825)
);

BUFx3_ASAP7_75t_L g2826 ( 
.A(n_2053),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_1976),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2830)
);

OAI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_1661),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2836)
);

AOI21x1_ASAP7_75t_L g2837 ( 
.A1(n_1593),
.A2(n_2143),
.B(n_2023),
.Y(n_2837)
);

INVx2_ASAP7_75t_SL g2838 ( 
.A(n_1788),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2840)
);

AND2x4_ASAP7_75t_L g2841 ( 
.A(n_1728),
.B(n_1731),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_1644),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_1720),
.A2(n_1380),
.B(n_1374),
.Y(n_2843)
);

OAI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_1644),
.Y(n_2845)
);

OA22x2_ASAP7_75t_L g2846 ( 
.A1(n_1996),
.A2(n_1102),
.B1(n_2037),
.B2(n_2002),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_1693),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2849)
);

HB1xp67_ASAP7_75t_L g2850 ( 
.A(n_1767),
.Y(n_2850)
);

INVx1_ASAP7_75t_SL g2851 ( 
.A(n_1976),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_1999),
.A2(n_1466),
.B1(n_1490),
.B2(n_2018),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_1600),
.B(n_1614),
.Y(n_2854)
);

AOI21x1_ASAP7_75t_L g2855 ( 
.A1(n_1593),
.A2(n_2143),
.B(n_2023),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2857)
);

OAI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_1999),
.A2(n_1490),
.B1(n_1466),
.B2(n_1380),
.Y(n_2858)
);

NOR2xp67_ASAP7_75t_L g2859 ( 
.A(n_1750),
.B(n_1874),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2100),
.A2(n_1486),
.B(n_1545),
.C(n_1480),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2106),
.Y(n_2862)
);

OAI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_1644),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_1644),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2868)
);

OAI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_1616),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2872)
);

A2O1A1Ixp33_ASAP7_75t_L g2873 ( 
.A1(n_2042),
.A2(n_1490),
.B(n_1466),
.C(n_1374),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2874)
);

OAI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_1999),
.A2(n_1490),
.B(n_1466),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2877)
);

O2A1O1Ixp33_ASAP7_75t_L g2878 ( 
.A1(n_2100),
.A2(n_1486),
.B(n_1545),
.C(n_1480),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_1693),
.Y(n_2879)
);

NOR3xp33_ASAP7_75t_L g2880 ( 
.A(n_2100),
.B(n_1490),
.C(n_1466),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_1996),
.B(n_2002),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2176),
.B(n_1466),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2883)
);

INVx4_ASAP7_75t_L g2884 ( 
.A(n_2684),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2295),
.B(n_2750),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2553),
.B(n_2281),
.Y(n_2886)
);

NAND2x1_ASAP7_75t_L g2887 ( 
.A(n_2286),
.B(n_2278),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2314),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2749),
.B(n_2788),
.Y(n_2889)
);

OAI21x1_ASAP7_75t_SL g2890 ( 
.A1(n_2770),
.A2(n_2799),
.B(n_2792),
.Y(n_2890)
);

INVxp67_ASAP7_75t_SL g2891 ( 
.A(n_2477),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_SL g2892 ( 
.A1(n_2770),
.A2(n_2799),
.B(n_2792),
.Y(n_2892)
);

OAI221xp5_ASAP7_75t_L g2893 ( 
.A1(n_2264),
.A2(n_2254),
.B1(n_2271),
.B2(n_2761),
.C(n_2746),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2260),
.A2(n_2760),
.B(n_2753),
.Y(n_2894)
);

OAI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2259),
.A2(n_2285),
.B(n_2256),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_SL g2896 ( 
.A1(n_2275),
.A2(n_2784),
.B(n_2751),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2295),
.B(n_2750),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2812),
.B(n_2823),
.Y(n_2898)
);

AOI21x1_ASAP7_75t_L g2899 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_2899)
);

OAI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2760),
.A2(n_2776),
.B(n_2767),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2802),
.B(n_2816),
.Y(n_2902)
);

NAND3xp33_ASAP7_75t_L g2903 ( 
.A(n_2757),
.B(n_2773),
.C(n_2767),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2802),
.B(n_2816),
.Y(n_2904)
);

OAI21xp33_ASAP7_75t_L g2905 ( 
.A1(n_2776),
.A2(n_2795),
.B(n_2785),
.Y(n_2905)
);

BUFx2_ASAP7_75t_L g2906 ( 
.A(n_2344),
.Y(n_2906)
);

NAND2x1_ASAP7_75t_L g2907 ( 
.A(n_2286),
.B(n_2278),
.Y(n_2907)
);

OAI21xp33_ASAP7_75t_L g2908 ( 
.A1(n_2785),
.A2(n_2815),
.B(n_2795),
.Y(n_2908)
);

AOI221x1_ASAP7_75t_L g2909 ( 
.A1(n_2815),
.A2(n_2832),
.B1(n_2848),
.B2(n_2840),
.C(n_2839),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2314),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2289),
.B(n_2315),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2832),
.A2(n_2840),
.B(n_2839),
.Y(n_2912)
);

NAND2x1p5_ASAP7_75t_L g2913 ( 
.A(n_2346),
.B(n_2453),
.Y(n_2913)
);

NAND3xp33_ASAP7_75t_L g2914 ( 
.A(n_2848),
.B(n_2853),
.C(n_2289),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2853),
.A2(n_2761),
.B1(n_2820),
.B2(n_2746),
.Y(n_2915)
);

AO21x1_ASAP7_75t_L g2916 ( 
.A1(n_2765),
.A2(n_2806),
.B(n_2777),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2858),
.A2(n_2860),
.B(n_2810),
.Y(n_2917)
);

OAI22x1_ASAP7_75t_L g2918 ( 
.A1(n_2440),
.A2(n_2820),
.B1(n_2405),
.B2(n_2443),
.Y(n_2918)
);

INVx1_ASAP7_75t_SL g2919 ( 
.A(n_2405),
.Y(n_2919)
);

HB1xp67_ASAP7_75t_L g2920 ( 
.A(n_2527),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2824),
.B(n_2827),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2868),
.A2(n_2882),
.B(n_2876),
.Y(n_2922)
);

A2O1A1Ixp33_ASAP7_75t_L g2923 ( 
.A1(n_2313),
.A2(n_2273),
.B(n_2252),
.C(n_2288),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2500),
.B(n_2501),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2340),
.Y(n_2925)
);

INVx2_ASAP7_75t_SL g2926 ( 
.A(n_2514),
.Y(n_2926)
);

OAI222xp33_ASAP7_75t_L g2927 ( 
.A1(n_2438),
.A2(n_2355),
.B1(n_2266),
.B2(n_2440),
.C1(n_2846),
.C2(n_2775),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2786),
.A2(n_2873),
.B(n_2843),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2834),
.A2(n_2852),
.B(n_2849),
.Y(n_2929)
);

AO32x1_ASAP7_75t_L g2930 ( 
.A1(n_2355),
.A2(n_2302),
.A3(n_2639),
.B1(n_2647),
.B2(n_2721),
.Y(n_2930)
);

AOI21x1_ASAP7_75t_SL g2931 ( 
.A1(n_2255),
.A2(n_2748),
.B(n_2251),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2831),
.A2(n_2863),
.B(n_2844),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2378),
.B(n_2478),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_2344),
.Y(n_2934)
);

OAI21xp33_ASAP7_75t_L g2935 ( 
.A1(n_2854),
.A2(n_2844),
.B(n_2831),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2805),
.A2(n_2284),
.B1(n_2315),
.B2(n_2438),
.Y(n_2936)
);

OAI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2552),
.A2(n_2299),
.B(n_2616),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2863),
.A2(n_2875),
.B(n_2869),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2335),
.B(n_2350),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_2346),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2869),
.A2(n_2875),
.B(n_2774),
.Y(n_2941)
);

CKINVDCx20_ASAP7_75t_R g2942 ( 
.A(n_2809),
.Y(n_2942)
);

OAI21x1_ASAP7_75t_L g2943 ( 
.A1(n_2389),
.A2(n_2549),
.B(n_2547),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2258),
.A2(n_2267),
.B(n_2747),
.Y(n_2944)
);

NAND2x1p5_ASAP7_75t_L g2945 ( 
.A(n_2346),
.B(n_2453),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2752),
.A2(n_2300),
.B(n_2808),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2335),
.B(n_2350),
.Y(n_2947)
);

INVx1_ASAP7_75t_SL g2948 ( 
.A(n_2443),
.Y(n_2948)
);

OAI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2880),
.A2(n_2283),
.B(n_2296),
.Y(n_2949)
);

INVx3_ASAP7_75t_L g2950 ( 
.A(n_2274),
.Y(n_2950)
);

OAI21xp33_ASAP7_75t_SL g2951 ( 
.A1(n_2747),
.A2(n_2859),
.B(n_2394),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2859),
.A2(n_2360),
.B(n_2351),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2447),
.B(n_2456),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2579),
.Y(n_2954)
);

AOI21xp33_ASAP7_75t_L g2955 ( 
.A1(n_2294),
.A2(n_2805),
.B(n_2284),
.Y(n_2955)
);

AOI221xp5_ASAP7_75t_SL g2956 ( 
.A1(n_2755),
.A2(n_2825),
.B1(n_2878),
.B2(n_2861),
.C(n_2793),
.Y(n_2956)
);

A2O1A1Ixp33_ASAP7_75t_L g2957 ( 
.A1(n_2313),
.A2(n_2394),
.B(n_2323),
.C(n_2320),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_SL g2958 ( 
.A(n_2453),
.B(n_2504),
.Y(n_2958)
);

OR2x2_ASAP7_75t_L g2959 ( 
.A(n_2468),
.B(n_2529),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2340),
.Y(n_2960)
);

AOI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_2961)
);

NOR2x1_ASAP7_75t_SL g2962 ( 
.A(n_2486),
.B(n_2513),
.Y(n_2962)
);

OA21x2_ASAP7_75t_L g2963 ( 
.A1(n_2436),
.A2(n_2373),
.B(n_2638),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2425),
.A2(n_2505),
.B(n_2608),
.Y(n_2964)
);

OAI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2302),
.A2(n_2283),
.B1(n_2316),
.B2(n_2329),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2364),
.A2(n_2349),
.B(n_2778),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2484),
.B(n_2451),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_2579),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2312),
.A2(n_2328),
.B(n_2388),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2447),
.B(n_2456),
.Y(n_2970)
);

OAI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2294),
.A2(n_2297),
.B(n_2292),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2410),
.B(n_2265),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2297),
.B(n_2306),
.Y(n_2973)
);

AOI221x1_ASAP7_75t_L g2974 ( 
.A1(n_2803),
.A2(n_2463),
.B1(n_2329),
.B2(n_2306),
.C(n_2331),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2348),
.B(n_2358),
.Y(n_2975)
);

NOR3xp33_ASAP7_75t_L g2976 ( 
.A(n_2800),
.B(n_2303),
.C(n_2301),
.Y(n_2976)
);

OAI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2762),
.A2(n_2763),
.B1(n_2766),
.B2(n_2764),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2467),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2463),
.A2(n_2411),
.B(n_2338),
.C(n_2430),
.Y(n_2979)
);

INVx3_ASAP7_75t_L g2980 ( 
.A(n_2274),
.Y(n_2980)
);

INVx2_ASAP7_75t_SL g2981 ( 
.A(n_2514),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2348),
.Y(n_2982)
);

AO31x2_ASAP7_75t_L g2983 ( 
.A1(n_2471),
.A2(n_2373),
.A3(n_2647),
.B(n_2639),
.Y(n_2983)
);

OAI22x1_ASAP7_75t_L g2984 ( 
.A1(n_2437),
.A2(n_2262),
.B1(n_2403),
.B2(n_2837),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_L g2985 ( 
.A(n_2417),
.B(n_2343),
.C(n_2311),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2486),
.B(n_2397),
.Y(n_2986)
);

INVx5_ASAP7_75t_L g2987 ( 
.A(n_2772),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2358),
.B(n_2367),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2367),
.B(n_2370),
.Y(n_2989)
);

AO21x1_ASAP7_75t_L g2990 ( 
.A1(n_2426),
.A2(n_2324),
.B(n_2303),
.Y(n_2990)
);

OAI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2417),
.A2(n_2301),
.B(n_2343),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2370),
.B(n_2374),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2374),
.B(n_2377),
.Y(n_2993)
);

AO21x1_ASAP7_75t_L g2994 ( 
.A1(n_2426),
.A2(n_2855),
.B(n_2309),
.Y(n_2994)
);

OR2x6_ASAP7_75t_L g2995 ( 
.A(n_2479),
.B(n_2513),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2768),
.B(n_2782),
.Y(n_2996)
);

AO21x1_ASAP7_75t_L g2997 ( 
.A1(n_2436),
.A2(n_2489),
.B(n_2361),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2483),
.B(n_2263),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_SL g2999 ( 
.A1(n_2325),
.A2(n_2624),
.B(n_2605),
.Y(n_2999)
);

OAI21x1_ASAP7_75t_SL g3000 ( 
.A1(n_2627),
.A2(n_2567),
.B(n_2558),
.Y(n_3000)
);

BUFx6f_ASAP7_75t_L g3001 ( 
.A(n_2504),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2504),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2452),
.A2(n_2450),
.B(n_2446),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2754),
.B(n_2779),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2779),
.B(n_2783),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2783),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2410),
.B(n_2265),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2883),
.B(n_2790),
.Y(n_3008)
);

AO21x1_ASAP7_75t_L g3009 ( 
.A1(n_2356),
.A2(n_2379),
.B(n_2476),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2794),
.B(n_2842),
.Y(n_3010)
);

AND2x4_ASAP7_75t_L g3011 ( 
.A(n_2553),
.B(n_2281),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2541),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2467),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2796),
.B(n_2797),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2645),
.A2(n_2623),
.B(n_2603),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2794),
.B(n_2842),
.Y(n_3016)
);

INVx3_ASAP7_75t_SL g3017 ( 
.A(n_2578),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_2548),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2631),
.A2(n_2637),
.B(n_2671),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2413),
.A2(n_2434),
.B(n_2362),
.Y(n_3020)
);

INVx2_ASAP7_75t_SL g3021 ( 
.A(n_2541),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2578),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2845),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2807),
.A2(n_2814),
.B(n_2813),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2413),
.A2(n_2434),
.B(n_2362),
.Y(n_3025)
);

A2O1A1Ixp33_ASAP7_75t_L g3026 ( 
.A1(n_2369),
.A2(n_2354),
.B(n_2455),
.C(n_2819),
.Y(n_3026)
);

AOI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2623),
.A2(n_2654),
.B(n_2603),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2845),
.B(n_2864),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2603),
.A2(n_2654),
.B(n_2382),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2371),
.B(n_2366),
.Y(n_3030)
);

OAI22x1_ASAP7_75t_L g3031 ( 
.A1(n_2572),
.A2(n_2653),
.B1(n_2472),
.B2(n_2525),
.Y(n_3031)
);

BUFx6f_ASAP7_75t_L g3032 ( 
.A(n_2578),
.Y(n_3032)
);

BUFx4f_ASAP7_75t_SL g3033 ( 
.A(n_2422),
.Y(n_3033)
);

BUFx6f_ASAP7_75t_L g3034 ( 
.A(n_2291),
.Y(n_3034)
);

AO21x1_ASAP7_75t_L g3035 ( 
.A1(n_2476),
.A2(n_2466),
.B(n_2475),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2291),
.Y(n_3036)
);

BUFx6f_ASAP7_75t_L g3037 ( 
.A(n_2291),
.Y(n_3037)
);

A2O1A1Ixp33_ASAP7_75t_L g3038 ( 
.A1(n_2829),
.A2(n_2833),
.B(n_2836),
.C(n_2830),
.Y(n_3038)
);

INVx1_ASAP7_75t_SL g3039 ( 
.A(n_2594),
.Y(n_3039)
);

BUFx3_ASAP7_75t_L g3040 ( 
.A(n_2424),
.Y(n_3040)
);

NOR2x1_ASAP7_75t_L g3041 ( 
.A(n_2581),
.B(n_2568),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2268),
.B(n_2290),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2856),
.B(n_2857),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2654),
.A2(n_2384),
.B(n_2376),
.Y(n_3044)
);

OAI21x1_ASAP7_75t_L g3045 ( 
.A1(n_2644),
.A2(n_2789),
.B(n_2287),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2865),
.B(n_2866),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_2468),
.B(n_2529),
.Y(n_3047)
);

AOI21x1_ASAP7_75t_SL g3048 ( 
.A1(n_2870),
.A2(n_2874),
.B(n_2872),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2548),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2497),
.Y(n_3050)
);

OAI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2877),
.A2(n_2261),
.B(n_2257),
.Y(n_3051)
);

CKINVDCx6p67_ASAP7_75t_R g3052 ( 
.A(n_2270),
.Y(n_3052)
);

OAI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2272),
.A2(n_2280),
.B(n_2277),
.Y(n_3053)
);

OAI21x1_ASAP7_75t_L g3054 ( 
.A1(n_2287),
.A2(n_2791),
.B(n_2789),
.Y(n_3054)
);

HB1xp67_ASAP7_75t_L g3055 ( 
.A(n_2818),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2864),
.Y(n_3056)
);

AO31x2_ASAP7_75t_L g3057 ( 
.A1(n_2742),
.A2(n_2592),
.A3(n_2721),
.B(n_2714),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2268),
.B(n_2290),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2461),
.A2(n_2522),
.B(n_2588),
.Y(n_3059)
);

AND2x2_ASAP7_75t_SL g3060 ( 
.A(n_2737),
.B(n_2538),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_SL g3061 ( 
.A(n_2263),
.B(n_2828),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2381),
.B(n_2490),
.Y(n_3062)
);

AO31x2_ASAP7_75t_L g3063 ( 
.A1(n_2592),
.A2(n_2721),
.A3(n_2731),
.B(n_2728),
.Y(n_3063)
);

INVxp67_ASAP7_75t_SL g3064 ( 
.A(n_2732),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2850),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2494),
.B(n_2298),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2319),
.B(n_2321),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2393),
.B(n_2409),
.Y(n_3068)
);

OAI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2322),
.A2(n_2327),
.B(n_2326),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2333),
.A2(n_2339),
.B(n_2334),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2867),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_SL g3072 ( 
.A1(n_2510),
.A2(n_2524),
.B(n_2517),
.Y(n_3072)
);

OAI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2580),
.A2(n_2511),
.B(n_2571),
.Y(n_3073)
);

AOI21x1_ASAP7_75t_L g3074 ( 
.A1(n_2433),
.A2(n_2442),
.B(n_2613),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2867),
.Y(n_3075)
);

AO31x2_ASAP7_75t_L g3076 ( 
.A1(n_2721),
.A2(n_2735),
.A3(n_2707),
.B(n_2308),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2341),
.B(n_2342),
.Y(n_3077)
);

AO31x2_ASAP7_75t_L g3078 ( 
.A1(n_2707),
.A2(n_2308),
.A3(n_2399),
.B(n_2365),
.Y(n_3078)
);

OAI21x1_ASAP7_75t_SL g3079 ( 
.A1(n_2445),
.A2(n_2492),
.B(n_2564),
.Y(n_3079)
);

AO31x2_ASAP7_75t_L g3080 ( 
.A1(n_2308),
.A2(n_2365),
.A3(n_2402),
.B(n_2399),
.Y(n_3080)
);

NAND2x1p5_ASAP7_75t_L g3081 ( 
.A(n_2526),
.B(n_2535),
.Y(n_3081)
);

AOI21x1_ASAP7_75t_L g3082 ( 
.A1(n_2433),
.A2(n_2442),
.B(n_2622),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2400),
.B(n_2408),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2404),
.Y(n_3084)
);

NAND2x1p5_ASAP7_75t_L g3085 ( 
.A(n_2526),
.B(n_2535),
.Y(n_3085)
);

OAI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2345),
.A2(n_2353),
.B(n_2352),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2427),
.B(n_2828),
.Y(n_3087)
);

OAI21xp5_ASAP7_75t_L g3088 ( 
.A1(n_2398),
.A2(n_2330),
.B(n_2279),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2439),
.B(n_2431),
.Y(n_3089)
);

CKINVDCx6p67_ASAP7_75t_R g3090 ( 
.A(n_2270),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2497),
.Y(n_3091)
);

AOI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_2438),
.A2(n_2709),
.B1(n_2846),
.B2(n_2396),
.Y(n_3092)
);

O2A1O1Ixp5_ASAP7_75t_L g3093 ( 
.A1(n_2459),
.A2(n_2502),
.B(n_2595),
.C(n_2576),
.Y(n_3093)
);

AOI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2692),
.A2(n_2698),
.B(n_2669),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2499),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2546),
.A2(n_2543),
.B(n_2538),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2546),
.A2(n_2543),
.B(n_2479),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2706),
.A2(n_2680),
.B(n_2675),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2706),
.A2(n_2554),
.B(n_2561),
.Y(n_3099)
);

AND3x2_ASAP7_75t_L g3100 ( 
.A(n_2562),
.B(n_2590),
.C(n_2372),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2684),
.A2(n_2737),
.B(n_2565),
.Y(n_3101)
);

AOI221xp5_ASAP7_75t_L g3102 ( 
.A1(n_2276),
.A2(n_2811),
.B1(n_2419),
.B2(n_2421),
.C(n_2457),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2393),
.B(n_2409),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2684),
.A2(n_2737),
.B(n_2432),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2780),
.B(n_2801),
.Y(n_3105)
);

NOR2xp67_ASAP7_75t_L g3106 ( 
.A(n_2643),
.B(n_2485),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2684),
.A2(n_2586),
.B(n_2507),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2415),
.B(n_2416),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2383),
.A2(n_2458),
.B(n_2332),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2684),
.A2(n_2586),
.B(n_2506),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2502),
.A2(n_2545),
.B(n_2401),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2415),
.B(n_2416),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2499),
.Y(n_3113)
);

NAND2x1_ASAP7_75t_L g3114 ( 
.A(n_2688),
.B(n_2359),
.Y(n_3114)
);

OA21x2_ASAP7_75t_L g3115 ( 
.A1(n_2733),
.A2(n_2726),
.B(n_2719),
.Y(n_3115)
);

NAND2x1p5_ASAP7_75t_L g3116 ( 
.A(n_2526),
.B(n_2535),
.Y(n_3116)
);

BUFx4_ASAP7_75t_SL g3117 ( 
.A(n_2771),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2418),
.B(n_2454),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2359),
.A2(n_2470),
.B(n_2391),
.Y(n_3119)
);

AO31x2_ASAP7_75t_L g3120 ( 
.A1(n_2365),
.A2(n_2399),
.A3(n_2414),
.B(n_2402),
.Y(n_3120)
);

NAND2x1_ASAP7_75t_L g3121 ( 
.A(n_2688),
.B(n_2359),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2291),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2621),
.A2(n_2642),
.B(n_2559),
.Y(n_3123)
);

OAI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2536),
.A2(n_2537),
.B(n_2512),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2291),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2499),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2418),
.B(n_2454),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2460),
.B(n_2487),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2460),
.B(n_2487),
.Y(n_3129)
);

AND3x2_ASAP7_75t_L g3130 ( 
.A(n_2569),
.B(n_2575),
.C(n_2551),
.Y(n_3130)
);

OAI21x1_ASAP7_75t_L g3131 ( 
.A1(n_2391),
.A2(n_2496),
.B(n_2470),
.Y(n_3131)
);

OAI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_2851),
.A2(n_2412),
.B1(n_2846),
.B2(n_2525),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_2307),
.A2(n_2653),
.B1(n_2572),
.B2(n_2429),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2583),
.B(n_2598),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_2496),
.A2(n_2509),
.B(n_2503),
.Y(n_3135)
);

OAI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2493),
.A2(n_2515),
.B(n_2444),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2583),
.B(n_2598),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2609),
.B(n_2619),
.Y(n_3138)
);

A2O1A1Ixp33_ASAP7_75t_L g3139 ( 
.A1(n_2305),
.A2(n_2556),
.B(n_2533),
.C(n_2508),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2851),
.A2(n_2472),
.B1(n_2406),
.B2(n_2582),
.Y(n_3140)
);

OAI21x1_ASAP7_75t_L g3141 ( 
.A1(n_2496),
.A2(n_2509),
.B(n_2503),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_SL g3142 ( 
.A(n_2395),
.B(n_2528),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2759),
.Y(n_3143)
);

O2A1O1Ixp5_ASAP7_75t_L g3144 ( 
.A1(n_2576),
.A2(n_2595),
.B(n_2491),
.C(n_2530),
.Y(n_3144)
);

OAI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2485),
.A2(n_2581),
.B(n_2696),
.Y(n_3145)
);

INVxp67_ASAP7_75t_L g3146 ( 
.A(n_2386),
.Y(n_3146)
);

HB1xp67_ASAP7_75t_L g3147 ( 
.A(n_2407),
.Y(n_3147)
);

OAI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2532),
.A2(n_2686),
.B(n_2615),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2609),
.Y(n_3149)
);

CKINVDCx20_ASAP7_75t_R g3150 ( 
.A(n_2435),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2518),
.Y(n_3151)
);

AO221x2_ASAP7_75t_L g3152 ( 
.A1(n_2318),
.A2(n_2582),
.B1(n_2307),
.B2(n_2699),
.C(n_2682),
.Y(n_3152)
);

A2O1A1Ixp33_ASAP7_75t_L g3153 ( 
.A1(n_2305),
.A2(n_2596),
.B(n_2682),
.C(n_2304),
.Y(n_3153)
);

OAI21xp33_ASAP7_75t_L g3154 ( 
.A1(n_2307),
.A2(n_2862),
.B(n_2771),
.Y(n_3154)
);

OAI21x1_ASAP7_75t_L g3155 ( 
.A1(n_2847),
.A2(n_2879),
.B(n_2688),
.Y(n_3155)
);

NOR2x1_ASAP7_75t_L g3156 ( 
.A(n_2697),
.B(n_2576),
.Y(n_3156)
);

OAI21x1_ASAP7_75t_L g3157 ( 
.A1(n_2879),
.A2(n_2688),
.B(n_2595),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2620),
.B(n_2625),
.Y(n_3158)
);

OAI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2599),
.A2(n_2634),
.B(n_2666),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2518),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2666),
.A2(n_2687),
.B(n_2591),
.Y(n_3161)
);

AND2x4_ASAP7_75t_SL g3162 ( 
.A(n_2772),
.B(n_2269),
.Y(n_3162)
);

AO31x2_ASAP7_75t_L g3163 ( 
.A1(n_2402),
.A2(n_2414),
.A3(n_2756),
.B(n_2449),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2687),
.A2(n_2838),
.B(n_2591),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2518),
.Y(n_3165)
);

NOR2x1_ASAP7_75t_SL g3166 ( 
.A(n_2772),
.B(n_2304),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2626),
.B(n_2628),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2628),
.B(n_2652),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_2780),
.B(n_2801),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_2652),
.Y(n_3170)
);

AND3x2_ASAP7_75t_L g3171 ( 
.A(n_2357),
.B(n_2385),
.C(n_2363),
.Y(n_3171)
);

A2O1A1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_2448),
.A2(n_2462),
.B(n_2482),
.C(n_2474),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2656),
.B(n_2481),
.Y(n_3173)
);

OAI21xp5_ASAP7_75t_SL g3174 ( 
.A1(n_2441),
.A2(n_2465),
.B(n_2420),
.Y(n_3174)
);

AOI21x1_ASAP7_75t_L g3175 ( 
.A1(n_2646),
.A2(n_2649),
.B(n_2614),
.Y(n_3175)
);

AND2x6_ASAP7_75t_L g3176 ( 
.A(n_2448),
.B(n_2462),
.Y(n_3176)
);

AOI21xp33_ASAP7_75t_L g3177 ( 
.A1(n_2681),
.A2(n_2740),
.B(n_2724),
.Y(n_3177)
);

AO31x2_ASAP7_75t_L g3178 ( 
.A1(n_2414),
.A2(n_2756),
.A3(n_2787),
.B(n_2449),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2881),
.B(n_2387),
.Y(n_3179)
);

OR2x6_ASAP7_75t_L g3180 ( 
.A(n_2448),
.B(n_2462),
.Y(n_3180)
);

A2O1A1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_2474),
.A2(n_2482),
.B(n_2781),
.C(n_2826),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2862),
.B(n_2392),
.Y(n_3182)
);

OAI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2838),
.A2(n_2690),
.B(n_2704),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_2395),
.B(n_2495),
.Y(n_3184)
);

AO31x2_ASAP7_75t_L g3185 ( 
.A1(n_2449),
.A2(n_2756),
.A3(n_2804),
.B(n_2871),
.Y(n_3185)
);

OAI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2716),
.A2(n_2722),
.B(n_2718),
.Y(n_3186)
);

OAI22x1_ASAP7_75t_L g3187 ( 
.A1(n_2269),
.A2(n_2429),
.B1(n_2881),
.B2(n_2253),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2481),
.B(n_2516),
.Y(n_3188)
);

OAI22x1_ASAP7_75t_L g3189 ( 
.A1(n_2269),
.A2(n_2429),
.B1(n_2310),
.B2(n_2841),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2516),
.B(n_2539),
.Y(n_3190)
);

O2A1O1Ixp5_ASAP7_75t_L g3191 ( 
.A1(n_2540),
.A2(n_2542),
.B(n_2664),
.C(n_2544),
.Y(n_3191)
);

OAI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2719),
.A2(n_2741),
.B(n_2726),
.Y(n_3192)
);

AND2x4_ASAP7_75t_L g3193 ( 
.A(n_2474),
.B(n_2482),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_2640),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2733),
.A2(n_2681),
.B(n_2695),
.Y(n_3195)
);

AOI21x1_ASAP7_75t_SL g3196 ( 
.A1(n_2480),
.A2(n_2318),
.B(n_2337),
.Y(n_3196)
);

AND2x4_ASAP7_75t_L g3197 ( 
.A(n_2781),
.B(n_2821),
.Y(n_3197)
);

OAI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_2700),
.A2(n_2681),
.B(n_2557),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2550),
.Y(n_3199)
);

INVxp67_ASAP7_75t_L g3200 ( 
.A(n_2560),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2587),
.B(n_2610),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2587),
.B(n_2610),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_2759),
.Y(n_3203)
);

OAI22x1_ASAP7_75t_L g3204 ( 
.A1(n_2253),
.A2(n_2310),
.B1(n_2841),
.B2(n_2336),
.Y(n_3204)
);

HB1xp67_ASAP7_75t_L g3205 ( 
.A(n_2607),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2423),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_2253),
.B(n_2310),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2712),
.B(n_2725),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2310),
.B(n_2336),
.Y(n_3209)
);

NAND2x1p5_ASAP7_75t_L g3210 ( 
.A(n_2821),
.B(n_2822),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2730),
.B(n_2734),
.Y(n_3211)
);

BUFx12f_ASAP7_75t_L g3212 ( 
.A(n_2495),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2694),
.B(n_2702),
.Y(n_3213)
);

INVx2_ASAP7_75t_SL g3214 ( 
.A(n_2336),
.Y(n_3214)
);

OAI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2700),
.A2(n_2745),
.B(n_2670),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2694),
.B(n_2702),
.Y(n_3216)
);

HB1xp67_ASAP7_75t_L g3217 ( 
.A(n_2607),
.Y(n_3217)
);

HB1xp67_ASAP7_75t_L g3218 ( 
.A(n_2657),
.Y(n_3218)
);

A2O1A1Ixp33_ASAP7_75t_L g3219 ( 
.A1(n_2821),
.A2(n_2822),
.B(n_2826),
.C(n_2835),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2480),
.A2(n_2826),
.B1(n_2822),
.B2(n_2375),
.Y(n_3220)
);

OAI21x1_ASAP7_75t_L g3221 ( 
.A1(n_2732),
.A2(n_2738),
.B(n_2736),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2336),
.B(n_2347),
.Y(n_3222)
);

HAxp5_ASAP7_75t_L g3223 ( 
.A(n_2337),
.B(n_2390),
.CON(n_3223),
.SN(n_3223)
);

NAND2x1p5_ASAP7_75t_L g3224 ( 
.A(n_2380),
.B(n_2759),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_SL g3225 ( 
.A1(n_2759),
.A2(n_2835),
.B(n_2772),
.Y(n_3225)
);

NAND3xp33_ASAP7_75t_L g3226 ( 
.A(n_2606),
.B(n_2641),
.C(n_2633),
.Y(n_3226)
);

OAI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_2347),
.A2(n_2841),
.B1(n_2368),
.B2(n_2375),
.Y(n_3227)
);

OAI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2674),
.A2(n_2679),
.B(n_2685),
.Y(n_3228)
);

OAI21x1_ASAP7_75t_L g3229 ( 
.A1(n_2732),
.A2(n_2738),
.B(n_2736),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_2347),
.B(n_2368),
.Y(n_3230)
);

OAI21x1_ASAP7_75t_SL g3231 ( 
.A1(n_2563),
.A2(n_2600),
.B(n_2584),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2566),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2705),
.B(n_2683),
.Y(n_3233)
);

OAI21x1_ASAP7_75t_L g3234 ( 
.A1(n_2732),
.A2(n_2729),
.B(n_2674),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2423),
.Y(n_3235)
);

OAI21x1_ASAP7_75t_L g3236 ( 
.A1(n_2679),
.A2(n_2729),
.B(n_2685),
.Y(n_3236)
);

AO21x1_ASAP7_75t_L g3237 ( 
.A1(n_2570),
.A2(n_2611),
.B(n_2660),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_2317),
.Y(n_3238)
);

BUFx4f_ASAP7_75t_L g3239 ( 
.A(n_2835),
.Y(n_3239)
);

NAND2x1p5_ASAP7_75t_L g3240 ( 
.A(n_2380),
.B(n_2835),
.Y(n_3240)
);

OAI21x1_ASAP7_75t_L g3241 ( 
.A1(n_2672),
.A2(n_2710),
.B(n_2701),
.Y(n_3241)
);

AND3x4_ASAP7_75t_L g3242 ( 
.A(n_2368),
.B(n_2375),
.C(n_2841),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_2566),
.Y(n_3243)
);

A2O1A1Ixp33_ASAP7_75t_L g3244 ( 
.A1(n_2835),
.A2(n_2375),
.B(n_2758),
.C(n_2523),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2423),
.Y(n_3245)
);

AOI21x1_ASAP7_75t_L g3246 ( 
.A1(n_2573),
.A2(n_2651),
.B(n_2655),
.Y(n_3246)
);

OAI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_2708),
.A2(n_2711),
.B(n_2604),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2566),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2661),
.A2(n_2758),
.B(n_2618),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2612),
.Y(n_3250)
);

OAI22x1_ASAP7_75t_L g3251 ( 
.A1(n_2758),
.A2(n_2667),
.B1(n_2663),
.B2(n_2665),
.Y(n_3251)
);

OA21x2_ASAP7_75t_L g3252 ( 
.A1(n_2673),
.A2(n_2723),
.B(n_2715),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2661),
.A2(n_2758),
.B(n_2618),
.Y(n_3253)
);

OAI21x1_ASAP7_75t_SL g3254 ( 
.A1(n_2574),
.A2(n_2635),
.B(n_2659),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2395),
.B(n_2422),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2663),
.B(n_2665),
.Y(n_3256)
);

OR2x6_ASAP7_75t_L g3257 ( 
.A(n_2597),
.B(n_2717),
.Y(n_3257)
);

OAI21x1_ASAP7_75t_L g3258 ( 
.A1(n_2713),
.A2(n_2720),
.B(n_2585),
.Y(n_3258)
);

BUFx2_ASAP7_75t_R g3259 ( 
.A(n_2662),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2612),
.Y(n_3260)
);

AOI21x1_ASAP7_75t_SL g3261 ( 
.A1(n_2390),
.A2(n_2555),
.B(n_2488),
.Y(n_3261)
);

OAI21x1_ASAP7_75t_L g3262 ( 
.A1(n_2577),
.A2(n_2589),
.B(n_2602),
.Y(n_3262)
);

OAI21x1_ASAP7_75t_L g3263 ( 
.A1(n_2593),
.A2(n_2629),
.B(n_2601),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2618),
.A2(n_2689),
.B(n_2691),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2612),
.Y(n_3265)
);

AO221x2_ASAP7_75t_L g3266 ( 
.A1(n_2435),
.A2(n_2488),
.B1(n_2555),
.B2(n_2597),
.C(n_2618),
.Y(n_3266)
);

INVx4_ASAP7_75t_L g3267 ( 
.A(n_2648),
.Y(n_3267)
);

NAND3xp33_ASAP7_75t_L g3268 ( 
.A(n_2435),
.B(n_2555),
.C(n_2488),
.Y(n_3268)
);

OAI22x1_ASAP7_75t_L g3269 ( 
.A1(n_2667),
.A2(n_2668),
.B1(n_2521),
.B2(n_2520),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_SL g3270 ( 
.A1(n_2469),
.A2(n_2519),
.B(n_2498),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2617),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2668),
.Y(n_3272)
);

AOI21xp33_ASAP7_75t_L g3273 ( 
.A1(n_2717),
.A2(n_2727),
.B(n_2691),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2618),
.Y(n_3274)
);

OA21x2_ASAP7_75t_L g3275 ( 
.A1(n_2617),
.A2(n_2658),
.B(n_2632),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2630),
.B(n_2658),
.Y(n_3276)
);

BUFx8_ASAP7_75t_L g3277 ( 
.A(n_2648),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2630),
.B(n_2632),
.Y(n_3278)
);

A2O1A1Ixp33_ASAP7_75t_L g3279 ( 
.A1(n_2469),
.A2(n_2519),
.B(n_2498),
.C(n_2534),
.Y(n_3279)
);

INVx4_ASAP7_75t_L g3280 ( 
.A(n_2691),
.Y(n_3280)
);

AO21x2_ASAP7_75t_L g3281 ( 
.A1(n_2636),
.A2(n_2650),
.B(n_2743),
.Y(n_3281)
);

AOI21x1_ASAP7_75t_L g3282 ( 
.A1(n_2650),
.A2(n_2739),
.B(n_2677),
.Y(n_3282)
);

OAI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_2464),
.A2(n_2473),
.B1(n_2534),
.B2(n_2519),
.Y(n_3283)
);

OAI21xp33_ASAP7_75t_L g3284 ( 
.A1(n_2498),
.A2(n_2534),
.B(n_2531),
.Y(n_3284)
);

BUFx3_ASAP7_75t_L g3285 ( 
.A(n_2424),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2676),
.B(n_2693),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_SL g3287 ( 
.A(n_2424),
.B(n_2428),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_SL g3288 ( 
.A(n_2519),
.B(n_2534),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2677),
.B(n_2703),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2787),
.Y(n_3290)
);

A2O1A1Ixp33_ASAP7_75t_L g3291 ( 
.A1(n_2531),
.A2(n_2804),
.B(n_2787),
.C(n_2817),
.Y(n_3291)
);

BUFx2_ASAP7_75t_SL g3292 ( 
.A(n_2424),
.Y(n_3292)
);

OAI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_2804),
.A2(n_2817),
.B(n_2428),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2717),
.B(n_2727),
.Y(n_3294)
);

AOI21x1_ASAP7_75t_SL g3295 ( 
.A1(n_2435),
.A2(n_2488),
.B(n_2555),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_2531),
.A2(n_2817),
.B(n_2727),
.C(n_2464),
.Y(n_3296)
);

OAI21x1_ASAP7_75t_L g3297 ( 
.A1(n_2678),
.A2(n_2424),
.B(n_2428),
.Y(n_3297)
);

AOI21x1_ASAP7_75t_L g3298 ( 
.A1(n_2678),
.A2(n_2424),
.B(n_2428),
.Y(n_3298)
);

INVx3_ASAP7_75t_SL g3299 ( 
.A(n_2424),
.Y(n_3299)
);

AND2x4_ASAP7_75t_L g3300 ( 
.A(n_2428),
.B(n_2678),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_2428),
.B(n_2678),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2428),
.A2(n_1380),
.B(n_1374),
.Y(n_3302)
);

BUFx2_ASAP7_75t_L g3303 ( 
.A(n_2473),
.Y(n_3303)
);

INVxp33_ASAP7_75t_SL g3304 ( 
.A(n_2317),
.Y(n_3304)
);

NAND2x1p5_ASAP7_75t_L g3305 ( 
.A(n_2346),
.B(n_2453),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_SL g3306 ( 
.A(n_2289),
.B(n_2259),
.Y(n_3306)
);

NOR2xp67_ASAP7_75t_L g3307 ( 
.A(n_2260),
.B(n_2299),
.Y(n_3307)
);

AOI21xp33_ASAP7_75t_L g3308 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2744),
.Y(n_3309)
);

AO31x2_ASAP7_75t_L g3310 ( 
.A1(n_2471),
.A2(n_1447),
.A3(n_2373),
.B(n_2805),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3312)
);

AOI21xp33_ASAP7_75t_L g3313 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2744),
.Y(n_3314)
);

AOI21xp5_ASAP7_75t_L g3315 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_SL g3316 ( 
.A1(n_2271),
.A2(n_1380),
.B(n_1374),
.Y(n_3316)
);

AOI21x1_ASAP7_75t_L g3317 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3319)
);

INVx3_ASAP7_75t_L g3320 ( 
.A(n_2293),
.Y(n_3320)
);

INVxp67_ASAP7_75t_L g3321 ( 
.A(n_2439),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2744),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_2744),
.Y(n_3323)
);

OAI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_2254),
.A2(n_2264),
.B1(n_2761),
.B2(n_2746),
.Y(n_3324)
);

BUFx5_ASAP7_75t_L g3325 ( 
.A(n_2578),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3326)
);

BUFx4f_ASAP7_75t_L g3327 ( 
.A(n_2291),
.Y(n_3327)
);

OAI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3329)
);

AO31x2_ASAP7_75t_L g3330 ( 
.A1(n_2471),
.A2(n_1447),
.A3(n_2373),
.B(n_2805),
.Y(n_3330)
);

AOI221xp5_ASAP7_75t_L g3331 ( 
.A1(n_2259),
.A2(n_2254),
.B1(n_2271),
.B2(n_2760),
.C(n_2753),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_2314),
.Y(n_3333)
);

AND2x2_ASAP7_75t_SL g3334 ( 
.A(n_2737),
.B(n_2346),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2314),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3336)
);

BUFx12f_ASAP7_75t_L g3337 ( 
.A(n_2809),
.Y(n_3337)
);

INVxp67_ASAP7_75t_L g3338 ( 
.A(n_2439),
.Y(n_3338)
);

OAI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2744),
.Y(n_3340)
);

A2O1A1Ixp33_ASAP7_75t_L g3341 ( 
.A1(n_2757),
.A2(n_2773),
.B(n_2254),
.C(n_2264),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_SL g3342 ( 
.A1(n_2264),
.A2(n_2254),
.B(n_2289),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2744),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3344)
);

NAND2x1p5_ASAP7_75t_L g3345 ( 
.A(n_2346),
.B(n_2453),
.Y(n_3345)
);

CKINVDCx20_ASAP7_75t_R g3346 ( 
.A(n_2809),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2314),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3348)
);

AO31x2_ASAP7_75t_L g3349 ( 
.A1(n_2471),
.A2(n_1447),
.A3(n_2373),
.B(n_2805),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_SL g3350 ( 
.A(n_2289),
.B(n_2259),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_2346),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2749),
.B(n_2788),
.Y(n_3353)
);

HB1xp67_ASAP7_75t_L g3354 ( 
.A(n_2527),
.Y(n_3354)
);

BUFx4f_ASAP7_75t_L g3355 ( 
.A(n_2291),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2314),
.Y(n_3356)
);

INVx4_ASAP7_75t_L g3357 ( 
.A(n_2684),
.Y(n_3357)
);

INVx1_ASAP7_75t_SL g3358 ( 
.A(n_2295),
.Y(n_3358)
);

AO21x1_ASAP7_75t_L g3359 ( 
.A1(n_2256),
.A2(n_2760),
.B(n_2753),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_SL g3360 ( 
.A1(n_2271),
.A2(n_1380),
.B(n_1374),
.Y(n_3360)
);

INVx3_ASAP7_75t_L g3361 ( 
.A(n_2293),
.Y(n_3361)
);

NAND2x1p5_ASAP7_75t_L g3362 ( 
.A(n_2346),
.B(n_2453),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2744),
.Y(n_3363)
);

AOI21x1_ASAP7_75t_L g3364 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_3364)
);

NOR2x1_ASAP7_75t_SL g3365 ( 
.A(n_2486),
.B(n_2513),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_2289),
.B(n_2259),
.Y(n_3366)
);

AO31x2_ASAP7_75t_L g3367 ( 
.A1(n_2471),
.A2(n_1447),
.A3(n_2373),
.B(n_2805),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_2346),
.B(n_2453),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_2744),
.Y(n_3369)
);

A2O1A1Ixp33_ASAP7_75t_L g3370 ( 
.A1(n_2757),
.A2(n_2773),
.B(n_2254),
.C(n_2264),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3371)
);

HB1xp67_ASAP7_75t_L g3372 ( 
.A(n_2527),
.Y(n_3372)
);

AOI21x1_ASAP7_75t_L g3373 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_3373)
);

AOI21x1_ASAP7_75t_L g3374 ( 
.A1(n_2282),
.A2(n_2798),
.B(n_2769),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3376)
);

NAND2xp33_ASAP7_75t_L g3377 ( 
.A(n_2285),
.B(n_1480),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2314),
.Y(n_3378)
);

BUFx3_ASAP7_75t_L g3379 ( 
.A(n_2579),
.Y(n_3379)
);

OAI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3382)
);

AOI21xp33_ASAP7_75t_L g3383 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2744),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_2527),
.Y(n_3385)
);

OAI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3387)
);

OAI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3388)
);

INVxp67_ASAP7_75t_SL g3389 ( 
.A(n_2477),
.Y(n_3389)
);

NAND3xp33_ASAP7_75t_L g3390 ( 
.A(n_2254),
.B(n_2264),
.C(n_2271),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3392)
);

OAI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_2254),
.A2(n_2264),
.B1(n_2761),
.B2(n_2746),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3395)
);

O2A1O1Ixp5_ASAP7_75t_L g3396 ( 
.A1(n_2256),
.A2(n_2285),
.B(n_2777),
.C(n_2765),
.Y(n_3396)
);

OR2x6_ASAP7_75t_L g3397 ( 
.A(n_2479),
.B(n_2513),
.Y(n_3397)
);

AOI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3398)
);

NAND3xp33_ASAP7_75t_L g3399 ( 
.A(n_2254),
.B(n_2264),
.C(n_2271),
.Y(n_3399)
);

INVx5_ASAP7_75t_L g3400 ( 
.A(n_2772),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3402)
);

AO21x1_ASAP7_75t_L g3403 ( 
.A1(n_2256),
.A2(n_2760),
.B(n_2753),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3404)
);

AO21x2_ASAP7_75t_L g3405 ( 
.A1(n_2426),
.A2(n_1447),
.B(n_2373),
.Y(n_3405)
);

OAI21x1_ASAP7_75t_SL g3406 ( 
.A1(n_2770),
.A2(n_2799),
.B(n_2792),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3407)
);

OAI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_2254),
.A2(n_2264),
.B1(n_2761),
.B2(n_2746),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_2744),
.Y(n_3409)
);

INVx3_ASAP7_75t_L g3410 ( 
.A(n_2293),
.Y(n_3410)
);

AND2x4_ASAP7_75t_L g3411 ( 
.A(n_2553),
.B(n_2281),
.Y(n_3411)
);

OAI21x1_ASAP7_75t_SL g3412 ( 
.A1(n_2770),
.A2(n_2799),
.B(n_2792),
.Y(n_3412)
);

A2O1A1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_2757),
.A2(n_2773),
.B(n_2254),
.C(n_2264),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3414)
);

OAI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_2254),
.A2(n_2264),
.B1(n_2761),
.B2(n_2746),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2314),
.Y(n_3418)
);

OAI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_2254),
.A2(n_1490),
.B(n_1466),
.Y(n_3419)
);

AND2x2_ASAP7_75t_L g3420 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2314),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_2548),
.Y(n_3422)
);

AND2x4_ASAP7_75t_L g3423 ( 
.A(n_2553),
.B(n_2281),
.Y(n_3423)
);

OR2x2_ASAP7_75t_L g3424 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3424)
);

A2O1A1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_2757),
.A2(n_2773),
.B(n_2254),
.C(n_2264),
.Y(n_3425)
);

NAND2xp33_ASAP7_75t_L g3426 ( 
.A(n_2285),
.B(n_1480),
.Y(n_3426)
);

INVxp67_ASAP7_75t_L g3427 ( 
.A(n_2439),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3428)
);

AO21x1_ASAP7_75t_L g3429 ( 
.A1(n_2256),
.A2(n_2760),
.B(n_2753),
.Y(n_3429)
);

AND2x2_ASAP7_75t_SL g3430 ( 
.A(n_2737),
.B(n_2346),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_2293),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3435)
);

BUFx12f_ASAP7_75t_L g3436 ( 
.A(n_2809),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3439)
);

NAND3xp33_ASAP7_75t_L g3440 ( 
.A(n_2254),
.B(n_2264),
.C(n_2271),
.Y(n_3440)
);

AOI21xp5_ASAP7_75t_L g3441 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3441)
);

HB1xp67_ASAP7_75t_L g3442 ( 
.A(n_2527),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_2346),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_2447),
.B(n_2456),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_2757),
.A2(n_2773),
.B(n_2254),
.C(n_2264),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3448)
);

NAND2x1p5_ASAP7_75t_L g3449 ( 
.A(n_2346),
.B(n_2453),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2264),
.A2(n_2256),
.B1(n_2254),
.B2(n_2753),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_2260),
.A2(n_1380),
.B(n_1374),
.Y(n_3452)
);

AOI21xp33_ASAP7_75t_L g3453 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_3453)
);

INVxp67_ASAP7_75t_L g3454 ( 
.A(n_2439),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_2295),
.B(n_2750),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_2749),
.B(n_2788),
.Y(n_3456)
);

BUFx6f_ASAP7_75t_L g3457 ( 
.A(n_2346),
.Y(n_3457)
);

AO31x2_ASAP7_75t_L g3458 ( 
.A1(n_2471),
.A2(n_1447),
.A3(n_2373),
.B(n_2805),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2314),
.Y(n_3459)
);

CKINVDCx5p33_ASAP7_75t_R g3460 ( 
.A(n_2548),
.Y(n_3460)
);

AOI21xp33_ASAP7_75t_L g3461 ( 
.A1(n_2259),
.A2(n_2264),
.B(n_2753),
.Y(n_3461)
);

INVx6_ASAP7_75t_SL g3462 ( 
.A(n_2995),
.Y(n_3462)
);

INVx3_ASAP7_75t_SL g3463 ( 
.A(n_2911),
.Y(n_3463)
);

BUFx2_ASAP7_75t_SL g3464 ( 
.A(n_3359),
.Y(n_3464)
);

OR2x6_ASAP7_75t_L g3465 ( 
.A(n_2995),
.B(n_3397),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2888),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3282),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_2939),
.B(n_2947),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_2953),
.B(n_2970),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2888),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_2910),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2910),
.Y(n_3472)
);

INVx3_ASAP7_75t_SL g3473 ( 
.A(n_3017),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_2939),
.B(n_2947),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2905),
.B(n_2908),
.Y(n_3475)
);

BUFx3_ASAP7_75t_L g3476 ( 
.A(n_3297),
.Y(n_3476)
);

BUFx12f_ASAP7_75t_L g3477 ( 
.A(n_3018),
.Y(n_3477)
);

INVx2_ASAP7_75t_SL g3478 ( 
.A(n_3266),
.Y(n_3478)
);

INVx3_ASAP7_75t_L g3479 ( 
.A(n_3114),
.Y(n_3479)
);

INVxp67_ASAP7_75t_SL g3480 ( 
.A(n_2891),
.Y(n_3480)
);

BUFx3_ASAP7_75t_L g3481 ( 
.A(n_3297),
.Y(n_3481)
);

INVx5_ASAP7_75t_L g3482 ( 
.A(n_2995),
.Y(n_3482)
);

BUFx12f_ASAP7_75t_L g3483 ( 
.A(n_3049),
.Y(n_3483)
);

CKINVDCx20_ASAP7_75t_R g3484 ( 
.A(n_2942),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_2953),
.B(n_2970),
.Y(n_3485)
);

INVx5_ASAP7_75t_L g3486 ( 
.A(n_2995),
.Y(n_3486)
);

INVx5_ASAP7_75t_L g3487 ( 
.A(n_2995),
.Y(n_3487)
);

INVx5_ASAP7_75t_L g3488 ( 
.A(n_3397),
.Y(n_3488)
);

INVx4_ASAP7_75t_L g3489 ( 
.A(n_3300),
.Y(n_3489)
);

INVx3_ASAP7_75t_SL g3490 ( 
.A(n_2973),
.Y(n_3490)
);

INVx5_ASAP7_75t_L g3491 ( 
.A(n_3397),
.Y(n_3491)
);

INVx3_ASAP7_75t_L g3492 ( 
.A(n_3114),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3282),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_2905),
.B(n_2908),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3275),
.Y(n_3495)
);

BUFx3_ASAP7_75t_L g3496 ( 
.A(n_2887),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2901),
.B(n_2912),
.Y(n_3497)
);

NAND2x1p5_ASAP7_75t_L g3498 ( 
.A(n_3334),
.B(n_3430),
.Y(n_3498)
);

BUFx3_ASAP7_75t_L g3499 ( 
.A(n_2887),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2909),
.B(n_2932),
.Y(n_3500)
);

BUFx4_ASAP7_75t_SL g3501 ( 
.A(n_3346),
.Y(n_3501)
);

INVxp67_ASAP7_75t_SL g3502 ( 
.A(n_3389),
.Y(n_3502)
);

INVxp67_ASAP7_75t_SL g3503 ( 
.A(n_3035),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3318),
.B(n_3326),
.Y(n_3504)
);

BUFx2_ASAP7_75t_L g3505 ( 
.A(n_3156),
.Y(n_3505)
);

BUFx4_ASAP7_75t_SL g3506 ( 
.A(n_3268),
.Y(n_3506)
);

INVx3_ASAP7_75t_L g3507 ( 
.A(n_3121),
.Y(n_3507)
);

BUFx2_ASAP7_75t_L g3508 ( 
.A(n_3156),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3275),
.Y(n_3509)
);

NOR2x1_ASAP7_75t_SL g3510 ( 
.A(n_3397),
.B(n_3292),
.Y(n_3510)
);

INVx3_ASAP7_75t_L g3511 ( 
.A(n_3121),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_2906),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2925),
.Y(n_3513)
);

BUFx12f_ASAP7_75t_L g3514 ( 
.A(n_3422),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3358),
.B(n_2897),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3275),
.Y(n_3516)
);

INVx4_ASAP7_75t_L g3517 ( 
.A(n_3300),
.Y(n_3517)
);

INVx2_ASAP7_75t_SL g3518 ( 
.A(n_3266),
.Y(n_3518)
);

INVx2_ASAP7_75t_SL g3519 ( 
.A(n_3266),
.Y(n_3519)
);

INVx3_ASAP7_75t_L g3520 ( 
.A(n_2964),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3275),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3318),
.B(n_3326),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3281),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_2925),
.Y(n_3524)
);

INVx5_ASAP7_75t_L g3525 ( 
.A(n_3397),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_3117),
.Y(n_3526)
);

AND2x2_ASAP7_75t_L g3527 ( 
.A(n_3420),
.B(n_3432),
.Y(n_3527)
);

CKINVDCx20_ASAP7_75t_R g3528 ( 
.A(n_3150),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2909),
.B(n_2938),
.Y(n_3529)
);

CKINVDCx16_ASAP7_75t_R g3530 ( 
.A(n_3337),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3281),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_2960),
.Y(n_3532)
);

CKINVDCx20_ASAP7_75t_R g3533 ( 
.A(n_3033),
.Y(n_3533)
);

INVx3_ASAP7_75t_L g3534 ( 
.A(n_2964),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3266),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_2907),
.Y(n_3536)
);

BUFx2_ASAP7_75t_L g3537 ( 
.A(n_2906),
.Y(n_3537)
);

NAND2x1p5_ASAP7_75t_L g3538 ( 
.A(n_3334),
.B(n_3430),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3281),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2960),
.Y(n_3540)
);

BUFx2_ASAP7_75t_L g3541 ( 
.A(n_2934),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3420),
.B(n_3432),
.Y(n_3542)
);

CKINVDCx20_ASAP7_75t_R g3543 ( 
.A(n_3052),
.Y(n_3543)
);

BUFx3_ASAP7_75t_L g3544 ( 
.A(n_2907),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_2982),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_2967),
.B(n_2894),
.Y(n_3546)
);

BUFx3_ASAP7_75t_L g3547 ( 
.A(n_3176),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_2967),
.B(n_2914),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3324),
.A2(n_3393),
.B1(n_3416),
.B2(n_3408),
.Y(n_3549)
);

INVx3_ASAP7_75t_SL g3550 ( 
.A(n_3306),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_2982),
.Y(n_3551)
);

BUFx5_ASAP7_75t_L g3552 ( 
.A(n_3334),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2914),
.B(n_3358),
.Y(n_3553)
);

BUFx12f_ASAP7_75t_L g3554 ( 
.A(n_3460),
.Y(n_3554)
);

INVx1_ASAP7_75t_SL g3555 ( 
.A(n_3039),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_2934),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3006),
.Y(n_3557)
);

AND2x4_ASAP7_75t_L g3558 ( 
.A(n_3040),
.B(n_3285),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3006),
.Y(n_3559)
);

AND2x4_ASAP7_75t_L g3560 ( 
.A(n_3040),
.B(n_3285),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3359),
.B(n_3403),
.Y(n_3561)
);

BUFx12f_ASAP7_75t_L g3562 ( 
.A(n_3337),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3023),
.Y(n_3563)
);

HB1xp67_ASAP7_75t_L g3564 ( 
.A(n_3170),
.Y(n_3564)
);

BUFx6f_ASAP7_75t_L g3565 ( 
.A(n_3045),
.Y(n_3565)
);

OR2x6_ASAP7_75t_L g3566 ( 
.A(n_3292),
.B(n_3180),
.Y(n_3566)
);

INVx5_ASAP7_75t_L g3567 ( 
.A(n_3176),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_3176),
.Y(n_3568)
);

BUFx12f_ASAP7_75t_L g3569 ( 
.A(n_3337),
.Y(n_3569)
);

CKINVDCx16_ASAP7_75t_R g3570 ( 
.A(n_3436),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_3238),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3023),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3056),
.Y(n_3573)
);

INVx8_ASAP7_75t_L g3574 ( 
.A(n_3176),
.Y(n_3574)
);

BUFx3_ASAP7_75t_L g3575 ( 
.A(n_3176),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3056),
.Y(n_3576)
);

AO21x1_ASAP7_75t_L g3577 ( 
.A1(n_3350),
.A2(n_3366),
.B(n_3342),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3071),
.Y(n_3578)
);

INVx1_ASAP7_75t_SL g3579 ( 
.A(n_3039),
.Y(n_3579)
);

INVx3_ASAP7_75t_L g3580 ( 
.A(n_2943),
.Y(n_3580)
);

CKINVDCx20_ASAP7_75t_R g3581 ( 
.A(n_3052),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3445),
.B(n_2972),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3324),
.A2(n_3393),
.B1(n_3416),
.B2(n_3408),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_3176),
.Y(n_3584)
);

INVx1_ASAP7_75t_SL g3585 ( 
.A(n_2919),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_2935),
.B(n_2915),
.Y(n_3586)
);

OR2x6_ASAP7_75t_L g3587 ( 
.A(n_3180),
.B(n_3097),
.Y(n_3587)
);

HB1xp67_ASAP7_75t_L g3588 ( 
.A(n_2920),
.Y(n_3588)
);

INVx1_ASAP7_75t_SL g3589 ( 
.A(n_2919),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3071),
.Y(n_3590)
);

BUFx3_ASAP7_75t_L g3591 ( 
.A(n_3242),
.Y(n_3591)
);

BUFx3_ASAP7_75t_L g3592 ( 
.A(n_3242),
.Y(n_3592)
);

INVx1_ASAP7_75t_SL g3593 ( 
.A(n_2948),
.Y(n_3593)
);

INVx1_ASAP7_75t_SL g3594 ( 
.A(n_2948),
.Y(n_3594)
);

BUFx12f_ASAP7_75t_L g3595 ( 
.A(n_3436),
.Y(n_3595)
);

BUFx3_ASAP7_75t_L g3596 ( 
.A(n_3242),
.Y(n_3596)
);

INVx2_ASAP7_75t_SL g3597 ( 
.A(n_2926),
.Y(n_3597)
);

NAND2x1p5_ASAP7_75t_L g3598 ( 
.A(n_3430),
.B(n_3060),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3445),
.B(n_2972),
.Y(n_3599)
);

CKINVDCx6p67_ASAP7_75t_R g3600 ( 
.A(n_3436),
.Y(n_3600)
);

BUFx3_ASAP7_75t_L g3601 ( 
.A(n_3257),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_3090),
.Y(n_3602)
);

BUFx12f_ASAP7_75t_L g3603 ( 
.A(n_3212),
.Y(n_3603)
);

BUFx4_ASAP7_75t_SL g3604 ( 
.A(n_3268),
.Y(n_3604)
);

INVx5_ASAP7_75t_SL g3605 ( 
.A(n_3060),
.Y(n_3605)
);

OR2x6_ASAP7_75t_L g3606 ( 
.A(n_3180),
.B(n_3072),
.Y(n_3606)
);

INVx1_ASAP7_75t_SL g3607 ( 
.A(n_2897),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3257),
.Y(n_3608)
);

BUFx8_ASAP7_75t_SL g3609 ( 
.A(n_3212),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_2943),
.Y(n_3610)
);

BUFx6f_ASAP7_75t_SL g3611 ( 
.A(n_3060),
.Y(n_3611)
);

BUFx4f_ASAP7_75t_SL g3612 ( 
.A(n_3212),
.Y(n_3612)
);

INVx1_ASAP7_75t_SL g3613 ( 
.A(n_3392),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3075),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_2893),
.A2(n_2900),
.B1(n_3399),
.B2(n_3390),
.Y(n_3615)
);

CKINVDCx20_ASAP7_75t_R g3616 ( 
.A(n_3090),
.Y(n_3616)
);

BUFx12f_ASAP7_75t_L g3617 ( 
.A(n_3303),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3007),
.B(n_3042),
.Y(n_3618)
);

NAND2x1p5_ASAP7_75t_L g3619 ( 
.A(n_2987),
.B(n_3400),
.Y(n_3619)
);

INVx5_ASAP7_75t_SL g3620 ( 
.A(n_3180),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3075),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_3304),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3333),
.Y(n_3623)
);

BUFx5_ASAP7_75t_L g3624 ( 
.A(n_3040),
.Y(n_3624)
);

AND2x4_ASAP7_75t_L g3625 ( 
.A(n_3285),
.B(n_3230),
.Y(n_3625)
);

BUFx3_ASAP7_75t_L g3626 ( 
.A(n_2954),
.Y(n_3626)
);

NAND2x1p5_ASAP7_75t_L g3627 ( 
.A(n_2987),
.B(n_3400),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3333),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3403),
.B(n_3429),
.Y(n_3629)
);

NAND2x1p5_ASAP7_75t_L g3630 ( 
.A(n_2987),
.B(n_3400),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3335),
.Y(n_3631)
);

BUFx3_ASAP7_75t_L g3632 ( 
.A(n_2954),
.Y(n_3632)
);

INVx5_ASAP7_75t_L g3633 ( 
.A(n_3180),
.Y(n_3633)
);

INVx5_ASAP7_75t_L g3634 ( 
.A(n_2940),
.Y(n_3634)
);

BUFx6f_ASAP7_75t_L g3635 ( 
.A(n_3054),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3335),
.Y(n_3636)
);

INVx2_ASAP7_75t_SL g3637 ( 
.A(n_2926),
.Y(n_3637)
);

BUFx3_ASAP7_75t_L g3638 ( 
.A(n_2954),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3347),
.Y(n_3639)
);

INVx1_ASAP7_75t_SL g3640 ( 
.A(n_3392),
.Y(n_3640)
);

AO21x2_ASAP7_75t_L g3641 ( 
.A1(n_3206),
.A2(n_3245),
.B(n_3235),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_SL g3642 ( 
.A1(n_2900),
.A2(n_3399),
.B1(n_3440),
.B2(n_3390),
.Y(n_3642)
);

INVx1_ASAP7_75t_SL g3643 ( 
.A(n_3424),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3347),
.Y(n_3644)
);

BUFx3_ASAP7_75t_L g3645 ( 
.A(n_2968),
.Y(n_3645)
);

CKINVDCx14_ASAP7_75t_R g3646 ( 
.A(n_3142),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3007),
.B(n_3042),
.Y(n_3647)
);

BUFx6f_ASAP7_75t_L g3648 ( 
.A(n_3054),
.Y(n_3648)
);

INVx4_ASAP7_75t_L g3649 ( 
.A(n_3022),
.Y(n_3649)
);

BUFx3_ASAP7_75t_L g3650 ( 
.A(n_2968),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_2935),
.B(n_2915),
.Y(n_3651)
);

BUFx2_ASAP7_75t_R g3652 ( 
.A(n_2968),
.Y(n_3652)
);

INVx5_ASAP7_75t_L g3653 ( 
.A(n_2940),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3354),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3379),
.Y(n_3655)
);

INVx5_ASAP7_75t_L g3656 ( 
.A(n_2940),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3356),
.Y(n_3657)
);

INVxp33_ASAP7_75t_L g3658 ( 
.A(n_3182),
.Y(n_3658)
);

BUFx12f_ASAP7_75t_L g3659 ( 
.A(n_3303),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3451),
.A2(n_3342),
.B1(n_3331),
.B2(n_3440),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_2937),
.Y(n_3661)
);

INVx1_ASAP7_75t_SL g3662 ( 
.A(n_3424),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3356),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3378),
.Y(n_3664)
);

BUFx3_ASAP7_75t_L g3665 ( 
.A(n_3379),
.Y(n_3665)
);

BUFx12f_ASAP7_75t_L g3666 ( 
.A(n_3277),
.Y(n_3666)
);

BUFx2_ASAP7_75t_SL g3667 ( 
.A(n_3429),
.Y(n_3667)
);

AND2x4_ASAP7_75t_L g3668 ( 
.A(n_3230),
.B(n_3193),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3309),
.Y(n_3669)
);

INVx4_ASAP7_75t_L g3670 ( 
.A(n_3022),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3378),
.Y(n_3671)
);

INVx3_ASAP7_75t_SL g3672 ( 
.A(n_3280),
.Y(n_3672)
);

CKINVDCx20_ASAP7_75t_R g3673 ( 
.A(n_3194),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3418),
.Y(n_3674)
);

NOR2x1_ASAP7_75t_SL g3675 ( 
.A(n_3022),
.B(n_3032),
.Y(n_3675)
);

INVx4_ASAP7_75t_L g3676 ( 
.A(n_3022),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3205),
.B(n_3217),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3309),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3418),
.Y(n_3679)
);

BUFx12f_ASAP7_75t_L g3680 ( 
.A(n_3277),
.Y(n_3680)
);

BUFx3_ASAP7_75t_L g3681 ( 
.A(n_3379),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3218),
.B(n_3147),
.Y(n_3682)
);

BUFx12f_ASAP7_75t_L g3683 ( 
.A(n_3277),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_2981),
.Y(n_3684)
);

BUFx3_ASAP7_75t_L g3685 ( 
.A(n_3079),
.Y(n_3685)
);

INVx6_ASAP7_75t_SL g3686 ( 
.A(n_3193),
.Y(n_3686)
);

BUFx4_ASAP7_75t_SL g3687 ( 
.A(n_2985),
.Y(n_3687)
);

BUFx3_ASAP7_75t_L g3688 ( 
.A(n_3079),
.Y(n_3688)
);

INVx6_ASAP7_75t_L g3689 ( 
.A(n_3277),
.Y(n_3689)
);

BUFx12f_ASAP7_75t_L g3690 ( 
.A(n_3267),
.Y(n_3690)
);

BUFx2_ASAP7_75t_SL g3691 ( 
.A(n_2916),
.Y(n_3691)
);

INVx3_ASAP7_75t_L g3692 ( 
.A(n_3157),
.Y(n_3692)
);

BUFx12f_ASAP7_75t_L g3693 ( 
.A(n_3267),
.Y(n_3693)
);

INVx3_ASAP7_75t_L g3694 ( 
.A(n_3157),
.Y(n_3694)
);

AOI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3451),
.A2(n_2903),
.B1(n_2916),
.B2(n_2895),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3421),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3421),
.Y(n_3697)
);

CKINVDCx16_ASAP7_75t_R g3698 ( 
.A(n_3194),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_3255),
.Y(n_3699)
);

NAND2xp33_ASAP7_75t_SL g3700 ( 
.A(n_2929),
.B(n_2965),
.Y(n_3700)
);

INVx3_ASAP7_75t_L g3701 ( 
.A(n_2884),
.Y(n_3701)
);

CKINVDCx20_ASAP7_75t_R g3702 ( 
.A(n_3061),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3459),
.Y(n_3703)
);

INVxp67_ASAP7_75t_SL g3704 ( 
.A(n_3237),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3459),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_2885),
.B(n_2902),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_2903),
.A2(n_2895),
.B1(n_3313),
.B2(n_3308),
.Y(n_3707)
);

BUFx2_ASAP7_75t_SL g3708 ( 
.A(n_3325),
.Y(n_3708)
);

BUFx4_ASAP7_75t_SL g3709 ( 
.A(n_2985),
.Y(n_3709)
);

BUFx12f_ASAP7_75t_L g3710 ( 
.A(n_3267),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_2885),
.B(n_2902),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3314),
.Y(n_3712)
);

CKINVDCx20_ASAP7_75t_R g3713 ( 
.A(n_2998),
.Y(n_3713)
);

BUFx3_ASAP7_75t_L g3714 ( 
.A(n_3299),
.Y(n_3714)
);

BUFx3_ASAP7_75t_L g3715 ( 
.A(n_3299),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_2904),
.B(n_3311),
.Y(n_3716)
);

BUFx12f_ASAP7_75t_L g3717 ( 
.A(n_3267),
.Y(n_3717)
);

INVx3_ASAP7_75t_L g3718 ( 
.A(n_2884),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3236),
.Y(n_3719)
);

BUFx12f_ASAP7_75t_L g3720 ( 
.A(n_3001),
.Y(n_3720)
);

CKINVDCx5p33_ASAP7_75t_R g3721 ( 
.A(n_3184),
.Y(n_3721)
);

INVx3_ASAP7_75t_L g3722 ( 
.A(n_2884),
.Y(n_3722)
);

HB1xp67_ASAP7_75t_L g3723 ( 
.A(n_3372),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_2904),
.B(n_3311),
.Y(n_3724)
);

NAND2x1p5_ASAP7_75t_L g3725 ( 
.A(n_3298),
.B(n_2884),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3084),
.Y(n_3726)
);

CKINVDCx20_ASAP7_75t_R g3727 ( 
.A(n_3055),
.Y(n_3727)
);

CKINVDCx5p33_ASAP7_75t_R g3728 ( 
.A(n_2977),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3058),
.B(n_3068),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3084),
.Y(n_3730)
);

INVx6_ASAP7_75t_L g3731 ( 
.A(n_3032),
.Y(n_3731)
);

INVx1_ASAP7_75t_SL g3732 ( 
.A(n_3065),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3312),
.B(n_3332),
.Y(n_3733)
);

BUFx3_ASAP7_75t_L g3734 ( 
.A(n_3189),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3058),
.B(n_3068),
.Y(n_3735)
);

BUFx3_ASAP7_75t_L g3736 ( 
.A(n_3189),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3103),
.B(n_3105),
.Y(n_3737)
);

BUFx12f_ASAP7_75t_L g3738 ( 
.A(n_3001),
.Y(n_3738)
);

BUFx3_ASAP7_75t_L g3739 ( 
.A(n_3032),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3325),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_SL g3741 ( 
.A(n_2951),
.B(n_2941),
.Y(n_3741)
);

INVx1_ASAP7_75t_SL g3742 ( 
.A(n_3385),
.Y(n_3742)
);

INVx1_ASAP7_75t_SL g3743 ( 
.A(n_3442),
.Y(n_3743)
);

BUFx2_ASAP7_75t_L g3744 ( 
.A(n_3325),
.Y(n_3744)
);

NAND2x1p5_ASAP7_75t_L g3745 ( 
.A(n_3298),
.B(n_3357),
.Y(n_3745)
);

BUFx12f_ASAP7_75t_L g3746 ( 
.A(n_3001),
.Y(n_3746)
);

HB1xp67_ASAP7_75t_L g3747 ( 
.A(n_3234),
.Y(n_3747)
);

AND2x2_ASAP7_75t_SL g3748 ( 
.A(n_3287),
.B(n_2936),
.Y(n_3748)
);

BUFx2_ASAP7_75t_L g3749 ( 
.A(n_2951),
.Y(n_3749)
);

CKINVDCx5p33_ASAP7_75t_R g3750 ( 
.A(n_2977),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3314),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_SL g3752 ( 
.A1(n_2890),
.A2(n_3406),
.B1(n_3412),
.B2(n_2892),
.Y(n_3752)
);

HB1xp67_ASAP7_75t_L g3753 ( 
.A(n_3234),
.Y(n_3753)
);

CKINVDCx20_ASAP7_75t_R g3754 ( 
.A(n_3179),
.Y(n_3754)
);

BUFx4_ASAP7_75t_SL g3755 ( 
.A(n_3295),
.Y(n_3755)
);

CKINVDCx11_ASAP7_75t_R g3756 ( 
.A(n_3223),
.Y(n_3756)
);

OR2x6_ASAP7_75t_L g3757 ( 
.A(n_3072),
.B(n_3096),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3103),
.B(n_3105),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_L g3759 ( 
.A(n_2917),
.B(n_3377),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_2941),
.B(n_2971),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3322),
.Y(n_3761)
);

NAND2x1p5_ASAP7_75t_L g3762 ( 
.A(n_3002),
.B(n_3351),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3322),
.Y(n_3763)
);

BUFx2_ASAP7_75t_R g3764 ( 
.A(n_2986),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3312),
.B(n_3332),
.Y(n_3765)
);

INVx3_ASAP7_75t_L g3766 ( 
.A(n_3155),
.Y(n_3766)
);

CKINVDCx20_ASAP7_75t_R g3767 ( 
.A(n_3087),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3322),
.Y(n_3768)
);

INVxp67_ASAP7_75t_SL g3769 ( 
.A(n_2963),
.Y(n_3769)
);

INVx4_ASAP7_75t_L g3770 ( 
.A(n_3301),
.Y(n_3770)
);

INVx3_ASAP7_75t_L g3771 ( 
.A(n_3155),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3323),
.Y(n_3772)
);

BUFx6f_ASAP7_75t_SL g3773 ( 
.A(n_3443),
.Y(n_3773)
);

HB1xp67_ASAP7_75t_L g3774 ( 
.A(n_3228),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_L g3775 ( 
.A(n_3426),
.B(n_2896),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3323),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3323),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_3183),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3169),
.B(n_3221),
.Y(n_3779)
);

CKINVDCx20_ASAP7_75t_R g3780 ( 
.A(n_3089),
.Y(n_3780)
);

BUFx2_ASAP7_75t_L g3781 ( 
.A(n_3183),
.Y(n_3781)
);

INVxp67_ASAP7_75t_SL g3782 ( 
.A(n_2963),
.Y(n_3782)
);

BUFx3_ASAP7_75t_L g3783 ( 
.A(n_2886),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3149),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3149),
.Y(n_3785)
);

BUFx2_ASAP7_75t_SL g3786 ( 
.A(n_3009),
.Y(n_3786)
);

INVxp67_ASAP7_75t_SL g3787 ( 
.A(n_2963),
.Y(n_3787)
);

INVx1_ASAP7_75t_SL g3788 ( 
.A(n_3083),
.Y(n_3788)
);

BUFx2_ASAP7_75t_L g3789 ( 
.A(n_3064),
.Y(n_3789)
);

BUFx2_ASAP7_75t_SL g3790 ( 
.A(n_3009),
.Y(n_3790)
);

BUFx2_ASAP7_75t_R g3791 ( 
.A(n_3046),
.Y(n_3791)
);

CKINVDCx5p33_ASAP7_75t_R g3792 ( 
.A(n_3146),
.Y(n_3792)
);

CKINVDCx5p33_ASAP7_75t_R g3793 ( 
.A(n_2889),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3340),
.Y(n_3794)
);

INVx1_ASAP7_75t_SL g3795 ( 
.A(n_3083),
.Y(n_3795)
);

INVx1_ASAP7_75t_SL g3796 ( 
.A(n_3371),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_L g3797 ( 
.A(n_3457),
.Y(n_3797)
);

INVx4_ASAP7_75t_L g3798 ( 
.A(n_3301),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3164),
.Y(n_3799)
);

BUFx2_ASAP7_75t_L g3800 ( 
.A(n_3164),
.Y(n_3800)
);

BUFx4_ASAP7_75t_SL g3801 ( 
.A(n_3223),
.Y(n_3801)
);

INVx1_ASAP7_75t_SL g3802 ( 
.A(n_3375),
.Y(n_3802)
);

BUFx12f_ASAP7_75t_L g3803 ( 
.A(n_3034),
.Y(n_3803)
);

NAND2x1p5_ASAP7_75t_L g3804 ( 
.A(n_3041),
.B(n_3107),
.Y(n_3804)
);

INVx3_ASAP7_75t_L g3805 ( 
.A(n_3119),
.Y(n_3805)
);

BUFx2_ASAP7_75t_L g3806 ( 
.A(n_2950),
.Y(n_3806)
);

INVx2_ASAP7_75t_SL g3807 ( 
.A(n_3041),
.Y(n_3807)
);

CKINVDCx11_ASAP7_75t_R g3808 ( 
.A(n_3223),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_2896),
.B(n_2946),
.Y(n_3809)
);

INVx1_ASAP7_75t_SL g3810 ( 
.A(n_3375),
.Y(n_3810)
);

BUFx2_ASAP7_75t_SL g3811 ( 
.A(n_3059),
.Y(n_3811)
);

INVx2_ASAP7_75t_SL g3812 ( 
.A(n_3221),
.Y(n_3812)
);

HB1xp67_ASAP7_75t_L g3813 ( 
.A(n_3228),
.Y(n_3813)
);

BUFx2_ASAP7_75t_L g3814 ( 
.A(n_2950),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3340),
.Y(n_3815)
);

INVx1_ASAP7_75t_SL g3816 ( 
.A(n_3376),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3340),
.Y(n_3817)
);

BUFx12f_ASAP7_75t_L g3818 ( 
.A(n_3034),
.Y(n_3818)
);

INVx3_ASAP7_75t_L g3819 ( 
.A(n_3119),
.Y(n_3819)
);

BUFx2_ASAP7_75t_SL g3820 ( 
.A(n_2997),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3343),
.Y(n_3821)
);

CKINVDCx8_ASAP7_75t_R g3822 ( 
.A(n_3034),
.Y(n_3822)
);

BUFx2_ASAP7_75t_L g3823 ( 
.A(n_2950),
.Y(n_3823)
);

NOR2xp33_ASAP7_75t_L g3824 ( 
.A(n_2946),
.B(n_3308),
.Y(n_3824)
);

INVx1_ASAP7_75t_SL g3825 ( 
.A(n_3387),
.Y(n_3825)
);

BUFx12f_ASAP7_75t_L g3826 ( 
.A(n_3034),
.Y(n_3826)
);

AND2x4_ASAP7_75t_L g3827 ( 
.A(n_3197),
.B(n_3011),
.Y(n_3827)
);

BUFx12f_ASAP7_75t_L g3828 ( 
.A(n_3034),
.Y(n_3828)
);

NAND2x1p5_ASAP7_75t_L g3829 ( 
.A(n_3110),
.B(n_3020),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3343),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3343),
.Y(n_3831)
);

BUFx4f_ASAP7_75t_SL g3832 ( 
.A(n_3036),
.Y(n_3832)
);

OAI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3313),
.A2(n_3453),
.B1(n_3461),
.B2(n_3383),
.Y(n_3833)
);

CKINVDCx8_ASAP7_75t_R g3834 ( 
.A(n_3036),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2975),
.Y(n_3835)
);

INVx2_ASAP7_75t_SL g3836 ( 
.A(n_3229),
.Y(n_3836)
);

BUFx2_ASAP7_75t_L g3837 ( 
.A(n_2950),
.Y(n_3837)
);

INVx1_ASAP7_75t_SL g3838 ( 
.A(n_3391),
.Y(n_3838)
);

BUFx6f_ASAP7_75t_L g3839 ( 
.A(n_3073),
.Y(n_3839)
);

NAND2x1p5_ASAP7_75t_L g3840 ( 
.A(n_3020),
.B(n_3025),
.Y(n_3840)
);

NAND2x1p5_ASAP7_75t_L g3841 ( 
.A(n_3025),
.B(n_3098),
.Y(n_3841)
);

INVx3_ASAP7_75t_L g3842 ( 
.A(n_3131),
.Y(n_3842)
);

BUFx6f_ASAP7_75t_L g3843 ( 
.A(n_3073),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3363),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3363),
.Y(n_3845)
);

BUFx2_ASAP7_75t_L g3846 ( 
.A(n_2980),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_2975),
.Y(n_3847)
);

INVx4_ASAP7_75t_L g3848 ( 
.A(n_3036),
.Y(n_3848)
);

BUFx12f_ASAP7_75t_L g3849 ( 
.A(n_3036),
.Y(n_3849)
);

CKINVDCx16_ASAP7_75t_R g3850 ( 
.A(n_3287),
.Y(n_3850)
);

CKINVDCx5p33_ASAP7_75t_R g3851 ( 
.A(n_2898),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3363),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2988),
.Y(n_3853)
);

BUFx2_ASAP7_75t_L g3854 ( 
.A(n_2980),
.Y(n_3854)
);

OAI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3383),
.A2(n_3453),
.B1(n_3461),
.B2(n_2936),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_2988),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3369),
.Y(n_3857)
);

INVx2_ASAP7_75t_SL g3858 ( 
.A(n_3229),
.Y(n_3858)
);

AOI22xp33_ASAP7_75t_L g3859 ( 
.A1(n_2922),
.A2(n_2892),
.B1(n_3406),
.B2(n_2890),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_L g3860 ( 
.A1(n_3412),
.A2(n_2965),
.B1(n_3339),
.B2(n_3328),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_3135),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_2989),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_2989),
.Y(n_3863)
);

BUFx8_ASAP7_75t_SL g3864 ( 
.A(n_3030),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3328),
.A2(n_3339),
.B1(n_3386),
.B2(n_3380),
.Y(n_3865)
);

INVx2_ASAP7_75t_SL g3866 ( 
.A(n_3003),
.Y(n_3866)
);

INVx6_ASAP7_75t_SL g3867 ( 
.A(n_3411),
.Y(n_3867)
);

BUFx8_ASAP7_75t_L g3868 ( 
.A(n_3037),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_3135),
.Y(n_3869)
);

BUFx8_ASAP7_75t_L g3870 ( 
.A(n_3037),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3369),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3169),
.B(n_3274),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_2992),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_2992),
.Y(n_3874)
);

AOI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3341),
.A2(n_3413),
.B1(n_3425),
.B2(n_3370),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3423),
.B(n_3166),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3369),
.Y(n_3877)
);

BUFx10_ASAP7_75t_L g3878 ( 
.A(n_3130),
.Y(n_3878)
);

INVx4_ASAP7_75t_L g3879 ( 
.A(n_3037),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_2993),
.Y(n_3880)
);

INVx1_ASAP7_75t_SL g3881 ( 
.A(n_3394),
.Y(n_3881)
);

BUFx4_ASAP7_75t_SL g3882 ( 
.A(n_3261),
.Y(n_3882)
);

CKINVDCx5p33_ASAP7_75t_R g3883 ( 
.A(n_2921),
.Y(n_3883)
);

INVx4_ASAP7_75t_L g3884 ( 
.A(n_3122),
.Y(n_3884)
);

OR2x6_ASAP7_75t_L g3885 ( 
.A(n_3101),
.B(n_3099),
.Y(n_3885)
);

INVx1_ASAP7_75t_SL g3886 ( 
.A(n_3395),
.Y(n_3886)
);

INVx5_ASAP7_75t_L g3887 ( 
.A(n_3122),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3384),
.Y(n_3888)
);

BUFx3_ASAP7_75t_L g3889 ( 
.A(n_3210),
.Y(n_3889)
);

BUFx6f_ASAP7_75t_L g3890 ( 
.A(n_3019),
.Y(n_3890)
);

BUFx3_ASAP7_75t_L g3891 ( 
.A(n_3210),
.Y(n_3891)
);

OAI21xp33_ASAP7_75t_L g3892 ( 
.A1(n_2928),
.A2(n_2949),
.B(n_2923),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3384),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3384),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_3019),
.Y(n_3895)
);

CKINVDCx16_ASAP7_75t_R g3896 ( 
.A(n_2971),
.Y(n_3896)
);

NAND2x1p5_ASAP7_75t_L g3897 ( 
.A(n_2952),
.B(n_2969),
.Y(n_3897)
);

BUFx4_ASAP7_75t_SL g3898 ( 
.A(n_3196),
.Y(n_3898)
);

INVx4_ASAP7_75t_L g3899 ( 
.A(n_3122),
.Y(n_3899)
);

BUFx6f_ASAP7_75t_L g3900 ( 
.A(n_2899),
.Y(n_3900)
);

BUFx2_ASAP7_75t_SL g3901 ( 
.A(n_2997),
.Y(n_3901)
);

BUFx3_ASAP7_75t_L g3902 ( 
.A(n_3210),
.Y(n_3902)
);

BUFx4_ASAP7_75t_SL g3903 ( 
.A(n_3171),
.Y(n_3903)
);

AND2x4_ASAP7_75t_L g3904 ( 
.A(n_3166),
.B(n_3293),
.Y(n_3904)
);

INVx1_ASAP7_75t_SL g3905 ( 
.A(n_3401),
.Y(n_3905)
);

INVx3_ASAP7_75t_SL g3906 ( 
.A(n_3122),
.Y(n_3906)
);

BUFx6f_ASAP7_75t_L g3907 ( 
.A(n_2899),
.Y(n_3907)
);

INVx3_ASAP7_75t_L g3908 ( 
.A(n_3141),
.Y(n_3908)
);

BUFx4f_ASAP7_75t_SL g3909 ( 
.A(n_3122),
.Y(n_3909)
);

CKINVDCx5p33_ASAP7_75t_R g3910 ( 
.A(n_3353),
.Y(n_3910)
);

BUFx3_ASAP7_75t_L g3911 ( 
.A(n_3000),
.Y(n_3911)
);

INVx5_ASAP7_75t_L g3912 ( 
.A(n_3125),
.Y(n_3912)
);

BUFx3_ASAP7_75t_L g3913 ( 
.A(n_3000),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3404),
.B(n_3407),
.Y(n_3914)
);

BUFx10_ASAP7_75t_L g3915 ( 
.A(n_3125),
.Y(n_3915)
);

BUFx2_ASAP7_75t_SL g3916 ( 
.A(n_2990),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_3081),
.Y(n_3917)
);

AND2x4_ASAP7_75t_L g3918 ( 
.A(n_3293),
.B(n_3207),
.Y(n_3918)
);

INVx6_ASAP7_75t_SL g3919 ( 
.A(n_2958),
.Y(n_3919)
);

AOI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3447),
.A2(n_3386),
.B1(n_3388),
.B2(n_3380),
.Y(n_3920)
);

NOR2x1_ASAP7_75t_SL g3921 ( 
.A(n_3220),
.B(n_3227),
.Y(n_3921)
);

INVx2_ASAP7_75t_SL g3922 ( 
.A(n_3003),
.Y(n_3922)
);

AND2x4_ASAP7_75t_L g3923 ( 
.A(n_3207),
.B(n_3209),
.Y(n_3923)
);

BUFx3_ASAP7_75t_L g3924 ( 
.A(n_3081),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3141),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_3081),
.Y(n_3926)
);

NAND2x1p5_ASAP7_75t_L g3927 ( 
.A(n_3104),
.B(n_3115),
.Y(n_3927)
);

BUFx3_ASAP7_75t_L g3928 ( 
.A(n_3085),
.Y(n_3928)
);

BUFx6f_ASAP7_75t_L g3929 ( 
.A(n_2961),
.Y(n_3929)
);

BUFx3_ASAP7_75t_L g3930 ( 
.A(n_3085),
.Y(n_3930)
);

BUFx6f_ASAP7_75t_L g3931 ( 
.A(n_2961),
.Y(n_3931)
);

INVx1_ASAP7_75t_SL g3932 ( 
.A(n_3404),
.Y(n_3932)
);

CKINVDCx20_ASAP7_75t_R g3933 ( 
.A(n_2929),
.Y(n_3933)
);

CKINVDCx20_ASAP7_75t_R g3934 ( 
.A(n_3321),
.Y(n_3934)
);

BUFx3_ASAP7_75t_L g3935 ( 
.A(n_3085),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3793),
.B(n_3456),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3466),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3495),
.Y(n_3938)
);

AOI32xp33_ASAP7_75t_L g3939 ( 
.A1(n_3700),
.A2(n_3396),
.A3(n_3140),
.B1(n_2996),
.B2(n_3043),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3549),
.A2(n_2974),
.B(n_2944),
.Y(n_3940)
);

OAI22xp5_ASAP7_75t_L g3941 ( 
.A1(n_3865),
.A2(n_3402),
.B1(n_3415),
.B2(n_3388),
.Y(n_3941)
);

AND2x4_ASAP7_75t_L g3942 ( 
.A(n_3567),
.B(n_3249),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3466),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3577),
.A2(n_3152),
.B1(n_3092),
.B2(n_2918),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3567),
.B(n_3253),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3546),
.B(n_3405),
.Y(n_3946)
);

AND2x6_ASAP7_75t_SL g3947 ( 
.A(n_3759),
.B(n_3008),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3495),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3577),
.A2(n_3642),
.B1(n_3660),
.B2(n_3865),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3470),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3470),
.Y(n_3951)
);

NAND2x1p5_ASAP7_75t_L g3952 ( 
.A(n_3749),
.B(n_3106),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_L g3953 ( 
.A(n_3851),
.B(n_3014),
.Y(n_3953)
);

NAND3xp33_ASAP7_75t_L g3954 ( 
.A(n_3892),
.B(n_2974),
.C(n_2949),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_3577),
.A2(n_3642),
.B1(n_3660),
.B2(n_3651),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_3501),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3749),
.B(n_3407),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3779),
.B(n_3274),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3471),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3471),
.Y(n_3960)
);

INVx3_ASAP7_75t_L g3961 ( 
.A(n_3479),
.Y(n_3961)
);

CKINVDCx11_ASAP7_75t_R g3962 ( 
.A(n_3484),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3549),
.A2(n_3583),
.B(n_3920),
.Y(n_3963)
);

NOR2xp67_ASAP7_75t_L g3964 ( 
.A(n_3567),
.B(n_3805),
.Y(n_3964)
);

BUFx6f_ASAP7_75t_L g3965 ( 
.A(n_3890),
.Y(n_3965)
);

OAI22xp5_ASAP7_75t_L g3966 ( 
.A1(n_3860),
.A2(n_3415),
.B1(n_3419),
.B2(n_3402),
.Y(n_3966)
);

BUFx3_ASAP7_75t_L g3967 ( 
.A(n_3562),
.Y(n_3967)
);

A2O1A1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3892),
.A2(n_3809),
.B(n_3775),
.C(n_3695),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3472),
.Y(n_3969)
);

OAI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3583),
.A2(n_3092),
.B1(n_3419),
.B2(n_2955),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3472),
.Y(n_3971)
);

OAI22xp33_ASAP7_75t_L g3972 ( 
.A1(n_3920),
.A2(n_2955),
.B1(n_3140),
.B2(n_2918),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3741),
.A2(n_2930),
.B(n_3316),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_3867),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3651),
.A2(n_3152),
.B1(n_3132),
.B2(n_2990),
.Y(n_3975)
);

BUFx6f_ASAP7_75t_L g3976 ( 
.A(n_3890),
.Y(n_3976)
);

INVx2_ASAP7_75t_SL g3977 ( 
.A(n_3496),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3509),
.Y(n_3978)
);

NAND2xp33_ASAP7_75t_SL g3979 ( 
.A(n_3728),
.B(n_3750),
.Y(n_3979)
);

INVx3_ASAP7_75t_SL g3980 ( 
.A(n_3600),
.Y(n_3980)
);

AO31x2_ASAP7_75t_L g3981 ( 
.A1(n_3500),
.A2(n_2994),
.A3(n_3251),
.B(n_3269),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3741),
.A2(n_2930),
.B(n_3316),
.Y(n_3982)
);

BUFx6f_ASAP7_75t_L g3983 ( 
.A(n_3890),
.Y(n_3983)
);

AO21x2_ASAP7_75t_L g3984 ( 
.A1(n_3503),
.A2(n_2994),
.B(n_3409),
.Y(n_3984)
);

INVx3_ASAP7_75t_L g3985 ( 
.A(n_3479),
.Y(n_3985)
);

OR2x2_ASAP7_75t_L g3986 ( 
.A(n_3607),
.B(n_3414),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3860),
.A2(n_3360),
.B1(n_2979),
.B2(n_2957),
.Y(n_3987)
);

INVxp67_ASAP7_75t_L g3988 ( 
.A(n_3774),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3546),
.B(n_3405),
.Y(n_3989)
);

CKINVDCx6p67_ASAP7_75t_R g3990 ( 
.A(n_3562),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_3562),
.Y(n_3991)
);

AO31x2_ASAP7_75t_L g3992 ( 
.A1(n_3500),
.A2(n_3251),
.A3(n_3269),
.B(n_3195),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3516),
.Y(n_3993)
);

OA21x2_ASAP7_75t_L g3994 ( 
.A1(n_3769),
.A2(n_3787),
.B(n_3782),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3468),
.B(n_3405),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3516),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3479),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3513),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3513),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3524),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3524),
.Y(n_4001)
);

HB1xp67_ASAP7_75t_L g4002 ( 
.A(n_3564),
.Y(n_4002)
);

A2O1A1Ixp33_ASAP7_75t_L g4003 ( 
.A1(n_3809),
.A2(n_3026),
.B(n_3154),
.C(n_2956),
.Y(n_4003)
);

CKINVDCx11_ASAP7_75t_R g4004 ( 
.A(n_3528),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_L g4005 ( 
.A(n_3824),
.B(n_2956),
.C(n_2991),
.Y(n_4005)
);

BUFx3_ASAP7_75t_L g4006 ( 
.A(n_3569),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3883),
.B(n_3038),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3521),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3521),
.Y(n_4009)
);

OAI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3494),
.A2(n_3132),
.B1(n_3109),
.B2(n_3106),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3532),
.Y(n_4011)
);

OAI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3561),
.A2(n_2991),
.B(n_3360),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3521),
.Y(n_4013)
);

CKINVDCx16_ASAP7_75t_R g4014 ( 
.A(n_3530),
.Y(n_4014)
);

OR2x2_ASAP7_75t_L g4015 ( 
.A(n_3607),
.B(n_3414),
.Y(n_4015)
);

A2O1A1Ixp33_ASAP7_75t_L g4016 ( 
.A1(n_3775),
.A2(n_3695),
.B(n_3824),
.C(n_3629),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3532),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3540),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3464),
.A2(n_3152),
.B1(n_3154),
.B2(n_3031),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3468),
.B(n_3405),
.Y(n_4020)
);

OR2x2_ASAP7_75t_L g4021 ( 
.A(n_3613),
.B(n_3417),
.Y(n_4021)
);

CKINVDCx14_ASAP7_75t_R g4022 ( 
.A(n_3543),
.Y(n_4022)
);

AOI221xp5_ASAP7_75t_L g4023 ( 
.A1(n_3833),
.A2(n_3855),
.B1(n_3475),
.B2(n_3494),
.C(n_3586),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3540),
.Y(n_4024)
);

CKINVDCx20_ASAP7_75t_R g4025 ( 
.A(n_3533),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3545),
.Y(n_4026)
);

O2A1O1Ixp33_ASAP7_75t_L g4027 ( 
.A1(n_3759),
.A2(n_3109),
.B(n_2976),
.C(n_2927),
.Y(n_4027)
);

BUFx3_ASAP7_75t_L g4028 ( 
.A(n_3569),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3545),
.Y(n_4029)
);

NAND2x1_ASAP7_75t_L g4030 ( 
.A(n_3606),
.B(n_2999),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3779),
.B(n_3320),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_SL g4032 ( 
.A1(n_3529),
.A2(n_3586),
.B(n_3139),
.Y(n_4032)
);

BUFx6f_ASAP7_75t_L g4033 ( 
.A(n_3890),
.Y(n_4033)
);

INVx6_ASAP7_75t_L g4034 ( 
.A(n_3567),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3551),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3474),
.B(n_3417),
.Y(n_4036)
);

HB1xp67_ASAP7_75t_L g4037 ( 
.A(n_3564),
.Y(n_4037)
);

CKINVDCx16_ASAP7_75t_R g4038 ( 
.A(n_3530),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3529),
.A2(n_2930),
.B(n_3315),
.Y(n_4039)
);

OAI221xp5_ASAP7_75t_L g4040 ( 
.A1(n_3875),
.A2(n_3088),
.B1(n_2966),
.B2(n_3136),
.C(n_3186),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_3501),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3615),
.A2(n_3329),
.B(n_3319),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3551),
.Y(n_4043)
);

HB1xp67_ASAP7_75t_L g4044 ( 
.A(n_3774),
.Y(n_4044)
);

BUFx6f_ASAP7_75t_L g4045 ( 
.A(n_3890),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3557),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3615),
.A2(n_3152),
.B1(n_2984),
.B2(n_3226),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3779),
.B(n_3361),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3557),
.Y(n_4049)
);

BUFx3_ASAP7_75t_L g4050 ( 
.A(n_3569),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3497),
.A2(n_2930),
.B(n_3704),
.Y(n_4051)
);

A2O1A1Ixp33_ASAP7_75t_L g4052 ( 
.A1(n_3707),
.A2(n_3088),
.B(n_3136),
.C(n_3198),
.Y(n_4052)
);

AO31x2_ASAP7_75t_L g4053 ( 
.A1(n_3799),
.A2(n_3291),
.A3(n_3365),
.B(n_2962),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_L g4054 ( 
.A(n_3910),
.B(n_3024),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3855),
.A2(n_2984),
.B1(n_3226),
.B2(n_3031),
.Y(n_4055)
);

AND2x6_ASAP7_75t_SL g4056 ( 
.A(n_3903),
.B(n_3077),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3559),
.Y(n_4057)
);

AOI22x1_ASAP7_75t_L g4058 ( 
.A1(n_3570),
.A2(n_3336),
.B1(n_3348),
.B2(n_3344),
.Y(n_4058)
);

OAI21xp5_ASAP7_75t_L g4059 ( 
.A1(n_3707),
.A2(n_3833),
.B(n_3760),
.Y(n_4059)
);

AO32x2_ASAP7_75t_L g4060 ( 
.A1(n_3597),
.A2(n_3227),
.A3(n_3021),
.B1(n_3012),
.B2(n_3214),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3559),
.Y(n_4061)
);

O2A1O1Ixp33_ASAP7_75t_SL g4062 ( 
.A1(n_3581),
.A2(n_3024),
.B(n_3124),
.C(n_3338),
.Y(n_4062)
);

BUFx3_ASAP7_75t_L g4063 ( 
.A(n_3595),
.Y(n_4063)
);

O2A1O1Ixp33_ASAP7_75t_L g4064 ( 
.A1(n_3497),
.A2(n_3381),
.B(n_3382),
.C(n_3352),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3563),
.Y(n_4065)
);

CKINVDCx16_ASAP7_75t_R g4066 ( 
.A(n_3570),
.Y(n_4066)
);

OAI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_3752),
.A2(n_3428),
.B(n_3398),
.Y(n_4067)
);

OAI21x1_ASAP7_75t_L g4068 ( 
.A1(n_3580),
.A2(n_3364),
.B(n_3317),
.Y(n_4068)
);

INVxp67_ASAP7_75t_SL g4069 ( 
.A(n_3480),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3563),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3572),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3464),
.A2(n_3215),
.B1(n_3133),
.B2(n_3177),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3580),
.A2(n_3610),
.B(n_3534),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3667),
.A2(n_3215),
.B1(n_3177),
.B2(n_3247),
.Y(n_4074)
);

BUFx2_ASAP7_75t_L g4075 ( 
.A(n_3867),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3469),
.B(n_3361),
.Y(n_4076)
);

BUFx3_ASAP7_75t_L g4077 ( 
.A(n_3595),
.Y(n_4077)
);

AOI21x1_ASAP7_75t_L g4078 ( 
.A1(n_3747),
.A2(n_3374),
.B(n_3373),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3469),
.B(n_3361),
.Y(n_4079)
);

A2O1A1Ixp33_ASAP7_75t_L g4080 ( 
.A1(n_3667),
.A2(n_3198),
.B(n_3153),
.C(n_3123),
.Y(n_4080)
);

HB1xp67_ASAP7_75t_L g4081 ( 
.A(n_3813),
.Y(n_4081)
);

AOI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_3875),
.A2(n_3933),
.B1(n_3550),
.B2(n_3896),
.Y(n_4082)
);

NOR2x1_ASAP7_75t_R g4083 ( 
.A(n_3595),
.B(n_2931),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3572),
.Y(n_4084)
);

INVx2_ASAP7_75t_SL g4085 ( 
.A(n_3496),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3469),
.B(n_3361),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3474),
.B(n_3438),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_3548),
.B(n_3438),
.Y(n_4088)
);

A2O1A1Ixp33_ASAP7_75t_L g4089 ( 
.A1(n_3691),
.A2(n_3790),
.B(n_3786),
.C(n_3518),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3573),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3573),
.Y(n_4091)
);

INVx3_ASAP7_75t_L g4092 ( 
.A(n_3479),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3666),
.Y(n_4093)
);

OAI21x1_ASAP7_75t_L g4094 ( 
.A1(n_3520),
.A2(n_3433),
.B(n_3410),
.Y(n_4094)
);

INVx6_ASAP7_75t_L g4095 ( 
.A(n_3567),
.Y(n_4095)
);

OAI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3752),
.A2(n_3434),
.B(n_3431),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3576),
.Y(n_4097)
);

OAI21x1_ASAP7_75t_L g4098 ( 
.A1(n_3534),
.A2(n_3433),
.B(n_3410),
.Y(n_4098)
);

CKINVDCx11_ASAP7_75t_R g4099 ( 
.A(n_3616),
.Y(n_4099)
);

BUFx3_ASAP7_75t_L g4100 ( 
.A(n_3666),
.Y(n_4100)
);

OAI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_3859),
.A2(n_3437),
.B(n_3435),
.Y(n_4101)
);

OAI21x1_ASAP7_75t_SL g4102 ( 
.A1(n_3921),
.A2(n_3365),
.B(n_2962),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3576),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_3613),
.B(n_3439),
.Y(n_4104)
);

AOI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3747),
.A2(n_3307),
.B(n_3264),
.Y(n_4105)
);

BUFx10_ASAP7_75t_L g4106 ( 
.A(n_3689),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3548),
.B(n_3439),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_SL g4108 ( 
.A1(n_3921),
.A2(n_3220),
.B(n_2999),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_3813),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3658),
.B(n_3864),
.Y(n_4110)
);

OAI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3859),
.A2(n_3448),
.B(n_3441),
.Y(n_4111)
);

NOR2xp33_ASAP7_75t_L g4112 ( 
.A(n_3721),
.B(n_3100),
.Y(n_4112)
);

INVxp67_ASAP7_75t_SL g4113 ( 
.A(n_3480),
.Y(n_4113)
);

OAI211xp5_ASAP7_75t_L g4114 ( 
.A1(n_3911),
.A2(n_3450),
.B(n_3452),
.C(n_3302),
.Y(n_4114)
);

INVx2_ASAP7_75t_SL g4115 ( 
.A(n_3496),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3578),
.Y(n_4116)
);

CKINVDCx20_ASAP7_75t_R g4117 ( 
.A(n_3673),
.Y(n_4117)
);

AND2x4_ASAP7_75t_L g4118 ( 
.A(n_3547),
.B(n_3222),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_3547),
.B(n_3222),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_3463),
.A2(n_3454),
.B1(n_3427),
.B2(n_3446),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3856),
.B(n_3444),
.Y(n_4121)
);

OAI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_3896),
.A2(n_2930),
.B1(n_2958),
.B2(n_3186),
.Y(n_4122)
);

OAI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3897),
.A2(n_3111),
.B(n_3192),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_L g4124 ( 
.A1(n_3550),
.A2(n_3247),
.B1(n_3051),
.B2(n_3069),
.Y(n_4124)
);

BUFx6f_ASAP7_75t_L g4125 ( 
.A(n_3890),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3578),
.Y(n_4126)
);

OA21x2_ASAP7_75t_L g4127 ( 
.A1(n_3523),
.A2(n_3539),
.B(n_3531),
.Y(n_4127)
);

AO21x2_ASAP7_75t_L g4128 ( 
.A1(n_3467),
.A2(n_3493),
.B(n_3523),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3590),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_3588),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3590),
.Y(n_4131)
);

NAND3xp33_ASAP7_75t_L g4132 ( 
.A(n_3553),
.B(n_3102),
.C(n_3051),
.Y(n_4132)
);

BUFx2_ASAP7_75t_L g4133 ( 
.A(n_3867),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3463),
.B(n_3208),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_3614),
.Y(n_4135)
);

INVx3_ASAP7_75t_L g4136 ( 
.A(n_3492),
.Y(n_4136)
);

AOI221xp5_ASAP7_75t_L g4137 ( 
.A1(n_3786),
.A2(n_3211),
.B1(n_3053),
.B2(n_3070),
.C(n_3086),
.Y(n_4137)
);

CKINVDCx5p33_ASAP7_75t_R g4138 ( 
.A(n_3571),
.Y(n_4138)
);

NAND2x1p5_ASAP7_75t_L g4139 ( 
.A(n_3633),
.B(n_3115),
.Y(n_4139)
);

OAI21x1_ASAP7_75t_L g4140 ( 
.A1(n_3661),
.A2(n_3082),
.B(n_3074),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3614),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_3621),
.Y(n_4142)
);

OAI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_3897),
.A2(n_3111),
.B(n_3192),
.Y(n_4143)
);

OR2x2_ASAP7_75t_L g4144 ( 
.A(n_3640),
.B(n_3444),
.Y(n_4144)
);

INVx3_ASAP7_75t_L g4145 ( 
.A(n_3492),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_3661),
.A2(n_3082),
.B(n_3074),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_3526),
.Y(n_4147)
);

BUFx2_ASAP7_75t_L g4148 ( 
.A(n_3867),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3621),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3623),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_3485),
.B(n_2983),
.Y(n_4151)
);

INVx2_ASAP7_75t_SL g4152 ( 
.A(n_3499),
.Y(n_4152)
);

INVx2_ASAP7_75t_SL g4153 ( 
.A(n_3499),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3856),
.B(n_3446),
.Y(n_4154)
);

OAI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3897),
.A2(n_3093),
.B(n_3161),
.Y(n_4155)
);

AND2x2_ASAP7_75t_L g4156 ( 
.A(n_3485),
.B(n_2983),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3623),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_3477),
.Y(n_4158)
);

OR2x6_ASAP7_75t_L g4159 ( 
.A(n_3574),
.B(n_3204),
.Y(n_4159)
);

OAI21x1_ASAP7_75t_SL g4160 ( 
.A1(n_3478),
.A2(n_3124),
.B(n_3231),
.Y(n_4160)
);

OAI22xp5_ASAP7_75t_SL g4161 ( 
.A1(n_3698),
.A2(n_3187),
.B1(n_3283),
.B2(n_3116),
.Y(n_4161)
);

CKINVDCx5p33_ASAP7_75t_R g4162 ( 
.A(n_3477),
.Y(n_4162)
);

BUFx2_ASAP7_75t_L g4163 ( 
.A(n_3867),
.Y(n_4163)
);

NAND2xp33_ASAP7_75t_SL g4164 ( 
.A(n_3463),
.B(n_3283),
.Y(n_4164)
);

OAI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3550),
.A2(n_3062),
.B1(n_3066),
.B2(n_3174),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3628),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_3485),
.B(n_2983),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3628),
.Y(n_4168)
);

NOR2xp67_ASAP7_75t_L g4169 ( 
.A(n_3805),
.B(n_3015),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_3631),
.Y(n_4170)
);

A2O1A1Ixp33_ASAP7_75t_L g4171 ( 
.A1(n_3691),
.A2(n_3790),
.B(n_3518),
.C(n_3519),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3502),
.B(n_3455),
.Y(n_4172)
);

NOR2x1_ASAP7_75t_R g4173 ( 
.A(n_3666),
.B(n_3048),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3631),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_3748),
.A2(n_2959),
.B1(n_3047),
.B2(n_3145),
.Y(n_4175)
);

AOI21x1_ASAP7_75t_L g4176 ( 
.A1(n_3753),
.A2(n_3094),
.B(n_3175),
.Y(n_4176)
);

OAI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_3757),
.A2(n_3455),
.B1(n_3200),
.B2(n_3259),
.Y(n_4177)
);

BUFx3_ASAP7_75t_L g4178 ( 
.A(n_3680),
.Y(n_4178)
);

OAI22xp33_ASAP7_75t_L g4179 ( 
.A1(n_3757),
.A2(n_3174),
.B1(n_3067),
.B2(n_3044),
.Y(n_4179)
);

BUFx3_ASAP7_75t_L g4180 ( 
.A(n_3680),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3636),
.Y(n_4181)
);

OAI21x1_ASAP7_75t_SL g4182 ( 
.A1(n_3478),
.A2(n_3254),
.B(n_3231),
.Y(n_4182)
);

BUFx2_ASAP7_75t_L g4183 ( 
.A(n_3686),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3636),
.Y(n_4184)
);

CKINVDCx6p67_ASAP7_75t_R g4185 ( 
.A(n_3600),
.Y(n_4185)
);

BUFx2_ASAP7_75t_L g4186 ( 
.A(n_3686),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3639),
.Y(n_4187)
);

AND2x6_ASAP7_75t_L g4188 ( 
.A(n_3605),
.B(n_3125),
.Y(n_4188)
);

OAI21xp5_ASAP7_75t_SL g4189 ( 
.A1(n_3478),
.A2(n_3519),
.B(n_3518),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_3748),
.A2(n_3086),
.B1(n_3053),
.B2(n_3069),
.Y(n_4190)
);

OAI21x1_ASAP7_75t_L g4191 ( 
.A1(n_3841),
.A2(n_3144),
.B(n_3094),
.Y(n_4191)
);

OAI21x1_ASAP7_75t_L g4192 ( 
.A1(n_3841),
.A2(n_3829),
.B(n_3819),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3639),
.Y(n_4193)
);

AO31x2_ASAP7_75t_L g4194 ( 
.A1(n_3800),
.A2(n_3028),
.A3(n_3016),
.B(n_3010),
.Y(n_4194)
);

INVx1_ASAP7_75t_SL g4195 ( 
.A(n_3585),
.Y(n_4195)
);

BUFx3_ASAP7_75t_L g4196 ( 
.A(n_3680),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3644),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3644),
.Y(n_4198)
);

OAI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_3757),
.A2(n_3161),
.B(n_3070),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_3504),
.B(n_2983),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3748),
.A2(n_2933),
.B1(n_2924),
.B2(n_3162),
.Y(n_4201)
);

BUFx3_ASAP7_75t_L g4202 ( 
.A(n_3683),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_3502),
.B(n_2933),
.Y(n_4203)
);

INVx8_ASAP7_75t_L g4204 ( 
.A(n_3574),
.Y(n_4204)
);

CKINVDCx20_ASAP7_75t_R g4205 ( 
.A(n_3609),
.Y(n_4205)
);

CKINVDCx5p33_ASAP7_75t_R g4206 ( 
.A(n_3477),
.Y(n_4206)
);

BUFx2_ASAP7_75t_SL g4207 ( 
.A(n_3499),
.Y(n_4207)
);

AO21x2_ASAP7_75t_L g4208 ( 
.A1(n_3493),
.A2(n_3254),
.B(n_3246),
.Y(n_4208)
);

AO21x2_ASAP7_75t_L g4209 ( 
.A1(n_3641),
.A2(n_3678),
.B(n_3669),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3796),
.B(n_3173),
.Y(n_4210)
);

INVx1_ASAP7_75t_SL g4211 ( 
.A(n_3585),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_3698),
.B(n_3148),
.Y(n_4212)
);

CKINVDCx6p67_ASAP7_75t_R g4213 ( 
.A(n_3600),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3657),
.Y(n_4214)
);

OAI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_3757),
.A2(n_3191),
.B(n_3027),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3657),
.Y(n_4216)
);

OAI21xp5_ASAP7_75t_SL g4217 ( 
.A1(n_3519),
.A2(n_3029),
.B(n_3159),
.Y(n_4217)
);

NOR2xp67_ASAP7_75t_L g4218 ( 
.A(n_3819),
.B(n_3148),
.Y(n_4218)
);

INVxp67_ASAP7_75t_L g4219 ( 
.A(n_3778),
.Y(n_4219)
);

OAI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_3757),
.A2(n_3244),
.B(n_3296),
.Y(n_4220)
);

INVx2_ASAP7_75t_SL g4221 ( 
.A(n_3536),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3796),
.B(n_3173),
.Y(n_4222)
);

A2O1A1Ixp33_ASAP7_75t_L g4223 ( 
.A1(n_3535),
.A2(n_3181),
.B(n_3172),
.C(n_3219),
.Y(n_4223)
);

CKINVDCx6p67_ASAP7_75t_R g4224 ( 
.A(n_3683),
.Y(n_4224)
);

OAI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_3757),
.A2(n_3764),
.B1(n_3535),
.B2(n_3791),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3504),
.B(n_3522),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3663),
.Y(n_4227)
);

O2A1O1Ixp33_ASAP7_75t_SL g4228 ( 
.A1(n_3903),
.A2(n_3279),
.B(n_3159),
.C(n_2924),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3663),
.Y(n_4229)
);

AOI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_3885),
.A2(n_3270),
.B(n_3284),
.Y(n_4230)
);

AOI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_3916),
.A2(n_3047),
.B1(n_2959),
.B2(n_2945),
.Y(n_4231)
);

OAI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_3764),
.A2(n_3213),
.B1(n_3188),
.B2(n_3216),
.Y(n_4232)
);

NOR2xp33_ASAP7_75t_L g4233 ( 
.A(n_3699),
.B(n_3190),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_3504),
.B(n_2983),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3522),
.B(n_2983),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3664),
.Y(n_4236)
);

OAI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_3553),
.A2(n_3241),
.B(n_3262),
.Y(n_4237)
);

OR2x6_ASAP7_75t_L g4238 ( 
.A(n_3574),
.B(n_3270),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_3522),
.B(n_3076),
.Y(n_4239)
);

O2A1O1Ixp33_ASAP7_75t_SL g4240 ( 
.A1(n_3732),
.A2(n_3028),
.B(n_3016),
.C(n_3010),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_3527),
.B(n_3076),
.Y(n_4241)
);

INVx4_ASAP7_75t_L g4242 ( 
.A(n_3689),
.Y(n_4242)
);

AOI21x1_ASAP7_75t_L g4243 ( 
.A1(n_3753),
.A2(n_3005),
.B(n_3004),
.Y(n_4243)
);

AOI22xp5_ASAP7_75t_L g4244 ( 
.A1(n_3780),
.A2(n_3162),
.B1(n_2945),
.B2(n_3449),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_3885),
.A2(n_3284),
.B(n_3294),
.Y(n_4245)
);

CKINVDCx20_ASAP7_75t_R g4246 ( 
.A(n_3767),
.Y(n_4246)
);

INVx5_ASAP7_75t_L g4247 ( 
.A(n_3606),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_3527),
.B(n_3076),
.Y(n_4248)
);

NOR2xp33_ASAP7_75t_SL g4249 ( 
.A(n_3791),
.B(n_2913),
.Y(n_4249)
);

HB1xp67_ASAP7_75t_L g4250 ( 
.A(n_3588),
.Y(n_4250)
);

AOI22xp33_ASAP7_75t_SL g4251 ( 
.A1(n_3820),
.A2(n_3458),
.B1(n_3367),
.B2(n_3349),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3664),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_3483),
.Y(n_4253)
);

AND2x2_ASAP7_75t_SL g4254 ( 
.A(n_3800),
.B(n_3162),
.Y(n_4254)
);

AOI22xp33_ASAP7_75t_L g4255 ( 
.A1(n_3611),
.A2(n_3252),
.B1(n_2945),
.B2(n_3449),
.Y(n_4255)
);

CKINVDCx11_ASAP7_75t_R g4256 ( 
.A(n_3483),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3671),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_3885),
.A2(n_3294),
.B(n_3288),
.Y(n_4258)
);

O2A1O1Ixp33_ASAP7_75t_SL g4259 ( 
.A1(n_3732),
.A2(n_3233),
.B(n_3167),
.C(n_3168),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3671),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_L g4261 ( 
.A(n_3654),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3674),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_3527),
.B(n_3076),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3674),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3679),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_3643),
.B(n_3662),
.Y(n_4266)
);

OAI221xp5_ASAP7_75t_L g4267 ( 
.A1(n_3820),
.A2(n_3224),
.B1(n_3240),
.B2(n_3158),
.C(n_3167),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3802),
.B(n_3310),
.Y(n_4268)
);

AOI22xp33_ASAP7_75t_L g4269 ( 
.A1(n_3611),
.A2(n_3252),
.B1(n_3449),
.B2(n_3368),
.Y(n_4269)
);

OAI21x1_ASAP7_75t_SL g4270 ( 
.A1(n_3535),
.A2(n_3134),
.B(n_3168),
.Y(n_4270)
);

OAI22x1_ASAP7_75t_L g4271 ( 
.A1(n_3598),
.A2(n_3272),
.B1(n_3202),
.B2(n_3201),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3679),
.Y(n_4272)
);

NAND2x1_ASAP7_75t_L g4273 ( 
.A(n_3606),
.B(n_3225),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_3802),
.B(n_3810),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_3591),
.B(n_3143),
.Y(n_4275)
);

AOI22xp33_ASAP7_75t_L g4276 ( 
.A1(n_3611),
.A2(n_3252),
.B1(n_3368),
.B2(n_3362),
.Y(n_4276)
);

AO21x1_ASAP7_75t_L g4277 ( 
.A1(n_3927),
.A2(n_3108),
.B(n_3138),
.Y(n_4277)
);

OAI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_3778),
.A2(n_3258),
.B(n_3263),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_3696),
.Y(n_4279)
);

AOI21xp33_ASAP7_75t_SL g4280 ( 
.A1(n_3602),
.A2(n_2913),
.B(n_3368),
.Y(n_4280)
);

AOI22xp33_ASAP7_75t_L g4281 ( 
.A1(n_3611),
.A2(n_3252),
.B1(n_3362),
.B2(n_3345),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3696),
.Y(n_4282)
);

AOI22xp33_ASAP7_75t_L g4283 ( 
.A1(n_3916),
.A2(n_3362),
.B1(n_3345),
.B2(n_3305),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3810),
.B(n_3367),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_3568),
.B(n_3076),
.Y(n_4285)
);

BUFx2_ASAP7_75t_L g4286 ( 
.A(n_3686),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_3483),
.B(n_3112),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_3542),
.B(n_3458),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3816),
.B(n_3458),
.Y(n_4289)
);

OAI21x1_ASAP7_75t_L g4290 ( 
.A1(n_3842),
.A2(n_3286),
.B(n_3276),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_3542),
.B(n_3458),
.Y(n_4291)
);

INVx4_ASAP7_75t_L g4292 ( 
.A(n_3689),
.Y(n_4292)
);

AOI22xp33_ASAP7_75t_L g4293 ( 
.A1(n_3901),
.A2(n_3256),
.B1(n_3327),
.B2(n_3355),
.Y(n_4293)
);

OAI21x1_ASAP7_75t_L g4294 ( 
.A1(n_3842),
.A2(n_3289),
.B(n_3278),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3697),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_3885),
.A2(n_3273),
.B(n_3327),
.Y(n_4296)
);

INVx4_ASAP7_75t_L g4297 ( 
.A(n_3689),
.Y(n_4297)
);

AOI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_3754),
.A2(n_3355),
.B1(n_3327),
.B2(n_3239),
.Y(n_4298)
);

AOI22xp33_ASAP7_75t_L g4299 ( 
.A1(n_3901),
.A2(n_3256),
.B1(n_3327),
.B2(n_3355),
.Y(n_4299)
);

BUFx12f_ASAP7_75t_L g4300 ( 
.A(n_3514),
.Y(n_4300)
);

OAI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_3781),
.A2(n_3239),
.B(n_3355),
.Y(n_4301)
);

CKINVDCx20_ASAP7_75t_R g4302 ( 
.A(n_3622),
.Y(n_4302)
);

A2O1A1Ixp33_ASAP7_75t_L g4303 ( 
.A1(n_3591),
.A2(n_3239),
.B(n_3127),
.C(n_3137),
.Y(n_4303)
);

OR2x2_ASAP7_75t_L g4304 ( 
.A(n_3643),
.B(n_3137),
.Y(n_4304)
);

AND2x4_ASAP7_75t_L g4305 ( 
.A(n_3568),
.B(n_3458),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3703),
.Y(n_4306)
);

OAI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3781),
.A2(n_3804),
.B(n_3709),
.Y(n_4307)
);

NOR2xp67_ASAP7_75t_L g4308 ( 
.A(n_3842),
.B(n_3158),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_3514),
.Y(n_4309)
);

NAND2x1p5_ASAP7_75t_L g4310 ( 
.A(n_3633),
.B(n_3203),
.Y(n_4310)
);

AOI22xp33_ASAP7_75t_L g4311 ( 
.A1(n_3605),
.A2(n_3239),
.B1(n_3203),
.B2(n_3143),
.Y(n_4311)
);

NAND2x2_ASAP7_75t_L g4312 ( 
.A(n_3911),
.B(n_3108),
.Y(n_4312)
);

AOI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_3885),
.A2(n_3129),
.B(n_3118),
.Y(n_4313)
);

AO21x2_ASAP7_75t_L g4314 ( 
.A1(n_3641),
.A2(n_2978),
.B(n_3013),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3703),
.Y(n_4315)
);

AOI22xp33_ASAP7_75t_L g4316 ( 
.A1(n_3605),
.A2(n_3203),
.B1(n_3143),
.B2(n_3128),
.Y(n_4316)
);

OAI21x1_ASAP7_75t_L g4317 ( 
.A1(n_3861),
.A2(n_3908),
.B(n_3869),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3705),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_3816),
.B(n_3367),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3705),
.Y(n_4320)
);

AND2x4_ASAP7_75t_L g4321 ( 
.A(n_3568),
.B(n_3458),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_3825),
.B(n_3367),
.Y(n_4322)
);

HB1xp67_ASAP7_75t_L g4323 ( 
.A(n_3654),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3726),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3825),
.B(n_3349),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3726),
.Y(n_4326)
);

HB1xp67_ASAP7_75t_L g4327 ( 
.A(n_3723),
.Y(n_4327)
);

INVxp67_ASAP7_75t_SL g4328 ( 
.A(n_3789),
.Y(n_4328)
);

BUFx3_ASAP7_75t_L g4329 ( 
.A(n_3683),
.Y(n_4329)
);

OAI21x1_ASAP7_75t_SL g4330 ( 
.A1(n_3510),
.A2(n_3050),
.B(n_3290),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_3662),
.B(n_3367),
.Y(n_4331)
);

AO21x1_ASAP7_75t_L g4332 ( 
.A1(n_3927),
.A2(n_3367),
.B(n_3349),
.Y(n_4332)
);

OAI22xp33_ASAP7_75t_L g4333 ( 
.A1(n_3606),
.A2(n_3203),
.B1(n_3143),
.B2(n_3330),
.Y(n_4333)
);

BUFx12f_ASAP7_75t_L g4334 ( 
.A(n_3514),
.Y(n_4334)
);

AOI21x1_ASAP7_75t_L g4335 ( 
.A1(n_3719),
.A2(n_3151),
.B(n_3232),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_3838),
.B(n_3881),
.Y(n_4336)
);

INVx3_ASAP7_75t_L g4337 ( 
.A(n_3507),
.Y(n_4337)
);

AOI21xp5_ASAP7_75t_L g4338 ( 
.A1(n_3885),
.A2(n_3143),
.B(n_3248),
.Y(n_4338)
);

AO21x2_ASAP7_75t_L g4339 ( 
.A1(n_3641),
.A2(n_3160),
.B(n_3232),
.Y(n_4339)
);

HB1xp67_ASAP7_75t_L g4340 ( 
.A(n_3723),
.Y(n_4340)
);

CKINVDCx6p67_ASAP7_75t_R g4341 ( 
.A(n_3603),
.Y(n_4341)
);

OR2x2_ASAP7_75t_L g4342 ( 
.A(n_3515),
.B(n_3349),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_3730),
.Y(n_4343)
);

AOI21x1_ASAP7_75t_L g4344 ( 
.A1(n_3712),
.A2(n_3160),
.B(n_3243),
.Y(n_4344)
);

BUFx3_ASAP7_75t_L g4345 ( 
.A(n_3603),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3730),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_3554),
.B(n_3126),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_3542),
.B(n_3349),
.Y(n_4348)
);

OR2x2_ASAP7_75t_L g4349 ( 
.A(n_3515),
.B(n_3349),
.Y(n_4349)
);

OAI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_3606),
.A2(n_3330),
.B1(n_3310),
.B2(n_3265),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_3554),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_3713),
.A2(n_3330),
.B1(n_3310),
.B2(n_3165),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_3925),
.A2(n_3771),
.B(n_3766),
.Y(n_4353)
);

NOR2xp33_ASAP7_75t_L g4354 ( 
.A(n_3554),
.B(n_3165),
.Y(n_4354)
);

OAI22xp5_ASAP7_75t_L g4355 ( 
.A1(n_3591),
.A2(n_3330),
.B1(n_3310),
.B2(n_3165),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_3582),
.B(n_3330),
.Y(n_4356)
);

AOI21x1_ASAP7_75t_L g4357 ( 
.A1(n_3712),
.A2(n_3095),
.B(n_3250),
.Y(n_4357)
);

O2A1O1Ixp33_ASAP7_75t_SL g4358 ( 
.A1(n_3702),
.A2(n_3330),
.B(n_3310),
.C(n_3091),
.Y(n_4358)
);

CKINVDCx20_ASAP7_75t_R g4359 ( 
.A(n_3612),
.Y(n_4359)
);

A2O1A1Ixp33_ASAP7_75t_L g4360 ( 
.A1(n_3592),
.A2(n_3271),
.B(n_3265),
.C(n_3260),
.Y(n_4360)
);

AOI22xp5_ASAP7_75t_L g4361 ( 
.A1(n_3605),
.A2(n_3552),
.B1(n_3598),
.B2(n_3538),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_3582),
.B(n_3063),
.Y(n_4362)
);

AND2x6_ASAP7_75t_L g4363 ( 
.A(n_3620),
.B(n_3271),
.Y(n_4363)
);

O2A1O1Ixp33_ASAP7_75t_SL g4364 ( 
.A1(n_3742),
.A2(n_3260),
.B(n_3199),
.C(n_3113),
.Y(n_4364)
);

BUFx3_ASAP7_75t_L g4365 ( 
.A(n_3603),
.Y(n_4365)
);

OAI221xp5_ASAP7_75t_L g4366 ( 
.A1(n_3490),
.A2(n_3260),
.B1(n_3199),
.B2(n_3091),
.C(n_3063),
.Y(n_4366)
);

OAI21x1_ASAP7_75t_L g4367 ( 
.A1(n_3766),
.A2(n_3057),
.B(n_3063),
.Y(n_4367)
);

OA21x2_ASAP7_75t_L g4368 ( 
.A1(n_3812),
.A2(n_3063),
.B(n_3057),
.Y(n_4368)
);

OAI21x1_ASAP7_75t_L g4369 ( 
.A1(n_3771),
.A2(n_3057),
.B(n_3063),
.Y(n_4369)
);

INVxp67_ASAP7_75t_SL g4370 ( 
.A(n_3789),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_3838),
.B(n_3063),
.Y(n_4371)
);

BUFx3_ASAP7_75t_L g4372 ( 
.A(n_3617),
.Y(n_4372)
);

OAI21x1_ASAP7_75t_L g4373 ( 
.A1(n_3771),
.A2(n_3057),
.B(n_3078),
.Y(n_4373)
);

OAI21x1_ASAP7_75t_L g4374 ( 
.A1(n_3771),
.A2(n_3057),
.B(n_3078),
.Y(n_4374)
);

AOI22xp33_ASAP7_75t_L g4375 ( 
.A1(n_3552),
.A2(n_3078),
.B1(n_3057),
.B2(n_3185),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_3575),
.B(n_3078),
.Y(n_4376)
);

AND2x4_ASAP7_75t_L g4377 ( 
.A(n_3575),
.B(n_3080),
.Y(n_4377)
);

AO21x2_ASAP7_75t_L g4378 ( 
.A1(n_3751),
.A2(n_3080),
.B(n_3120),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_3582),
.B(n_3080),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_3599),
.B(n_3080),
.Y(n_4380)
);

OAI22xp33_ASAP7_75t_L g4381 ( 
.A1(n_3598),
.A2(n_3120),
.B1(n_3163),
.B2(n_3178),
.Y(n_4381)
);

OAI21x1_ASAP7_75t_L g4382 ( 
.A1(n_3692),
.A2(n_3120),
.B(n_3163),
.Y(n_4382)
);

AOI221xp5_ASAP7_75t_L g4383 ( 
.A1(n_3811),
.A2(n_3120),
.B1(n_3163),
.B2(n_3178),
.C(n_3185),
.Y(n_4383)
);

OAI21x1_ASAP7_75t_L g4384 ( 
.A1(n_3692),
.A2(n_3120),
.B(n_3163),
.Y(n_4384)
);

OAI21x1_ASAP7_75t_L g4385 ( 
.A1(n_3692),
.A2(n_3163),
.B(n_3178),
.Y(n_4385)
);

AO21x2_ASAP7_75t_L g4386 ( 
.A1(n_3761),
.A2(n_3163),
.B(n_3178),
.Y(n_4386)
);

BUFx3_ASAP7_75t_L g4387 ( 
.A(n_3617),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_3599),
.B(n_3178),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_L g4389 ( 
.A1(n_3552),
.A2(n_3185),
.B1(n_3462),
.B2(n_3465),
.Y(n_4389)
);

A2O1A1Ixp33_ASAP7_75t_L g4390 ( 
.A1(n_3592),
.A2(n_3185),
.B(n_3596),
.C(n_3911),
.Y(n_4390)
);

BUFx3_ASAP7_75t_L g4391 ( 
.A(n_3617),
.Y(n_4391)
);

NOR2xp33_ASAP7_75t_L g4392 ( 
.A(n_3612),
.B(n_3659),
.Y(n_4392)
);

OAI21x1_ASAP7_75t_L g4393 ( 
.A1(n_3692),
.A2(n_3694),
.B(n_3804),
.Y(n_4393)
);

AOI22xp33_ASAP7_75t_L g4394 ( 
.A1(n_3552),
.A2(n_3490),
.B1(n_3538),
.B2(n_3498),
.Y(n_4394)
);

INVxp67_ASAP7_75t_SL g4395 ( 
.A(n_3900),
.Y(n_4395)
);

OAI21x1_ASAP7_75t_L g4396 ( 
.A1(n_3694),
.A2(n_3804),
.B(n_3840),
.Y(n_4396)
);

OAI21x1_ASAP7_75t_L g4397 ( 
.A1(n_3694),
.A2(n_3804),
.B(n_3840),
.Y(n_4397)
);

OAI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_3687),
.A2(n_3709),
.B(n_3913),
.Y(n_4398)
);

OAI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_3592),
.A2(n_3596),
.B1(n_3490),
.B2(n_3913),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_3659),
.Y(n_4400)
);

INVx3_ASAP7_75t_SL g4401 ( 
.A(n_3689),
.Y(n_4401)
);

AOI21x1_ASAP7_75t_L g4402 ( 
.A1(n_3763),
.A2(n_3772),
.B(n_3768),
.Y(n_4402)
);

BUFx3_ASAP7_75t_L g4403 ( 
.A(n_3659),
.Y(n_4403)
);

OAI21x1_ASAP7_75t_L g4404 ( 
.A1(n_3694),
.A2(n_3840),
.B(n_3745),
.Y(n_4404)
);

AO21x2_ASAP7_75t_L g4405 ( 
.A1(n_3763),
.A2(n_3772),
.B(n_3768),
.Y(n_4405)
);

INVxp67_ASAP7_75t_L g4406 ( 
.A(n_3512),
.Y(n_4406)
);

BUFx8_ASAP7_75t_SL g4407 ( 
.A(n_3727),
.Y(n_4407)
);

OAI21x1_ASAP7_75t_L g4408 ( 
.A1(n_3840),
.A2(n_3745),
.B(n_3725),
.Y(n_4408)
);

AOI22x1_ASAP7_75t_L g4409 ( 
.A1(n_3811),
.A2(n_3693),
.B1(n_3710),
.B2(n_3690),
.Y(n_4409)
);

AO21x2_ASAP7_75t_L g4410 ( 
.A1(n_3768),
.A2(n_3776),
.B(n_3772),
.Y(n_4410)
);

CKINVDCx20_ASAP7_75t_R g4411 ( 
.A(n_3934),
.Y(n_4411)
);

O2A1O1Ixp33_ASAP7_75t_SL g4412 ( 
.A1(n_3742),
.A2(n_3743),
.B(n_3604),
.C(n_3506),
.Y(n_4412)
);

AOI21xp5_ASAP7_75t_L g4413 ( 
.A1(n_3866),
.A2(n_3922),
.B(n_3895),
.Y(n_4413)
);

AOI22xp5_ASAP7_75t_L g4414 ( 
.A1(n_3552),
.A2(n_3498),
.B1(n_3538),
.B2(n_3792),
.Y(n_4414)
);

INVx2_ASAP7_75t_SL g4415 ( 
.A(n_3536),
.Y(n_4415)
);

OAI21x1_ASAP7_75t_L g4416 ( 
.A1(n_3725),
.A2(n_3745),
.B(n_3511),
.Y(n_4416)
);

CKINVDCx11_ASAP7_75t_R g4417 ( 
.A(n_3756),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_3599),
.B(n_3618),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_3618),
.B(n_3647),
.Y(n_4419)
);

AO21x2_ASAP7_75t_L g4420 ( 
.A1(n_3776),
.A2(n_3794),
.B(n_3777),
.Y(n_4420)
);

BUFx3_ASAP7_75t_L g4421 ( 
.A(n_3536),
.Y(n_4421)
);

OAI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_3687),
.A2(n_3913),
.B(n_3538),
.Y(n_4422)
);

AOI21x1_ASAP7_75t_L g4423 ( 
.A1(n_3776),
.A2(n_3794),
.B(n_3777),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_L g4424 ( 
.A1(n_3725),
.A2(n_3745),
.B(n_3511),
.Y(n_4424)
);

HB1xp67_ASAP7_75t_L g4425 ( 
.A(n_3512),
.Y(n_4425)
);

INVx4_ASAP7_75t_L g4426 ( 
.A(n_3544),
.Y(n_4426)
);

OR2x2_ASAP7_75t_L g4427 ( 
.A(n_3515),
.B(n_3886),
.Y(n_4427)
);

AO21x2_ASAP7_75t_L g4428 ( 
.A1(n_3777),
.A2(n_3815),
.B(n_3794),
.Y(n_4428)
);

NAND2xp33_ASAP7_75t_R g4429 ( 
.A(n_3465),
.B(n_3668),
.Y(n_4429)
);

OAI21x1_ASAP7_75t_L g4430 ( 
.A1(n_3725),
.A2(n_3511),
.B(n_3507),
.Y(n_4430)
);

OAI22x1_ASAP7_75t_L g4431 ( 
.A1(n_3498),
.A2(n_3482),
.B1(n_3487),
.B2(n_3486),
.Y(n_4431)
);

OA21x2_ASAP7_75t_L g4432 ( 
.A1(n_3812),
.A2(n_3858),
.B(n_3836),
.Y(n_4432)
);

HB1xp67_ASAP7_75t_L g4433 ( 
.A(n_3537),
.Y(n_4433)
);

OAI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_3498),
.A2(n_3593),
.B(n_3589),
.Y(n_4434)
);

BUFx12f_ASAP7_75t_L g4435 ( 
.A(n_3808),
.Y(n_4435)
);

AO21x2_ASAP7_75t_L g4436 ( 
.A1(n_3815),
.A2(n_3821),
.B(n_3817),
.Y(n_4436)
);

BUFx2_ASAP7_75t_L g4437 ( 
.A(n_3686),
.Y(n_4437)
);

INVx4_ASAP7_75t_L g4438 ( 
.A(n_3544),
.Y(n_4438)
);

BUFx3_ASAP7_75t_L g4439 ( 
.A(n_3544),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_3626),
.Y(n_4440)
);

OAI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_3596),
.A2(n_3465),
.B1(n_3486),
.B2(n_3482),
.Y(n_4441)
);

OAI21x1_ASAP7_75t_L g4442 ( 
.A1(n_3619),
.A2(n_3630),
.B(n_3627),
.Y(n_4442)
);

OAI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_3618),
.A2(n_3729),
.B1(n_3735),
.B2(n_3647),
.Y(n_4443)
);

AOI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_3552),
.A2(n_3462),
.B1(n_3465),
.B2(n_3574),
.Y(n_4444)
);

AOI22x1_ASAP7_75t_L g4445 ( 
.A1(n_3690),
.A2(n_3693),
.B1(n_3717),
.B2(n_3710),
.Y(n_4445)
);

OA21x2_ASAP7_75t_L g4446 ( 
.A1(n_3812),
.A2(n_3858),
.B(n_3836),
.Y(n_4446)
);

BUFx8_ASAP7_75t_L g4447 ( 
.A(n_4435),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3937),
.Y(n_4448)
);

BUFx12f_ASAP7_75t_L g4449 ( 
.A(n_3962),
.Y(n_4449)
);

INVx6_ASAP7_75t_L g4450 ( 
.A(n_4056),
.Y(n_4450)
);

INVx2_ASAP7_75t_SL g4451 ( 
.A(n_4425),
.Y(n_4451)
);

BUFx2_ASAP7_75t_L g4452 ( 
.A(n_4069),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_3937),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4402),
.Y(n_4454)
);

HB1xp67_ASAP7_75t_L g4455 ( 
.A(n_4130),
.Y(n_4455)
);

OR2x2_ASAP7_75t_L g4456 ( 
.A(n_3957),
.B(n_3788),
.Y(n_4456)
);

AOI22xp33_ASAP7_75t_L g4457 ( 
.A1(n_3954),
.A2(n_3552),
.B1(n_3465),
.B2(n_3462),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4137),
.B(n_3743),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_4069),
.Y(n_4459)
);

INVx2_ASAP7_75t_L g4460 ( 
.A(n_4402),
.Y(n_4460)
);

BUFx12f_ASAP7_75t_L g4461 ( 
.A(n_4256),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_3943),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4423),
.Y(n_4463)
);

AOI222xp33_ASAP7_75t_L g4464 ( 
.A1(n_4059),
.A2(n_3734),
.B1(n_3736),
.B2(n_3932),
.C1(n_3905),
.C2(n_3886),
.Y(n_4464)
);

BUFx6f_ASAP7_75t_L g4465 ( 
.A(n_4093),
.Y(n_4465)
);

HB1xp67_ASAP7_75t_L g4466 ( 
.A(n_4130),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_3943),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4423),
.Y(n_4468)
);

CKINVDCx11_ASAP7_75t_R g4469 ( 
.A(n_4025),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_4004),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_3950),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4344),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4344),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4068),
.A2(n_3627),
.B(n_3619),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_4113),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4226),
.B(n_3647),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4357),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4357),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4209),
.Y(n_4479)
);

BUFx2_ASAP7_75t_L g4480 ( 
.A(n_4113),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4209),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4209),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3950),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_3951),
.Y(n_4484)
);

CKINVDCx20_ASAP7_75t_R g4485 ( 
.A(n_4117),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4209),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_3951),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_3959),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_3959),
.Y(n_4489)
);

AOI22xp33_ASAP7_75t_SL g4490 ( 
.A1(n_3941),
.A2(n_3552),
.B1(n_3482),
.B2(n_3487),
.Y(n_4490)
);

BUFx3_ASAP7_75t_L g4491 ( 
.A(n_4300),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_3960),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4137),
.B(n_3905),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_4093),
.Y(n_4494)
);

INVx3_ASAP7_75t_L g4495 ( 
.A(n_4432),
.Y(n_4495)
);

OAI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_3941),
.A2(n_3646),
.B1(n_3473),
.B2(n_3770),
.Y(n_4496)
);

OAI21x1_ASAP7_75t_L g4497 ( 
.A1(n_4068),
.A2(n_3627),
.B(n_3619),
.Y(n_4497)
);

CKINVDCx5p33_ASAP7_75t_R g4498 ( 
.A(n_4099),
.Y(n_4498)
);

AOI22xp33_ASAP7_75t_L g4499 ( 
.A1(n_3954),
.A2(n_3552),
.B1(n_3465),
.B2(n_3462),
.Y(n_4499)
);

HB1xp67_ASAP7_75t_L g4500 ( 
.A(n_4250),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_3960),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4405),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4405),
.Y(n_4503)
);

NAND2x1p5_ASAP7_75t_L g4504 ( 
.A(n_4273),
.B(n_3633),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_3969),
.Y(n_4505)
);

INVx3_ASAP7_75t_L g4506 ( 
.A(n_4432),
.Y(n_4506)
);

OR2x6_ASAP7_75t_L g4507 ( 
.A(n_4431),
.B(n_3574),
.Y(n_4507)
);

INVx6_ASAP7_75t_L g4508 ( 
.A(n_4056),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4405),
.Y(n_4509)
);

BUFx5_ASAP7_75t_L g4510 ( 
.A(n_4363),
.Y(n_4510)
);

BUFx6f_ASAP7_75t_L g4511 ( 
.A(n_4093),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4405),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_3969),
.Y(n_4513)
);

BUFx3_ASAP7_75t_L g4514 ( 
.A(n_4300),
.Y(n_4514)
);

AOI21x1_ASAP7_75t_L g4515 ( 
.A1(n_4078),
.A2(n_3508),
.B(n_3505),
.Y(n_4515)
);

BUFx2_ASAP7_75t_L g4516 ( 
.A(n_4328),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_4138),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_3971),
.Y(n_4518)
);

HB1xp67_ASAP7_75t_L g4519 ( 
.A(n_4250),
.Y(n_4519)
);

AOI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_3949),
.A2(n_3552),
.B1(n_3850),
.B2(n_3587),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4261),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_3971),
.Y(n_4522)
);

BUFx3_ASAP7_75t_L g4523 ( 
.A(n_4300),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4335),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3998),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3998),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4335),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4410),
.Y(n_4528)
);

BUFx3_ASAP7_75t_L g4529 ( 
.A(n_4334),
.Y(n_4529)
);

AOI22xp33_ASAP7_75t_SL g4530 ( 
.A1(n_3966),
.A2(n_3486),
.B1(n_3487),
.B2(n_3482),
.Y(n_4530)
);

INVx4_ASAP7_75t_L g4531 ( 
.A(n_3990),
.Y(n_4531)
);

A2O1A1Ixp33_ASAP7_75t_L g4532 ( 
.A1(n_4059),
.A2(n_3736),
.B(n_3734),
.C(n_3476),
.Y(n_4532)
);

INVx2_ASAP7_75t_SL g4533 ( 
.A(n_4425),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_SL g4534 ( 
.A1(n_3966),
.A2(n_3486),
.B1(n_3487),
.B2(n_3482),
.Y(n_4534)
);

INVx2_ASAP7_75t_SL g4535 ( 
.A(n_4433),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_3999),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3999),
.Y(n_4537)
);

INVxp67_ASAP7_75t_L g4538 ( 
.A(n_4007),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4226),
.B(n_3729),
.Y(n_4539)
);

AOI21x1_ASAP7_75t_L g4540 ( 
.A1(n_4078),
.A2(n_3508),
.B(n_3505),
.Y(n_4540)
);

INVx6_ASAP7_75t_L g4541 ( 
.A(n_4334),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4410),
.Y(n_4542)
);

HB1xp67_ASAP7_75t_L g4543 ( 
.A(n_4261),
.Y(n_4543)
);

NAND2x1p5_ASAP7_75t_L g4544 ( 
.A(n_4273),
.B(n_3482),
.Y(n_4544)
);

OR2x2_ASAP7_75t_L g4545 ( 
.A(n_3957),
.B(n_3788),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4410),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4410),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4000),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4000),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4001),
.Y(n_4550)
);

INVx3_ASAP7_75t_L g4551 ( 
.A(n_4432),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4420),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_4088),
.B(n_3932),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_4147),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4420),
.Y(n_4555)
);

INVx3_ASAP7_75t_L g4556 ( 
.A(n_4432),
.Y(n_4556)
);

AO21x1_ASAP7_75t_SL g4557 ( 
.A1(n_4123),
.A2(n_3847),
.B(n_3835),
.Y(n_4557)
);

AOI22xp33_ASAP7_75t_L g4558 ( 
.A1(n_4010),
.A2(n_3462),
.B1(n_3486),
.B2(n_3482),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4420),
.Y(n_4559)
);

BUFx4f_ASAP7_75t_SL g4560 ( 
.A(n_4302),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4088),
.B(n_3589),
.Y(n_4561)
);

AOI22xp33_ASAP7_75t_L g4562 ( 
.A1(n_4010),
.A2(n_3486),
.B1(n_3487),
.B2(n_3482),
.Y(n_4562)
);

INVx3_ASAP7_75t_L g4563 ( 
.A(n_4432),
.Y(n_4563)
);

INVx2_ASAP7_75t_L g4564 ( 
.A(n_4420),
.Y(n_4564)
);

INVx2_ASAP7_75t_SL g4565 ( 
.A(n_4433),
.Y(n_4565)
);

AO21x1_ASAP7_75t_L g4566 ( 
.A1(n_3973),
.A2(n_3682),
.B(n_3677),
.Y(n_4566)
);

AOI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_3970),
.A2(n_3487),
.B1(n_3488),
.B2(n_3486),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4001),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_4428),
.Y(n_4569)
);

INVxp67_ASAP7_75t_L g4570 ( 
.A(n_4212),
.Y(n_4570)
);

BUFx12f_ASAP7_75t_L g4571 ( 
.A(n_3956),
.Y(n_4571)
);

OAI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_3940),
.A2(n_3487),
.B1(n_3488),
.B2(n_3486),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4011),
.Y(n_4573)
);

HB1xp67_ASAP7_75t_L g4574 ( 
.A(n_4323),
.Y(n_4574)
);

OAI22xp33_ASAP7_75t_L g4575 ( 
.A1(n_3940),
.A2(n_3488),
.B1(n_3491),
.B2(n_3487),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4428),
.Y(n_4576)
);

INVx8_ASAP7_75t_L g4577 ( 
.A(n_4334),
.Y(n_4577)
);

OA21x2_ASAP7_75t_L g4578 ( 
.A1(n_4367),
.A2(n_4369),
.B(n_4353),
.Y(n_4578)
);

HB1xp67_ASAP7_75t_SL g4579 ( 
.A(n_4041),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4428),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4011),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4428),
.Y(n_4582)
);

BUFx2_ASAP7_75t_L g4583 ( 
.A(n_4328),
.Y(n_4583)
);

NAND2x1p5_ASAP7_75t_L g4584 ( 
.A(n_4030),
.B(n_3488),
.Y(n_4584)
);

AO21x1_ASAP7_75t_SL g4585 ( 
.A1(n_4123),
.A2(n_3847),
.B(n_3835),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4017),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4436),
.Y(n_4587)
);

HB1xp67_ASAP7_75t_L g4588 ( 
.A(n_4323),
.Y(n_4588)
);

INVx6_ASAP7_75t_L g4589 ( 
.A(n_4106),
.Y(n_4589)
);

BUFx3_ASAP7_75t_L g4590 ( 
.A(n_4435),
.Y(n_4590)
);

AOI22xp33_ASAP7_75t_L g4591 ( 
.A1(n_3970),
.A2(n_3491),
.B1(n_3525),
.B2(n_3488),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_4407),
.Y(n_4592)
);

BUFx4f_ASAP7_75t_SL g4593 ( 
.A(n_4411),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4017),
.Y(n_4594)
);

INVx3_ASAP7_75t_L g4595 ( 
.A(n_4446),
.Y(n_4595)
);

INVx3_ASAP7_75t_L g4596 ( 
.A(n_4446),
.Y(n_4596)
);

INVx1_ASAP7_75t_SL g4597 ( 
.A(n_4246),
.Y(n_4597)
);

OAI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_3949),
.A2(n_3955),
.B1(n_4005),
.B2(n_4047),
.Y(n_4598)
);

BUFx12f_ASAP7_75t_L g4599 ( 
.A(n_4417),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4018),
.Y(n_4600)
);

AND2x4_ASAP7_75t_L g4601 ( 
.A(n_3964),
.B(n_3876),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4436),
.Y(n_4602)
);

CKINVDCx20_ASAP7_75t_R g4603 ( 
.A(n_4205),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4018),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4024),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4024),
.Y(n_4606)
);

AND2x4_ASAP7_75t_L g4607 ( 
.A(n_3964),
.B(n_3876),
.Y(n_4607)
);

INVx2_ASAP7_75t_SL g4608 ( 
.A(n_4345),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4026),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4026),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4029),
.Y(n_4611)
);

INVx3_ASAP7_75t_L g4612 ( 
.A(n_4446),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4029),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4436),
.Y(n_4614)
);

HB1xp67_ASAP7_75t_L g4615 ( 
.A(n_4327),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4035),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4436),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4378),
.Y(n_4618)
);

OA21x2_ASAP7_75t_L g4619 ( 
.A1(n_4367),
.A2(n_3858),
.B(n_3836),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4327),
.Y(n_4620)
);

INVx3_ASAP7_75t_L g4621 ( 
.A(n_4446),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4035),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_4159),
.B(n_3876),
.Y(n_4623)
);

INVx3_ASAP7_75t_L g4624 ( 
.A(n_4446),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4127),
.Y(n_4625)
);

NAND2x1p5_ASAP7_75t_L g4626 ( 
.A(n_4030),
.B(n_3488),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_3957),
.B(n_3795),
.Y(n_4627)
);

INVxp67_ASAP7_75t_L g4628 ( 
.A(n_3936),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4127),
.Y(n_4629)
);

OR2x2_ASAP7_75t_L g4630 ( 
.A(n_4151),
.B(n_3795),
.Y(n_4630)
);

OAI22xp33_ASAP7_75t_L g4631 ( 
.A1(n_4082),
.A2(n_3491),
.B1(n_3525),
.B2(n_3488),
.Y(n_4631)
);

INVxp67_ASAP7_75t_L g4632 ( 
.A(n_3953),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4127),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4127),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4127),
.Y(n_4635)
);

BUFx4f_ASAP7_75t_SL g4636 ( 
.A(n_4359),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4043),
.Y(n_4637)
);

INVx3_ASAP7_75t_L g4638 ( 
.A(n_3965),
.Y(n_4638)
);

AOI22xp33_ASAP7_75t_L g4639 ( 
.A1(n_3944),
.A2(n_3491),
.B1(n_3525),
.B2(n_3488),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4043),
.Y(n_4640)
);

AOI22xp33_ASAP7_75t_L g4641 ( 
.A1(n_4023),
.A2(n_3525),
.B1(n_3491),
.B2(n_3574),
.Y(n_4641)
);

CKINVDCx20_ASAP7_75t_R g4642 ( 
.A(n_4022),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4107),
.B(n_3593),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4100),
.Y(n_4644)
);

AOI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4023),
.A2(n_3525),
.B1(n_3491),
.B2(n_3734),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4046),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4107),
.B(n_3594),
.Y(n_4647)
);

AOI22xp33_ASAP7_75t_SL g4648 ( 
.A1(n_3952),
.A2(n_3525),
.B1(n_3491),
.B2(n_3736),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4151),
.B(n_3677),
.Y(n_4649)
);

OR2x2_ASAP7_75t_L g4650 ( 
.A(n_4151),
.B(n_3682),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4046),
.Y(n_4651)
);

AOI22xp33_ASAP7_75t_L g4652 ( 
.A1(n_4047),
.A2(n_3525),
.B1(n_3491),
.B2(n_3575),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4378),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4378),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4378),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4049),
.Y(n_4656)
);

AOI22xp33_ASAP7_75t_L g4657 ( 
.A1(n_3975),
.A2(n_3525),
.B1(n_3584),
.B2(n_3587),
.Y(n_4657)
);

BUFx6f_ASAP7_75t_L g4658 ( 
.A(n_4100),
.Y(n_4658)
);

AOI22xp33_ASAP7_75t_L g4659 ( 
.A1(n_3975),
.A2(n_3584),
.B1(n_3587),
.B2(n_3904),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4226),
.B(n_3729),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4049),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4386),
.Y(n_4662)
);

AOI22xp33_ASAP7_75t_L g4663 ( 
.A1(n_3955),
.A2(n_3584),
.B1(n_3587),
.B2(n_3904),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_4340),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4057),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4057),
.Y(n_4666)
);

AOI22xp33_ASAP7_75t_SL g4667 ( 
.A1(n_3952),
.A2(n_3850),
.B1(n_3481),
.B2(n_3476),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4203),
.B(n_3594),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4386),
.Y(n_4669)
);

OAI22xp33_ASAP7_75t_L g4670 ( 
.A1(n_4082),
.A2(n_3587),
.B1(n_3566),
.B2(n_3476),
.Y(n_4670)
);

OAI22xp33_ASAP7_75t_L g4671 ( 
.A1(n_3952),
.A2(n_3587),
.B1(n_3566),
.B2(n_3481),
.Y(n_4671)
);

INVx3_ASAP7_75t_L g4672 ( 
.A(n_3965),
.Y(n_4672)
);

INVx8_ASAP7_75t_L g4673 ( 
.A(n_4435),
.Y(n_4673)
);

AOI22xp33_ASAP7_75t_L g4674 ( 
.A1(n_4055),
.A2(n_3904),
.B1(n_3481),
.B2(n_3624),
.Y(n_4674)
);

INVx2_ASAP7_75t_L g4675 ( 
.A(n_3938),
.Y(n_4675)
);

AOI21x1_ASAP7_75t_L g4676 ( 
.A1(n_4218),
.A2(n_3821),
.B(n_3817),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_L g4677 ( 
.A1(n_4055),
.A2(n_4005),
.B1(n_4074),
.B2(n_3987),
.Y(n_4677)
);

NAND2x1p5_ASAP7_75t_L g4678 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4061),
.Y(n_4679)
);

OAI22xp33_ASAP7_75t_L g4680 ( 
.A1(n_3952),
.A2(n_3566),
.B1(n_3473),
.B2(n_3626),
.Y(n_4680)
);

OAI22xp5_ASAP7_75t_L g4681 ( 
.A1(n_4040),
.A2(n_3473),
.B1(n_3798),
.B2(n_3770),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4061),
.Y(n_4682)
);

BUFx6f_ASAP7_75t_L g4683 ( 
.A(n_4100),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4203),
.B(n_3735),
.Y(n_4684)
);

OAI22xp5_ASAP7_75t_L g4685 ( 
.A1(n_4040),
.A2(n_3798),
.B1(n_3770),
.B2(n_3688),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4065),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_4340),
.Y(n_4687)
);

INVx4_ASAP7_75t_L g4688 ( 
.A(n_3990),
.Y(n_4688)
);

INVx3_ASAP7_75t_L g4689 ( 
.A(n_3965),
.Y(n_4689)
);

AOI21x1_ASAP7_75t_L g4690 ( 
.A1(n_4218),
.A2(n_3831),
.B(n_3830),
.Y(n_4690)
);

AOI22xp33_ASAP7_75t_L g4691 ( 
.A1(n_3987),
.A2(n_3904),
.B1(n_3624),
.B2(n_3878),
.Y(n_4691)
);

NAND2x1p5_ASAP7_75t_L g4692 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4692)
);

BUFx2_ASAP7_75t_L g4693 ( 
.A(n_4370),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_3938),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4065),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4070),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4070),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4386),
.Y(n_4698)
);

INVx4_ASAP7_75t_L g4699 ( 
.A(n_3990),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4156),
.B(n_3914),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4071),
.Y(n_4701)
);

HB1xp67_ASAP7_75t_L g4702 ( 
.A(n_4002),
.Y(n_4702)
);

OAI22xp5_ASAP7_75t_L g4703 ( 
.A1(n_4003),
.A2(n_3798),
.B1(n_3770),
.B2(n_3688),
.Y(n_4703)
);

BUFx8_ASAP7_75t_SL g4704 ( 
.A(n_4158),
.Y(n_4704)
);

INVx1_ASAP7_75t_SL g4705 ( 
.A(n_4014),
.Y(n_4705)
);

AOI22xp33_ASAP7_75t_L g4706 ( 
.A1(n_3972),
.A2(n_3904),
.B1(n_3624),
.B2(n_3878),
.Y(n_4706)
);

AOI22xp33_ASAP7_75t_SL g4707 ( 
.A1(n_3973),
.A2(n_3688),
.B1(n_3685),
.B2(n_3675),
.Y(n_4707)
);

BUFx4f_ASAP7_75t_SL g4708 ( 
.A(n_3967),
.Y(n_4708)
);

CKINVDCx11_ASAP7_75t_R g4709 ( 
.A(n_4014),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_3938),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4386),
.Y(n_4711)
);

AO21x1_ASAP7_75t_SL g4712 ( 
.A1(n_4143),
.A2(n_3862),
.B(n_3853),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4418),
.B(n_3735),
.Y(n_4713)
);

BUFx3_ASAP7_75t_L g4714 ( 
.A(n_3967),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4418),
.B(n_3737),
.Y(n_4715)
);

CKINVDCx20_ASAP7_75t_R g4716 ( 
.A(n_4038),
.Y(n_4716)
);

CKINVDCx20_ASAP7_75t_R g4717 ( 
.A(n_4038),
.Y(n_4717)
);

INVx4_ASAP7_75t_L g4718 ( 
.A(n_3980),
.Y(n_4718)
);

NAND2x1p5_ASAP7_75t_L g4719 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4719)
);

HB1xp67_ASAP7_75t_L g4720 ( 
.A(n_4002),
.Y(n_4720)
);

AOI22xp33_ASAP7_75t_L g4721 ( 
.A1(n_3972),
.A2(n_3624),
.B1(n_3878),
.B2(n_3560),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4071),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4314),
.Y(n_4723)
);

HB1xp67_ASAP7_75t_L g4724 ( 
.A(n_4037),
.Y(n_4724)
);

AO21x1_ASAP7_75t_L g4725 ( 
.A1(n_3982),
.A2(n_3862),
.B(n_3853),
.Y(n_4725)
);

OAI22xp33_ASAP7_75t_L g4726 ( 
.A1(n_3982),
.A2(n_3566),
.B1(n_3632),
.B2(n_3626),
.Y(n_4726)
);

AOI22xp5_ASAP7_75t_SL g4727 ( 
.A1(n_4225),
.A2(n_3638),
.B1(n_3645),
.B2(n_3632),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4314),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4084),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4084),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4036),
.B(n_4087),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4036),
.B(n_3737),
.Y(n_4732)
);

HB1xp67_ASAP7_75t_L g4733 ( 
.A(n_4037),
.Y(n_4733)
);

NOR2xp33_ASAP7_75t_SL g4734 ( 
.A(n_4066),
.B(n_3652),
.Y(n_4734)
);

NAND2x1p5_ASAP7_75t_L g4735 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4735)
);

INVx2_ASAP7_75t_SL g4736 ( 
.A(n_4345),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4314),
.Y(n_4737)
);

BUFx2_ASAP7_75t_L g4738 ( 
.A(n_4370),
.Y(n_4738)
);

BUFx6f_ASAP7_75t_L g4739 ( 
.A(n_4178),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4090),
.Y(n_4740)
);

OAI22xp5_ASAP7_75t_L g4741 ( 
.A1(n_3963),
.A2(n_3798),
.B1(n_3685),
.B2(n_3822),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4090),
.Y(n_4742)
);

INVx3_ASAP7_75t_L g4743 ( 
.A(n_3965),
.Y(n_4743)
);

INVx1_ASAP7_75t_SL g4744 ( 
.A(n_4066),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4418),
.B(n_3737),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4314),
.Y(n_4746)
);

AO21x2_ASAP7_75t_L g4747 ( 
.A1(n_4051),
.A2(n_3845),
.B(n_3844),
.Y(n_4747)
);

HB1xp67_ASAP7_75t_L g4748 ( 
.A(n_4406),
.Y(n_4748)
);

AOI21x1_ASAP7_75t_L g4749 ( 
.A1(n_4176),
.A2(n_3845),
.B(n_3844),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4091),
.Y(n_4750)
);

AOI22xp33_ASAP7_75t_L g4751 ( 
.A1(n_4122),
.A2(n_3624),
.B1(n_3878),
.B2(n_3560),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4091),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4097),
.Y(n_4753)
);

AOI22xp33_ASAP7_75t_L g4754 ( 
.A1(n_4122),
.A2(n_4352),
.B1(n_4019),
.B2(n_4072),
.Y(n_4754)
);

INVx8_ASAP7_75t_L g4755 ( 
.A(n_4204),
.Y(n_4755)
);

INVx4_ASAP7_75t_SL g4756 ( 
.A(n_3980),
.Y(n_4756)
);

INVx3_ASAP7_75t_L g4757 ( 
.A(n_3965),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4097),
.Y(n_4758)
);

OAI22xp33_ASAP7_75t_L g4759 ( 
.A1(n_4012),
.A2(n_3566),
.B1(n_3638),
.B2(n_3632),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4156),
.B(n_3914),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4339),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4103),
.Y(n_4762)
);

OAI22xp33_ASAP7_75t_L g4763 ( 
.A1(n_4012),
.A2(n_3566),
.B1(n_3645),
.B2(n_3638),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4103),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4339),
.Y(n_4765)
);

HB1xp67_ASAP7_75t_L g4766 ( 
.A(n_4406),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4116),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4339),
.Y(n_4768)
);

HB1xp67_ASAP7_75t_L g4769 ( 
.A(n_4044),
.Y(n_4769)
);

BUFx6f_ASAP7_75t_L g4770 ( 
.A(n_4178),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4116),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4126),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4126),
.Y(n_4773)
);

HB1xp67_ASAP7_75t_L g4774 ( 
.A(n_4044),
.Y(n_4774)
);

BUFx6f_ASAP7_75t_L g4775 ( 
.A(n_4178),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4339),
.Y(n_4776)
);

HB1xp67_ASAP7_75t_L g4777 ( 
.A(n_4081),
.Y(n_4777)
);

BUFx6f_ASAP7_75t_L g4778 ( 
.A(n_4180),
.Y(n_4778)
);

AOI21x1_ASAP7_75t_L g4779 ( 
.A1(n_4176),
.A2(n_3857),
.B(n_3852),
.Y(n_4779)
);

INVx1_ASAP7_75t_SL g4780 ( 
.A(n_4162),
.Y(n_4780)
);

NAND2x1p5_ASAP7_75t_L g4781 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4781)
);

BUFx2_ASAP7_75t_R g4782 ( 
.A(n_4206),
.Y(n_4782)
);

BUFx6f_ASAP7_75t_L g4783 ( 
.A(n_4180),
.Y(n_4783)
);

BUFx4f_ASAP7_75t_SL g4784 ( 
.A(n_3967),
.Y(n_4784)
);

AOI22xp33_ASAP7_75t_L g4785 ( 
.A1(n_4352),
.A2(n_4072),
.B1(n_4132),
.B2(n_4165),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4129),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4419),
.B(n_3758),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4156),
.B(n_3914),
.Y(n_4788)
);

BUFx6f_ASAP7_75t_L g4789 ( 
.A(n_4180),
.Y(n_4789)
);

OR2x2_ASAP7_75t_L g4790 ( 
.A(n_4167),
.B(n_3706),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4129),
.Y(n_4791)
);

INVx6_ASAP7_75t_L g4792 ( 
.A(n_4106),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4131),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4131),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4135),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_3948),
.Y(n_4796)
);

AOI22xp33_ASAP7_75t_SL g4797 ( 
.A1(n_4225),
.A2(n_3685),
.B1(n_3675),
.B2(n_3895),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4419),
.B(n_3758),
.Y(n_4798)
);

CKINVDCx5p33_ASAP7_75t_R g4799 ( 
.A(n_4253),
.Y(n_4799)
);

AO21x1_ASAP7_75t_SL g4800 ( 
.A1(n_4143),
.A2(n_3873),
.B(n_3863),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4135),
.Y(n_4801)
);

BUFx3_ASAP7_75t_L g4802 ( 
.A(n_3991),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4141),
.Y(n_4803)
);

OAI22xp5_ASAP7_75t_L g4804 ( 
.A1(n_3963),
.A2(n_3798),
.B1(n_3834),
.B2(n_3822),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4141),
.Y(n_4805)
);

NAND2x1p5_ASAP7_75t_L g4806 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_3948),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_SL g4808 ( 
.A(n_4102),
.B(n_3876),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_SL g4809 ( 
.A1(n_4108),
.A2(n_3517),
.B(n_3489),
.Y(n_4809)
);

AOI22xp33_ASAP7_75t_L g4810 ( 
.A1(n_4132),
.A2(n_4165),
.B1(n_4251),
.B2(n_4179),
.Y(n_4810)
);

HB1xp67_ASAP7_75t_L g4811 ( 
.A(n_4081),
.Y(n_4811)
);

OAI22xp33_ASAP7_75t_L g4812 ( 
.A1(n_4199),
.A2(n_3645),
.B1(n_3655),
.B2(n_3650),
.Y(n_4812)
);

HB1xp67_ASAP7_75t_L g4813 ( 
.A(n_4109),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_3948),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4142),
.Y(n_4815)
);

INVx2_ASAP7_75t_SL g4816 ( 
.A(n_4345),
.Y(n_4816)
);

AOI22xp5_ASAP7_75t_L g4817 ( 
.A1(n_4052),
.A2(n_3878),
.B1(n_3731),
.B2(n_3889),
.Y(n_4817)
);

BUFx6f_ASAP7_75t_L g4818 ( 
.A(n_4196),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4087),
.B(n_3758),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_4309),
.Y(n_4820)
);

AND2x2_ASAP7_75t_L g4821 ( 
.A(n_4419),
.B(n_3872),
.Y(n_4821)
);

OAI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4199),
.A2(n_3655),
.B1(n_3665),
.B2(n_3650),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4142),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4149),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4149),
.Y(n_4825)
);

HB1xp67_ASAP7_75t_L g4826 ( 
.A(n_4109),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4382),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4150),
.Y(n_4828)
);

BUFx2_ASAP7_75t_L g4829 ( 
.A(n_4421),
.Y(n_4829)
);

AOI22xp33_ASAP7_75t_SL g4830 ( 
.A1(n_4177),
.A2(n_4167),
.B1(n_4234),
.B2(n_4200),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4382),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4150),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4157),
.Y(n_4833)
);

BUFx2_ASAP7_75t_L g4834 ( 
.A(n_4421),
.Y(n_4834)
);

AOI22xp33_ASAP7_75t_L g4835 ( 
.A1(n_4251),
.A2(n_3624),
.B1(n_3560),
.B2(n_3558),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4382),
.Y(n_4836)
);

AOI21x1_ASAP7_75t_L g4837 ( 
.A1(n_4413),
.A2(n_4105),
.B(n_4243),
.Y(n_4837)
);

AOI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4179),
.A2(n_4332),
.B1(n_4124),
.B2(n_4051),
.Y(n_4838)
);

AOI21xp33_ASAP7_75t_L g4839 ( 
.A1(n_4027),
.A2(n_3807),
.B(n_3648),
.Y(n_4839)
);

AOI21x1_ASAP7_75t_L g4840 ( 
.A1(n_4413),
.A2(n_3857),
.B(n_3852),
.Y(n_4840)
);

AOI22xp5_ASAP7_75t_L g4841 ( 
.A1(n_4016),
.A2(n_4124),
.B1(n_3968),
.B2(n_4190),
.Y(n_4841)
);

BUFx2_ASAP7_75t_SL g4842 ( 
.A(n_3991),
.Y(n_4842)
);

AOI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_4190),
.A2(n_3731),
.B1(n_3891),
.B2(n_3889),
.Y(n_4843)
);

AOI22xp5_ASAP7_75t_L g4844 ( 
.A1(n_4177),
.A2(n_3731),
.B1(n_3891),
.B2(n_3889),
.Y(n_4844)
);

AOI22xp33_ASAP7_75t_SL g4845 ( 
.A1(n_4167),
.A2(n_3895),
.B1(n_3839),
.B2(n_3843),
.Y(n_4845)
);

AOI22xp33_ASAP7_75t_L g4846 ( 
.A1(n_4332),
.A2(n_3624),
.B1(n_3560),
.B2(n_3558),
.Y(n_4846)
);

AOI21x1_ASAP7_75t_L g4847 ( 
.A1(n_4105),
.A2(n_3877),
.B(n_3871),
.Y(n_4847)
);

AOI21x1_ASAP7_75t_L g4848 ( 
.A1(n_4243),
.A2(n_3877),
.B(n_3871),
.Y(n_4848)
);

OAI22xp5_ASAP7_75t_L g4849 ( 
.A1(n_4042),
.A2(n_3834),
.B1(n_3822),
.B2(n_3652),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_3995),
.B(n_3706),
.Y(n_4850)
);

INVx3_ASAP7_75t_L g4851 ( 
.A(n_3965),
.Y(n_4851)
);

AOI22xp33_ASAP7_75t_L g4852 ( 
.A1(n_4332),
.A2(n_3624),
.B1(n_3560),
.B2(n_3558),
.Y(n_4852)
);

NAND2x1p5_ASAP7_75t_L g4853 ( 
.A(n_4247),
.B(n_3887),
.Y(n_4853)
);

BUFx6f_ASAP7_75t_L g4854 ( 
.A(n_4196),
.Y(n_4854)
);

AOI22xp33_ASAP7_75t_SL g4855 ( 
.A1(n_4234),
.A2(n_3895),
.B1(n_3839),
.B2(n_3843),
.Y(n_4855)
);

BUFx2_ASAP7_75t_L g4856 ( 
.A(n_4421),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4384),
.Y(n_4857)
);

AOI22xp5_ASAP7_75t_L g4858 ( 
.A1(n_4042),
.A2(n_3731),
.B1(n_3902),
.B2(n_3891),
.Y(n_4858)
);

OAI22xp5_ASAP7_75t_L g4859 ( 
.A1(n_4217),
.A2(n_3834),
.B1(n_3670),
.B2(n_3676),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4157),
.Y(n_4860)
);

OA21x2_ASAP7_75t_L g4861 ( 
.A1(n_4367),
.A2(n_3922),
.B(n_3866),
.Y(n_4861)
);

BUFx6f_ASAP7_75t_L g4862 ( 
.A(n_4196),
.Y(n_4862)
);

AOI22xp33_ASAP7_75t_L g4863 ( 
.A1(n_4175),
.A2(n_3624),
.B1(n_3558),
.B2(n_3919),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4166),
.Y(n_4864)
);

OAI22xp33_ASAP7_75t_L g4865 ( 
.A1(n_4217),
.A2(n_3655),
.B1(n_3665),
.B2(n_3650),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4166),
.Y(n_4866)
);

HB1xp67_ASAP7_75t_L g4867 ( 
.A(n_4219),
.Y(n_4867)
);

AOI21x1_ASAP7_75t_L g4868 ( 
.A1(n_4169),
.A2(n_3893),
.B(n_3888),
.Y(n_4868)
);

CKINVDCx20_ASAP7_75t_R g4869 ( 
.A(n_4351),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4168),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4168),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4170),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4170),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4174),
.Y(n_4874)
);

AOI22xp33_ASAP7_75t_L g4875 ( 
.A1(n_4305),
.A2(n_3624),
.B1(n_3558),
.B2(n_3919),
.Y(n_4875)
);

AOI22x1_ASAP7_75t_L g4876 ( 
.A1(n_3980),
.A2(n_3898),
.B1(n_3541),
.B2(n_3556),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4174),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4181),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4181),
.Y(n_4879)
);

HB1xp67_ASAP7_75t_L g4880 ( 
.A(n_4219),
.Y(n_4880)
);

AO21x2_ASAP7_75t_L g4881 ( 
.A1(n_4039),
.A2(n_3893),
.B(n_3888),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4384),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4184),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4184),
.Y(n_4884)
);

OA21x2_ASAP7_75t_L g4885 ( 
.A1(n_4369),
.A2(n_3922),
.B(n_3866),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_3988),
.Y(n_4886)
);

OAI22xp5_ASAP7_75t_L g4887 ( 
.A1(n_3939),
.A2(n_3670),
.B1(n_3676),
.B2(n_3649),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4187),
.Y(n_4888)
);

AND2x2_ASAP7_75t_L g4889 ( 
.A(n_4200),
.B(n_3872),
.Y(n_4889)
);

INVx1_ASAP7_75t_SL g4890 ( 
.A(n_4195),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_SL g4891 ( 
.A1(n_4200),
.A2(n_3895),
.B1(n_3839),
.B2(n_3843),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4234),
.B(n_3872),
.Y(n_4892)
);

INVx1_ASAP7_75t_SL g4893 ( 
.A(n_4195),
.Y(n_4893)
);

AOI22xp33_ASAP7_75t_L g4894 ( 
.A1(n_4305),
.A2(n_3624),
.B1(n_3919),
.B2(n_3918),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4187),
.Y(n_4895)
);

OAI21x1_ASAP7_75t_L g4896 ( 
.A1(n_4140),
.A2(n_3894),
.B(n_3718),
.Y(n_4896)
);

BUFx6f_ASAP7_75t_L g4897 ( 
.A(n_4202),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4235),
.B(n_3711),
.Y(n_4898)
);

BUFx2_ASAP7_75t_SL g4899 ( 
.A(n_3991),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_4384),
.Y(n_4900)
);

OA21x2_ASAP7_75t_L g4901 ( 
.A1(n_4369),
.A2(n_3894),
.B(n_3807),
.Y(n_4901)
);

OAI22xp33_ASAP7_75t_L g4902 ( 
.A1(n_4201),
.A2(n_3681),
.B1(n_3665),
.B2(n_3902),
.Y(n_4902)
);

AOI22xp33_ASAP7_75t_L g4903 ( 
.A1(n_4305),
.A2(n_3919),
.B1(n_3918),
.B2(n_3917),
.Y(n_4903)
);

HB1xp67_ASAP7_75t_L g4904 ( 
.A(n_3988),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4193),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4193),
.Y(n_4906)
);

INVx1_ASAP7_75t_SL g4907 ( 
.A(n_4211),
.Y(n_4907)
);

OR2x2_ASAP7_75t_L g4908 ( 
.A(n_4235),
.B(n_3711),
.Y(n_4908)
);

INVx6_ASAP7_75t_L g4909 ( 
.A(n_4106),
.Y(n_4909)
);

CKINVDCx20_ASAP7_75t_R g4910 ( 
.A(n_4224),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4159),
.B(n_3876),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4197),
.Y(n_4912)
);

BUFx3_ASAP7_75t_L g4913 ( 
.A(n_4006),
.Y(n_4913)
);

OA21x2_ASAP7_75t_L g4914 ( 
.A1(n_4317),
.A2(n_3894),
.B(n_3807),
.Y(n_4914)
);

AO21x2_ASAP7_75t_L g4915 ( 
.A1(n_4039),
.A2(n_3785),
.B(n_3784),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4197),
.Y(n_4916)
);

OAI22xp5_ASAP7_75t_L g4917 ( 
.A1(n_3939),
.A2(n_3670),
.B1(n_3676),
.B2(n_3649),
.Y(n_4917)
);

OA21x2_ASAP7_75t_L g4918 ( 
.A1(n_4317),
.A2(n_3744),
.B(n_3740),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4385),
.Y(n_4919)
);

OAI21x1_ASAP7_75t_L g4920 ( 
.A1(n_4140),
.A2(n_3718),
.B(n_3701),
.Y(n_4920)
);

BUFx3_ASAP7_75t_L g4921 ( 
.A(n_4006),
.Y(n_4921)
);

INVx5_ASAP7_75t_L g4922 ( 
.A(n_4188),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4198),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_3995),
.B(n_3716),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4198),
.Y(n_4925)
);

INVx4_ASAP7_75t_L g4926 ( 
.A(n_4224),
.Y(n_4926)
);

AND2x2_ASAP7_75t_L g4927 ( 
.A(n_4235),
.B(n_3923),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4305),
.A2(n_3919),
.B1(n_3918),
.B2(n_3917),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4385),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4379),
.B(n_3923),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4214),
.Y(n_4931)
);

AND2x2_ASAP7_75t_L g4932 ( 
.A(n_4379),
.B(n_4380),
.Y(n_4932)
);

NOR2x1_ASAP7_75t_R g4933 ( 
.A(n_4006),
.B(n_3690),
.Y(n_4933)
);

AOI22xp33_ASAP7_75t_L g4934 ( 
.A1(n_4305),
.A2(n_3918),
.B1(n_3917),
.B2(n_3902),
.Y(n_4934)
);

AND2x2_ASAP7_75t_L g4935 ( 
.A(n_4379),
.B(n_3923),
.Y(n_4935)
);

INVx4_ASAP7_75t_L g4936 ( 
.A(n_4224),
.Y(n_4936)
);

INVx8_ASAP7_75t_L g4937 ( 
.A(n_4204),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4214),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4380),
.B(n_3923),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4020),
.B(n_3716),
.Y(n_4940)
);

INVx3_ASAP7_75t_L g4941 ( 
.A(n_3965),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4216),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_SL g4943 ( 
.A(n_4102),
.B(n_3668),
.Y(n_4943)
);

HB1xp67_ASAP7_75t_L g4944 ( 
.A(n_4211),
.Y(n_4944)
);

AOI22xp5_ASAP7_75t_L g4945 ( 
.A1(n_4080),
.A2(n_3731),
.B1(n_3926),
.B2(n_3924),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4385),
.Y(n_4946)
);

AOI22xp33_ASAP7_75t_L g4947 ( 
.A1(n_4321),
.A2(n_3918),
.B1(n_3926),
.B2(n_3924),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4216),
.Y(n_4948)
);

AND2x2_ASAP7_75t_L g4949 ( 
.A(n_4380),
.B(n_3923),
.Y(n_4949)
);

NAND2x1p5_ASAP7_75t_L g4950 ( 
.A(n_4442),
.B(n_3887),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_3978),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4227),
.Y(n_4952)
);

AOI21x1_ASAP7_75t_L g4953 ( 
.A1(n_4169),
.A2(n_3814),
.B(n_3806),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4227),
.Y(n_4954)
);

OAI22xp33_ASAP7_75t_L g4955 ( 
.A1(n_4201),
.A2(n_3681),
.B1(n_3926),
.B2(n_3924),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4229),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4229),
.Y(n_4957)
);

HB1xp67_ASAP7_75t_L g4958 ( 
.A(n_4194),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4236),
.Y(n_4959)
);

INVx1_ASAP7_75t_SL g4960 ( 
.A(n_4110),
.Y(n_4960)
);

NOR2xp33_ASAP7_75t_L g4961 ( 
.A(n_3947),
.B(n_3724),
.Y(n_4961)
);

NAND2x1p5_ASAP7_75t_L g4962 ( 
.A(n_4442),
.B(n_3912),
.Y(n_4962)
);

BUFx2_ASAP7_75t_R g4963 ( 
.A(n_4202),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4020),
.B(n_3724),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4236),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4252),
.Y(n_4966)
);

INVxp67_ASAP7_75t_L g4967 ( 
.A(n_4054),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4252),
.Y(n_4968)
);

OAI21xp5_ASAP7_75t_L g4969 ( 
.A1(n_4032),
.A2(n_3579),
.B(n_3555),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4257),
.Y(n_4970)
);

OAI22xp5_ASAP7_75t_L g4971 ( 
.A1(n_4058),
.A2(n_3670),
.B1(n_3676),
.B2(n_3649),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4388),
.B(n_4362),
.Y(n_4972)
);

AOI22xp33_ASAP7_75t_L g4973 ( 
.A1(n_4321),
.A2(n_3930),
.B1(n_3935),
.B2(n_3928),
.Y(n_4973)
);

INVx2_ASAP7_75t_SL g4974 ( 
.A(n_4365),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4257),
.Y(n_4975)
);

BUFx2_ASAP7_75t_L g4976 ( 
.A(n_4439),
.Y(n_4976)
);

BUFx2_ASAP7_75t_L g4977 ( 
.A(n_4439),
.Y(n_4977)
);

CKINVDCx16_ASAP7_75t_R g4978 ( 
.A(n_3979),
.Y(n_4978)
);

CKINVDCx11_ASAP7_75t_R g4979 ( 
.A(n_4341),
.Y(n_4979)
);

BUFx3_ASAP7_75t_L g4980 ( 
.A(n_4028),
.Y(n_4980)
);

BUFx6f_ASAP7_75t_L g4981 ( 
.A(n_4202),
.Y(n_4981)
);

AO21x1_ASAP7_75t_SL g4982 ( 
.A1(n_4155),
.A2(n_3873),
.B(n_3863),
.Y(n_4982)
);

OAI21xp5_ASAP7_75t_L g4983 ( 
.A1(n_4027),
.A2(n_3579),
.B(n_3555),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_L g4984 ( 
.A1(n_4321),
.A2(n_3930),
.B1(n_3935),
.B2(n_3928),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4260),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4260),
.Y(n_4986)
);

INVx2_ASAP7_75t_SL g4987 ( 
.A(n_4365),
.Y(n_4987)
);

INVx6_ASAP7_75t_L g4988 ( 
.A(n_4106),
.Y(n_4988)
);

AO21x1_ASAP7_75t_L g4989 ( 
.A1(n_3946),
.A2(n_3880),
.B(n_3874),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_3993),
.Y(n_4990)
);

BUFx3_ASAP7_75t_L g4991 ( 
.A(n_4028),
.Y(n_4991)
);

CKINVDCx5p33_ASAP7_75t_R g4992 ( 
.A(n_3947),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4062),
.A2(n_3684),
.B(n_3637),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4262),
.Y(n_4994)
);

INVx5_ASAP7_75t_L g4995 ( 
.A(n_4188),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_3993),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4262),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4264),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4264),
.Y(n_4999)
);

INVx6_ASAP7_75t_L g5000 ( 
.A(n_4242),
.Y(n_5000)
);

OAI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_4067),
.A2(n_3684),
.B(n_3637),
.Y(n_5001)
);

OR2x2_ASAP7_75t_L g5002 ( 
.A(n_4443),
.B(n_3733),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4265),
.Y(n_5003)
);

AOI21x1_ASAP7_75t_L g5004 ( 
.A1(n_3946),
.A2(n_3814),
.B(n_3806),
.Y(n_5004)
);

OAI21x1_ASAP7_75t_L g5005 ( 
.A1(n_4146),
.A2(n_3718),
.B(n_3701),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4265),
.Y(n_5006)
);

INVx3_ASAP7_75t_L g5007 ( 
.A(n_3976),
.Y(n_5007)
);

AOI22xp33_ASAP7_75t_L g5008 ( 
.A1(n_4321),
.A2(n_3930),
.B1(n_3935),
.B2(n_3928),
.Y(n_5008)
);

AOI21x1_ASAP7_75t_L g5009 ( 
.A1(n_3989),
.A2(n_3837),
.B(n_3823),
.Y(n_5009)
);

BUFx12f_ASAP7_75t_L g5010 ( 
.A(n_4028),
.Y(n_5010)
);

OAI21x1_ASAP7_75t_L g5011 ( 
.A1(n_4146),
.A2(n_3718),
.B(n_3701),
.Y(n_5011)
);

AOI21x1_ASAP7_75t_L g5012 ( 
.A1(n_3989),
.A2(n_3837),
.B(n_3823),
.Y(n_5012)
);

HB1xp67_ASAP7_75t_L g5013 ( 
.A(n_4194),
.Y(n_5013)
);

BUFx2_ASAP7_75t_SL g5014 ( 
.A(n_4050),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4272),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4272),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4279),
.Y(n_5017)
);

CKINVDCx11_ASAP7_75t_R g5018 ( 
.A(n_4341),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4279),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4282),
.Y(n_5020)
);

CKINVDCx5p33_ASAP7_75t_R g5021 ( 
.A(n_4050),
.Y(n_5021)
);

OAI22xp5_ASAP7_75t_L g5022 ( 
.A1(n_4058),
.A2(n_3670),
.B1(n_3676),
.B2(n_3649),
.Y(n_5022)
);

INVx2_ASAP7_75t_L g5023 ( 
.A(n_3996),
.Y(n_5023)
);

OAI21x1_ASAP7_75t_L g5024 ( 
.A1(n_4146),
.A2(n_3722),
.B(n_3701),
.Y(n_5024)
);

BUFx2_ASAP7_75t_L g5025 ( 
.A(n_4439),
.Y(n_5025)
);

AND2x2_ASAP7_75t_L g5026 ( 
.A(n_4388),
.B(n_3783),
.Y(n_5026)
);

OA21x2_ASAP7_75t_L g5027 ( 
.A1(n_4317),
.A2(n_3744),
.B(n_3740),
.Y(n_5027)
);

HB1xp67_ASAP7_75t_L g5028 ( 
.A(n_4194),
.Y(n_5028)
);

CKINVDCx20_ASAP7_75t_R g5029 ( 
.A(n_4341),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4172),
.B(n_3733),
.Y(n_5030)
);

BUFx2_ASAP7_75t_L g5031 ( 
.A(n_4060),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4295),
.Y(n_5032)
);

INVx8_ASAP7_75t_L g5033 ( 
.A(n_4204),
.Y(n_5033)
);

INVx6_ASAP7_75t_L g5034 ( 
.A(n_4242),
.Y(n_5034)
);

AOI22xp33_ASAP7_75t_L g5035 ( 
.A1(n_4321),
.A2(n_3681),
.B1(n_3620),
.B2(n_3739),
.Y(n_5035)
);

AOI22xp33_ASAP7_75t_L g5036 ( 
.A1(n_4285),
.A2(n_4350),
.B1(n_4376),
.B2(n_4355),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4295),
.Y(n_5037)
);

AOI22xp33_ASAP7_75t_SL g5038 ( 
.A1(n_4366),
.A2(n_4355),
.B1(n_4285),
.B2(n_4362),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4306),
.Y(n_5039)
);

AOI22xp5_ASAP7_75t_L g5040 ( 
.A1(n_4232),
.A2(n_3715),
.B1(n_3714),
.B2(n_3773),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4306),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4315),
.Y(n_5042)
);

NAND2x1p5_ASAP7_75t_L g5043 ( 
.A(n_4442),
.B(n_3912),
.Y(n_5043)
);

INVx8_ASAP7_75t_L g5044 ( 
.A(n_4204),
.Y(n_5044)
);

CKINVDCx5p33_ASAP7_75t_R g5045 ( 
.A(n_4050),
.Y(n_5045)
);

INVx6_ASAP7_75t_L g5046 ( 
.A(n_4242),
.Y(n_5046)
);

INVx4_ASAP7_75t_L g5047 ( 
.A(n_4185),
.Y(n_5047)
);

BUFx3_ASAP7_75t_L g5048 ( 
.A(n_4063),
.Y(n_5048)
);

CKINVDCx6p67_ASAP7_75t_R g5049 ( 
.A(n_4063),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4318),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4318),
.Y(n_5051)
);

BUFx10_ASAP7_75t_L g5052 ( 
.A(n_4392),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4320),
.Y(n_5053)
);

BUFx2_ASAP7_75t_SL g5054 ( 
.A(n_4063),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4008),
.Y(n_5055)
);

BUFx6f_ASAP7_75t_L g5056 ( 
.A(n_4329),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_4008),
.Y(n_5057)
);

INVx3_ASAP7_75t_L g5058 ( 
.A(n_3976),
.Y(n_5058)
);

AOI22xp5_ASAP7_75t_L g5059 ( 
.A1(n_4232),
.A2(n_3715),
.B1(n_3714),
.B2(n_3773),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_4060),
.Y(n_5060)
);

AOI22xp33_ASAP7_75t_L g5061 ( 
.A1(n_4285),
.A2(n_3620),
.B1(n_3739),
.B2(n_3648),
.Y(n_5061)
);

CKINVDCx5p33_ASAP7_75t_R g5062 ( 
.A(n_4077),
.Y(n_5062)
);

AOI22xp33_ASAP7_75t_L g5063 ( 
.A1(n_4285),
.A2(n_3620),
.B1(n_3739),
.B2(n_3648),
.Y(n_5063)
);

BUFx6f_ASAP7_75t_L g5064 ( 
.A(n_4329),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4320),
.Y(n_5065)
);

AOI22xp33_ASAP7_75t_SL g5066 ( 
.A1(n_4366),
.A2(n_3895),
.B1(n_3839),
.B2(n_3843),
.Y(n_5066)
);

INVx6_ASAP7_75t_L g5067 ( 
.A(n_4242),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4388),
.B(n_3783),
.Y(n_5068)
);

BUFx6f_ASAP7_75t_L g5069 ( 
.A(n_4329),
.Y(n_5069)
);

AOI22xp33_ASAP7_75t_SL g5070 ( 
.A1(n_4285),
.A2(n_4362),
.B1(n_4288),
.B2(n_4348),
.Y(n_5070)
);

AOI22xp33_ASAP7_75t_L g5071 ( 
.A1(n_4350),
.A2(n_3620),
.B1(n_3648),
.B2(n_3635),
.Y(n_5071)
);

AOI22xp33_ASAP7_75t_L g5072 ( 
.A1(n_4376),
.A2(n_3620),
.B1(n_3648),
.B2(n_3635),
.Y(n_5072)
);

OA21x2_ASAP7_75t_L g5073 ( 
.A1(n_4353),
.A2(n_3854),
.B(n_3846),
.Y(n_5073)
);

AND2x4_ASAP7_75t_L g5074 ( 
.A(n_4159),
.B(n_3625),
.Y(n_5074)
);

CKINVDCx11_ASAP7_75t_R g5075 ( 
.A(n_4185),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4324),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4008),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_4077),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4324),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_SL g5080 ( 
.A1(n_4288),
.A2(n_3843),
.B1(n_3839),
.B2(n_3565),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_4077),
.Y(n_5081)
);

INVx2_ASAP7_75t_L g5082 ( 
.A(n_4009),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4326),
.Y(n_5083)
);

INVx2_ASAP7_75t_L g5084 ( 
.A(n_4009),
.Y(n_5084)
);

HB1xp67_ASAP7_75t_L g5085 ( 
.A(n_4194),
.Y(n_5085)
);

INVx1_ASAP7_75t_SL g5086 ( 
.A(n_4266),
.Y(n_5086)
);

INVx3_ASAP7_75t_L g5087 ( 
.A(n_3976),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4326),
.Y(n_5088)
);

OAI21x1_ASAP7_75t_SL g5089 ( 
.A1(n_4108),
.A2(n_3517),
.B(n_3489),
.Y(n_5089)
);

INVx2_ASAP7_75t_L g5090 ( 
.A(n_4009),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_4172),
.B(n_3765),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4343),
.Y(n_5092)
);

BUFx10_ASAP7_75t_L g5093 ( 
.A(n_4112),
.Y(n_5093)
);

CKINVDCx6p67_ASAP7_75t_R g5094 ( 
.A(n_4185),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4343),
.Y(n_5095)
);

AOI22xp5_ASAP7_75t_L g5096 ( 
.A1(n_4249),
.A2(n_3714),
.B1(n_3715),
.B2(n_3773),
.Y(n_5096)
);

BUFx8_ASAP7_75t_SL g5097 ( 
.A(n_4365),
.Y(n_5097)
);

AO21x2_ASAP7_75t_L g5098 ( 
.A1(n_3984),
.A2(n_4374),
.B(n_4373),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4013),
.Y(n_5099)
);

AOI21x1_ASAP7_75t_L g5100 ( 
.A1(n_4371),
.A2(n_3854),
.B(n_3846),
.Y(n_5100)
);

AND2x4_ASAP7_75t_L g5101 ( 
.A(n_4159),
.B(n_3625),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4346),
.Y(n_5102)
);

OAI21xp5_ASAP7_75t_L g5103 ( 
.A1(n_4067),
.A2(n_3684),
.B(n_3637),
.Y(n_5103)
);

HB1xp67_ASAP7_75t_L g5104 ( 
.A(n_4194),
.Y(n_5104)
);

BUFx3_ASAP7_75t_L g5105 ( 
.A(n_4213),
.Y(n_5105)
);

AOI22xp33_ASAP7_75t_L g5106 ( 
.A1(n_4376),
.A2(n_3648),
.B1(n_3635),
.B2(n_3708),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_4121),
.B(n_3765),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4013),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4848),
.Y(n_5109)
);

OR2x2_ASAP7_75t_L g5110 ( 
.A(n_4700),
.B(n_4443),
.Y(n_5110)
);

BUFx2_ASAP7_75t_L g5111 ( 
.A(n_4716),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_4930),
.B(n_4288),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4848),
.Y(n_5113)
);

BUFx3_ASAP7_75t_L g5114 ( 
.A(n_4599),
.Y(n_5114)
);

AND2x2_ASAP7_75t_L g5115 ( 
.A(n_4930),
.B(n_4291),
.Y(n_5115)
);

NOR2xp33_ASAP7_75t_L g5116 ( 
.A(n_4599),
.B(n_4213),
.Y(n_5116)
);

AOI21x1_ASAP7_75t_L g5117 ( 
.A1(n_4515),
.A2(n_4013),
.B(n_4371),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4448),
.Y(n_5118)
);

OR2x6_ASAP7_75t_L g5119 ( 
.A(n_4725),
.B(n_4155),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4448),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4935),
.B(n_4291),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_4495),
.Y(n_5122)
);

BUFx6f_ASAP7_75t_SL g5123 ( 
.A(n_4590),
.Y(n_5123)
);

BUFx3_ASAP7_75t_L g5124 ( 
.A(n_4447),
.Y(n_5124)
);

INVx2_ASAP7_75t_L g5125 ( 
.A(n_4495),
.Y(n_5125)
);

INVx5_ASAP7_75t_SL g5126 ( 
.A(n_5094),
.Y(n_5126)
);

INVx2_ASAP7_75t_L g5127 ( 
.A(n_4495),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_4453),
.Y(n_5128)
);

INVx5_ASAP7_75t_SL g5129 ( 
.A(n_5094),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4495),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_4506),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4961),
.B(n_4291),
.Y(n_5132)
);

AO21x2_ASAP7_75t_L g5133 ( 
.A1(n_4725),
.A2(n_4284),
.B(n_4268),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_4506),
.Y(n_5134)
);

OAI21x1_ASAP7_75t_L g5135 ( 
.A1(n_4676),
.A2(n_4353),
.B(n_4393),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4453),
.Y(n_5136)
);

INVx2_ASAP7_75t_L g5137 ( 
.A(n_4506),
.Y(n_5137)
);

OA21x2_ASAP7_75t_L g5138 ( 
.A1(n_4838),
.A2(n_4393),
.B(n_4566),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_4506),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_4551),
.Y(n_5140)
);

HB1xp67_ASAP7_75t_L g5141 ( 
.A(n_4748),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4731),
.B(n_4348),
.Y(n_5142)
);

HB1xp67_ASAP7_75t_L g5143 ( 
.A(n_4766),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_4700),
.B(n_4760),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4462),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4462),
.Y(n_5146)
);

BUFx2_ASAP7_75t_L g5147 ( 
.A(n_4717),
.Y(n_5147)
);

BUFx6f_ASAP7_75t_L g5148 ( 
.A(n_4590),
.Y(n_5148)
);

OAI21x1_ASAP7_75t_L g5149 ( 
.A1(n_4676),
.A2(n_4393),
.B(n_4430),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4467),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_4551),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_4467),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4471),
.Y(n_5153)
);

BUFx6f_ASAP7_75t_L g5154 ( 
.A(n_4590),
.Y(n_5154)
);

HB1xp67_ASAP7_75t_L g5155 ( 
.A(n_4944),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4471),
.Y(n_5156)
);

OAI21x1_ASAP7_75t_L g5157 ( 
.A1(n_4690),
.A2(n_4430),
.B(n_4397),
.Y(n_5157)
);

AOI221xp5_ASAP7_75t_SL g5158 ( 
.A1(n_4598),
.A2(n_4096),
.B1(n_4111),
.B2(n_4101),
.C(n_4120),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4483),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4483),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4484),
.Y(n_5161)
);

INVx3_ASAP7_75t_L g5162 ( 
.A(n_4551),
.Y(n_5162)
);

O2A1O1Ixp5_ASAP7_75t_L g5163 ( 
.A1(n_4566),
.A2(n_4277),
.B(n_4096),
.C(n_4390),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4551),
.Y(n_5164)
);

BUFx6f_ASAP7_75t_L g5165 ( 
.A(n_4461),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_4935),
.B(n_4348),
.Y(n_5166)
);

BUFx6f_ASAP7_75t_L g5167 ( 
.A(n_4461),
.Y(n_5167)
);

OAI21x1_ASAP7_75t_L g5168 ( 
.A1(n_4690),
.A2(n_4430),
.B(n_4397),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4484),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4487),
.Y(n_5170)
);

AND2x4_ASAP7_75t_L g5171 ( 
.A(n_4922),
.B(n_4159),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4487),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_4939),
.B(n_4356),
.Y(n_5173)
);

OR2x2_ASAP7_75t_L g5174 ( 
.A(n_4760),
.B(n_4194),
.Y(n_5174)
);

BUFx6f_ASAP7_75t_L g5175 ( 
.A(n_4449),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4488),
.Y(n_5176)
);

AND2x2_ASAP7_75t_L g5177 ( 
.A(n_4939),
.B(n_4356),
.Y(n_5177)
);

INVx2_ASAP7_75t_L g5178 ( 
.A(n_4556),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4556),
.Y(n_5179)
);

CKINVDCx20_ASAP7_75t_R g5180 ( 
.A(n_4469),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_4949),
.B(n_4356),
.Y(n_5181)
);

AND2x4_ASAP7_75t_L g5182 ( 
.A(n_4922),
.B(n_4159),
.Y(n_5182)
);

INVx2_ASAP7_75t_L g5183 ( 
.A(n_4556),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4556),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4488),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_4563),
.Y(n_5186)
);

BUFx3_ASAP7_75t_L g5187 ( 
.A(n_4447),
.Y(n_5187)
);

INVx2_ASAP7_75t_SL g5188 ( 
.A(n_4673),
.Y(n_5188)
);

INVxp67_ASAP7_75t_SL g5189 ( 
.A(n_4989),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4489),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_4563),
.Y(n_5191)
);

NOR2x1_ASAP7_75t_R g5192 ( 
.A(n_4449),
.B(n_4372),
.Y(n_5192)
);

OA21x2_ASAP7_75t_L g5193 ( 
.A1(n_4896),
.A2(n_4073),
.B(n_4396),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4489),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_4492),
.Y(n_5195)
);

OR2x2_ASAP7_75t_L g5196 ( 
.A(n_4788),
.B(n_4194),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_4470),
.Y(n_5197)
);

AOI22xp33_ASAP7_75t_L g5198 ( 
.A1(n_4754),
.A2(n_4376),
.B1(n_4377),
.B2(n_4312),
.Y(n_5198)
);

INVx2_ASAP7_75t_L g5199 ( 
.A(n_4563),
.Y(n_5199)
);

INVx5_ASAP7_75t_L g5200 ( 
.A(n_4673),
.Y(n_5200)
);

HB1xp67_ASAP7_75t_L g5201 ( 
.A(n_4455),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_4563),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4492),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_4595),
.Y(n_5204)
);

AOI22xp33_ASAP7_75t_L g5205 ( 
.A1(n_4785),
.A2(n_4376),
.B1(n_4377),
.B2(n_4312),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4501),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4501),
.Y(n_5207)
);

NOR2x1p5_ASAP7_75t_L g5208 ( 
.A(n_4491),
.B(n_4213),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4505),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_4505),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4513),
.Y(n_5211)
);

OAI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4841),
.A2(n_4089),
.B(n_4101),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_4513),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4518),
.Y(n_5214)
);

HB1xp67_ASAP7_75t_L g5215 ( 
.A(n_4466),
.Y(n_5215)
);

AOI21x1_ASAP7_75t_L g5216 ( 
.A1(n_4515),
.A2(n_4308),
.B(n_4048),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_4595),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_4949),
.B(n_3958),
.Y(n_5218)
);

AOI22xp33_ASAP7_75t_L g5219 ( 
.A1(n_4677),
.A2(n_4377),
.B1(n_4312),
.B2(n_4349),
.Y(n_5219)
);

OR2x2_ASAP7_75t_L g5220 ( 
.A(n_4788),
.B(n_4121),
.Y(n_5220)
);

HB1xp67_ASAP7_75t_SL g5221 ( 
.A(n_4447),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_4595),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4518),
.Y(n_5223)
);

OAI21x1_ASAP7_75t_L g5224 ( 
.A1(n_4837),
.A2(n_4397),
.B(n_4396),
.Y(n_5224)
);

OR2x2_ASAP7_75t_L g5225 ( 
.A(n_5002),
.B(n_4154),
.Y(n_5225)
);

NOR2xp33_ASAP7_75t_R g5226 ( 
.A(n_4592),
.B(n_4372),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_4522),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_4595),
.Y(n_5228)
);

AO21x2_ASAP7_75t_L g5229 ( 
.A1(n_4837),
.A2(n_4284),
.B(n_4268),
.Y(n_5229)
);

INVx2_ASAP7_75t_SL g5230 ( 
.A(n_4673),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4522),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_4525),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4525),
.Y(n_5233)
);

BUFx2_ASAP7_75t_L g5234 ( 
.A(n_4993),
.Y(n_5234)
);

HB1xp67_ASAP7_75t_L g5235 ( 
.A(n_4500),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_4596),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_4596),
.Y(n_5237)
);

OAI22xp5_ASAP7_75t_L g5238 ( 
.A1(n_4810),
.A2(n_4189),
.B1(n_4171),
.B2(n_4111),
.Y(n_5238)
);

AND2x2_ASAP7_75t_L g5239 ( 
.A(n_4927),
.B(n_3958),
.Y(n_5239)
);

OAI21x1_ASAP7_75t_L g5240 ( 
.A1(n_4953),
.A2(n_4396),
.B(n_4073),
.Y(n_5240)
);

INVxp67_ASAP7_75t_SL g5241 ( 
.A(n_4989),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_4596),
.Y(n_5242)
);

CKINVDCx5p33_ASAP7_75t_R g5243 ( 
.A(n_4603),
.Y(n_5243)
);

OAI21x1_ASAP7_75t_L g5244 ( 
.A1(n_4953),
.A2(n_4073),
.B(n_4404),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_4596),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_4458),
.B(n_4239),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4526),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_4526),
.Y(n_5248)
);

HB1xp67_ASAP7_75t_L g5249 ( 
.A(n_4519),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4536),
.Y(n_5250)
);

INVx2_ASAP7_75t_SL g5251 ( 
.A(n_4673),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_4612),
.Y(n_5252)
);

INVx3_ASAP7_75t_L g5253 ( 
.A(n_4612),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4536),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_4967),
.B(n_4239),
.Y(n_5255)
);

OR2x2_ASAP7_75t_L g5256 ( 
.A(n_5002),
.B(n_4154),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_4498),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_4612),
.Y(n_5258)
);

BUFx10_ASAP7_75t_L g5259 ( 
.A(n_4541),
.Y(n_5259)
);

OAI21x1_ASAP7_75t_L g5260 ( 
.A1(n_4868),
.A2(n_4404),
.B(n_4416),
.Y(n_5260)
);

INVx2_ASAP7_75t_SL g5261 ( 
.A(n_4673),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_4612),
.Y(n_5262)
);

OAI21x1_ASAP7_75t_L g5263 ( 
.A1(n_4868),
.A2(n_4404),
.B(n_4416),
.Y(n_5263)
);

BUFx2_ASAP7_75t_L g5264 ( 
.A(n_4642),
.Y(n_5264)
);

BUFx3_ASAP7_75t_L g5265 ( 
.A(n_4447),
.Y(n_5265)
);

AO21x2_ASAP7_75t_L g5266 ( 
.A1(n_5098),
.A2(n_4319),
.B(n_4289),
.Y(n_5266)
);

OAI21x1_ASAP7_75t_L g5267 ( 
.A1(n_4840),
.A2(n_4424),
.B(n_4416),
.Y(n_5267)
);

AND2x2_ASAP7_75t_L g5268 ( 
.A(n_4927),
.B(n_3958),
.Y(n_5268)
);

BUFx5_ASAP7_75t_L g5269 ( 
.A(n_4601),
.Y(n_5269)
);

HB1xp67_ASAP7_75t_L g5270 ( 
.A(n_4521),
.Y(n_5270)
);

BUFx2_ASAP7_75t_L g5271 ( 
.A(n_4718),
.Y(n_5271)
);

OAI21x1_ASAP7_75t_L g5272 ( 
.A1(n_4840),
.A2(n_4424),
.B(n_4192),
.Y(n_5272)
);

HB1xp67_ASAP7_75t_L g5273 ( 
.A(n_4543),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_4537),
.Y(n_5274)
);

HB1xp67_ASAP7_75t_L g5275 ( 
.A(n_4574),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5107),
.B(n_4239),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_4621),
.Y(n_5277)
);

OAI22xp5_ASAP7_75t_L g5278 ( 
.A1(n_4841),
.A2(n_4189),
.B1(n_4398),
.B2(n_4298),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4537),
.Y(n_5279)
);

INVx3_ASAP7_75t_L g5280 ( 
.A(n_4621),
.Y(n_5280)
);

AOI22xp33_ASAP7_75t_L g5281 ( 
.A1(n_4830),
.A2(n_4377),
.B1(n_4349),
.B2(n_4342),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4548),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4548),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4549),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_4621),
.Y(n_5285)
);

AND2x4_ASAP7_75t_L g5286 ( 
.A(n_4922),
.B(n_4424),
.Y(n_5286)
);

INVx3_ASAP7_75t_L g5287 ( 
.A(n_4621),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_4549),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_4624),
.Y(n_5289)
);

BUFx6f_ASAP7_75t_L g5290 ( 
.A(n_4491),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_4972),
.B(n_4241),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4550),
.Y(n_5292)
);

OR2x2_ASAP7_75t_L g5293 ( 
.A(n_4790),
.B(n_4898),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_4624),
.Y(n_5294)
);

INVx2_ASAP7_75t_L g5295 ( 
.A(n_4624),
.Y(n_5295)
);

AOI21xp5_ASAP7_75t_L g5296 ( 
.A1(n_4493),
.A2(n_4228),
.B(n_4412),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_4550),
.Y(n_5297)
);

INVx3_ASAP7_75t_L g5298 ( 
.A(n_4624),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_4625),
.Y(n_5299)
);

INVx3_ASAP7_75t_L g5300 ( 
.A(n_5073),
.Y(n_5300)
);

INVx8_ASAP7_75t_L g5301 ( 
.A(n_4577),
.Y(n_5301)
);

OR2x2_ASAP7_75t_L g5302 ( 
.A(n_4790),
.B(n_4304),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_4568),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4568),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4573),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_4625),
.Y(n_5306)
);

AND2x2_ASAP7_75t_L g5307 ( 
.A(n_4972),
.B(n_4241),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_4573),
.Y(n_5308)
);

INVx2_ASAP7_75t_L g5309 ( 
.A(n_4629),
.Y(n_5309)
);

BUFx3_ASAP7_75t_L g5310 ( 
.A(n_4571),
.Y(n_5310)
);

BUFx4f_ASAP7_75t_SL g5311 ( 
.A(n_4485),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_4629),
.Y(n_5312)
);

AO21x2_ASAP7_75t_L g5313 ( 
.A1(n_5098),
.A2(n_4319),
.B(n_4289),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4633),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_4581),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_4633),
.Y(n_5316)
);

INVx1_ASAP7_75t_SL g5317 ( 
.A(n_4709),
.Y(n_5317)
);

XOR2xp5_ASAP7_75t_L g5318 ( 
.A(n_4992),
.B(n_4244),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_4476),
.B(n_4241),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4581),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4586),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_4586),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_4594),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_4594),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_4600),
.Y(n_5325)
);

AND2x2_ASAP7_75t_L g5326 ( 
.A(n_4476),
.B(n_4248),
.Y(n_5326)
);

HB1xp67_ASAP7_75t_L g5327 ( 
.A(n_4588),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_4600),
.Y(n_5328)
);

OR2x6_ASAP7_75t_L g5329 ( 
.A(n_4544),
.B(n_4431),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4604),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4604),
.Y(n_5331)
);

BUFx6f_ASAP7_75t_L g5332 ( 
.A(n_4491),
.Y(n_5332)
);

INVx2_ASAP7_75t_SL g5333 ( 
.A(n_4577),
.Y(n_5333)
);

INVx2_ASAP7_75t_L g5334 ( 
.A(n_4634),
.Y(n_5334)
);

OR2x6_ASAP7_75t_L g5335 ( 
.A(n_4544),
.B(n_4431),
.Y(n_5335)
);

INVx2_ASAP7_75t_L g5336 ( 
.A(n_4634),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_4703),
.A2(n_4358),
.B(n_4064),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_4605),
.Y(n_5338)
);

BUFx3_ASAP7_75t_L g5339 ( 
.A(n_4571),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_4635),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_4605),
.Y(n_5341)
);

CKINVDCx5p33_ASAP7_75t_R g5342 ( 
.A(n_4704),
.Y(n_5342)
);

INVx2_ASAP7_75t_L g5343 ( 
.A(n_4635),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_4606),
.Y(n_5344)
);

CKINVDCx20_ASAP7_75t_R g5345 ( 
.A(n_4593),
.Y(n_5345)
);

INVx2_ASAP7_75t_L g5346 ( 
.A(n_4901),
.Y(n_5346)
);

OAI22xp5_ASAP7_75t_L g5347 ( 
.A1(n_4978),
.A2(n_4398),
.B1(n_4298),
.B2(n_4120),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_4606),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_4901),
.Y(n_5349)
);

AO21x1_ASAP7_75t_L g5350 ( 
.A1(n_4983),
.A2(n_4164),
.B(n_4064),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4609),
.Y(n_5351)
);

INVx3_ASAP7_75t_L g5352 ( 
.A(n_5073),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_4901),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4609),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4610),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_4901),
.Y(n_5356)
);

BUFx6f_ASAP7_75t_L g5357 ( 
.A(n_4514),
.Y(n_5357)
);

INVx3_ASAP7_75t_L g5358 ( 
.A(n_5073),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_4610),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_4611),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4611),
.Y(n_5361)
);

AND2x4_ASAP7_75t_L g5362 ( 
.A(n_4922),
.B(n_4307),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_4613),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4613),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_4454),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_4616),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_4454),
.Y(n_5367)
);

INVx2_ASAP7_75t_L g5368 ( 
.A(n_4454),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_4616),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_4460),
.Y(n_5370)
);

OA21x2_ASAP7_75t_L g5371 ( 
.A1(n_4896),
.A2(n_4374),
.B(n_4373),
.Y(n_5371)
);

AOI22xp5_ASAP7_75t_L g5372 ( 
.A1(n_4538),
.A2(n_4249),
.B1(n_4220),
.B2(n_4161),
.Y(n_5372)
);

INVx4_ASAP7_75t_L g5373 ( 
.A(n_4577),
.Y(n_5373)
);

CKINVDCx5p33_ASAP7_75t_R g5374 ( 
.A(n_4554),
.Y(n_5374)
);

INVx6_ASAP7_75t_L g5375 ( 
.A(n_4756),
.Y(n_5375)
);

BUFx3_ASAP7_75t_L g5376 ( 
.A(n_4450),
.Y(n_5376)
);

AND2x2_ASAP7_75t_L g5377 ( 
.A(n_4539),
.B(n_4248),
.Y(n_5377)
);

HB1xp67_ASAP7_75t_L g5378 ( 
.A(n_4615),
.Y(n_5378)
);

INVx3_ASAP7_75t_L g5379 ( 
.A(n_5073),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_4622),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_4622),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_4460),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_4460),
.Y(n_5383)
);

BUFx2_ASAP7_75t_L g5384 ( 
.A(n_4718),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4637),
.Y(n_5385)
);

AO21x2_ASAP7_75t_L g5386 ( 
.A1(n_5098),
.A2(n_4325),
.B(n_4322),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_4637),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_5030),
.B(n_5091),
.Y(n_5388)
);

HB1xp67_ASAP7_75t_L g5389 ( 
.A(n_4620),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4561),
.B(n_4643),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_4463),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_4640),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_4560),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4463),
.Y(n_5394)
);

AND2x2_ASAP7_75t_L g5395 ( 
.A(n_4539),
.B(n_4248),
.Y(n_5395)
);

OR2x2_ASAP7_75t_L g5396 ( 
.A(n_4898),
.B(n_4304),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_4463),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_4468),
.Y(n_5398)
);

HB1xp67_ASAP7_75t_L g5399 ( 
.A(n_4664),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_4660),
.B(n_4263),
.Y(n_5400)
);

AO21x1_ASAP7_75t_SL g5401 ( 
.A1(n_5001),
.A2(n_4422),
.B(n_4307),
.Y(n_5401)
);

INVx3_ASAP7_75t_L g5402 ( 
.A(n_4918),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_4640),
.Y(n_5403)
);

INVx2_ASAP7_75t_L g5404 ( 
.A(n_4468),
.Y(n_5404)
);

OR2x2_ASAP7_75t_L g5405 ( 
.A(n_4908),
.B(n_4304),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4646),
.Y(n_5406)
);

INVx2_ASAP7_75t_SL g5407 ( 
.A(n_4577),
.Y(n_5407)
);

OR2x2_ASAP7_75t_L g5408 ( 
.A(n_4908),
.B(n_4266),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_4646),
.Y(n_5409)
);

HB1xp67_ASAP7_75t_L g5410 ( 
.A(n_4687),
.Y(n_5410)
);

INVx2_ASAP7_75t_SL g5411 ( 
.A(n_4577),
.Y(n_5411)
);

AND2x2_ASAP7_75t_L g5412 ( 
.A(n_4660),
.B(n_4263),
.Y(n_5412)
);

OR2x2_ASAP7_75t_L g5413 ( 
.A(n_4650),
.B(n_4266),
.Y(n_5413)
);

OAI21xp5_ASAP7_75t_L g5414 ( 
.A1(n_4969),
.A2(n_4114),
.B(n_4215),
.Y(n_5414)
);

INVx3_ASAP7_75t_L g5415 ( 
.A(n_4918),
.Y(n_5415)
);

AND2x2_ASAP7_75t_L g5416 ( 
.A(n_4713),
.B(n_4263),
.Y(n_5416)
);

HB1xp67_ASAP7_75t_L g5417 ( 
.A(n_4702),
.Y(n_5417)
);

INVx2_ASAP7_75t_L g5418 ( 
.A(n_4468),
.Y(n_5418)
);

OR2x2_ASAP7_75t_L g5419 ( 
.A(n_4650),
.B(n_3986),
.Y(n_5419)
);

BUFx2_ASAP7_75t_L g5420 ( 
.A(n_4718),
.Y(n_5420)
);

HB1xp67_ASAP7_75t_SL g5421 ( 
.A(n_4579),
.Y(n_5421)
);

AOI21x1_ASAP7_75t_L g5422 ( 
.A1(n_4540),
.A2(n_4308),
.B(n_4048),
.Y(n_5422)
);

INVx2_ASAP7_75t_L g5423 ( 
.A(n_4914),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_4651),
.Y(n_5424)
);

INVx4_ASAP7_75t_SL g5425 ( 
.A(n_4450),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_4651),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_4914),
.Y(n_5427)
);

BUFx2_ASAP7_75t_SL g5428 ( 
.A(n_4910),
.Y(n_5428)
);

OAI21x1_ASAP7_75t_L g5429 ( 
.A1(n_4540),
.A2(n_4192),
.B(n_4373),
.Y(n_5429)
);

AND2x4_ASAP7_75t_L g5430 ( 
.A(n_4922),
.B(n_3942),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_4914),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_4656),
.Y(n_5432)
);

INVx2_ASAP7_75t_L g5433 ( 
.A(n_4914),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_4656),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_4661),
.Y(n_5435)
);

INVx3_ASAP7_75t_L g5436 ( 
.A(n_4918),
.Y(n_5436)
);

INVx2_ASAP7_75t_SL g5437 ( 
.A(n_4541),
.Y(n_5437)
);

NOR2xp33_ASAP7_75t_L g5438 ( 
.A(n_4979),
.B(n_4083),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_4661),
.Y(n_5439)
);

BUFx2_ASAP7_75t_L g5440 ( 
.A(n_4718),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_4665),
.Y(n_5441)
);

INVx2_ASAP7_75t_L g5442 ( 
.A(n_4472),
.Y(n_5442)
);

OAI21x1_ASAP7_75t_L g5443 ( 
.A1(n_5004),
.A2(n_4192),
.B(n_4374),
.Y(n_5443)
);

BUFx2_ASAP7_75t_L g5444 ( 
.A(n_4756),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_4472),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_4472),
.Y(n_5446)
);

INVx2_ASAP7_75t_L g5447 ( 
.A(n_4473),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_4665),
.Y(n_5448)
);

INVx2_ASAP7_75t_SL g5449 ( 
.A(n_4541),
.Y(n_5449)
);

INVx2_ASAP7_75t_L g5450 ( 
.A(n_4473),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_4473),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_4649),
.B(n_3986),
.Y(n_5452)
);

OAI21x1_ASAP7_75t_L g5453 ( 
.A1(n_5004),
.A2(n_4294),
.B(n_4290),
.Y(n_5453)
);

HB1xp67_ASAP7_75t_L g5454 ( 
.A(n_4720),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_4477),
.Y(n_5455)
);

INVx2_ASAP7_75t_L g5456 ( 
.A(n_4477),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_4477),
.Y(n_5457)
);

AND2x2_ASAP7_75t_L g5458 ( 
.A(n_4713),
.B(n_4076),
.Y(n_5458)
);

BUFx3_ASAP7_75t_L g5459 ( 
.A(n_4450),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_4666),
.Y(n_5460)
);

NAND2x1p5_ASAP7_75t_L g5461 ( 
.A(n_4922),
.B(n_4254),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4666),
.Y(n_5462)
);

INVxp67_ASAP7_75t_L g5463 ( 
.A(n_4734),
.Y(n_5463)
);

AND2x4_ASAP7_75t_L g5464 ( 
.A(n_4995),
.B(n_3942),
.Y(n_5464)
);

HB1xp67_ASAP7_75t_L g5465 ( 
.A(n_4724),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_4679),
.Y(n_5466)
);

AOI21xp5_ASAP7_75t_L g5467 ( 
.A1(n_4943),
.A2(n_4808),
.B(n_5103),
.Y(n_5467)
);

INVx3_ASAP7_75t_L g5468 ( 
.A(n_4918),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_4478),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_4478),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_4679),
.Y(n_5471)
);

INVx2_ASAP7_75t_L g5472 ( 
.A(n_4524),
.Y(n_5472)
);

AND2x2_ASAP7_75t_L g5473 ( 
.A(n_4715),
.B(n_4076),
.Y(n_5473)
);

BUFx4f_ASAP7_75t_SL g5474 ( 
.A(n_4869),
.Y(n_5474)
);

AOI221xp5_ASAP7_75t_L g5475 ( 
.A1(n_5031),
.A2(n_4277),
.B1(n_4271),
.B2(n_4325),
.C(n_4322),
.Y(n_5475)
);

OR2x6_ASAP7_75t_L g5476 ( 
.A(n_4544),
.B(n_4215),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_4682),
.Y(n_5477)
);

INVx3_ASAP7_75t_L g5478 ( 
.A(n_5027),
.Y(n_5478)
);

AND2x2_ASAP7_75t_L g5479 ( 
.A(n_4715),
.B(n_4076),
.Y(n_5479)
);

AND2x4_ASAP7_75t_L g5480 ( 
.A(n_4995),
.B(n_3942),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_4682),
.Y(n_5481)
);

OAI21x1_ASAP7_75t_L g5482 ( 
.A1(n_5009),
.A2(n_4294),
.B(n_4290),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_4686),
.Y(n_5483)
);

OAI21x1_ASAP7_75t_L g5484 ( 
.A1(n_5009),
.A2(n_5012),
.B(n_5100),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_4524),
.Y(n_5485)
);

HB1xp67_ASAP7_75t_L g5486 ( 
.A(n_4733),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_4686),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_4695),
.Y(n_5488)
);

INVx2_ASAP7_75t_L g5489 ( 
.A(n_4524),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_4695),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_4527),
.Y(n_5491)
);

INVxp67_ASAP7_75t_L g5492 ( 
.A(n_4963),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_4696),
.Y(n_5493)
);

INVx3_ASAP7_75t_L g5494 ( 
.A(n_5027),
.Y(n_5494)
);

HB1xp67_ASAP7_75t_L g5495 ( 
.A(n_4867),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_4696),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_4697),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_4697),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_4527),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_4701),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_4527),
.Y(n_5501)
);

INVx2_ASAP7_75t_L g5502 ( 
.A(n_4847),
.Y(n_5502)
);

OAI21x1_ASAP7_75t_L g5503 ( 
.A1(n_5012),
.A2(n_4294),
.B(n_4290),
.Y(n_5503)
);

HB1xp67_ASAP7_75t_L g5504 ( 
.A(n_4880),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_4847),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_4701),
.Y(n_5506)
);

OR2x2_ASAP7_75t_L g5507 ( 
.A(n_4649),
.B(n_3986),
.Y(n_5507)
);

INVx2_ASAP7_75t_SL g5508 ( 
.A(n_4541),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_4722),
.Y(n_5509)
);

BUFx2_ASAP7_75t_L g5510 ( 
.A(n_4756),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_4502),
.Y(n_5511)
);

BUFx2_ASAP7_75t_L g5512 ( 
.A(n_4756),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_4722),
.Y(n_5513)
);

OAI21xp5_ASAP7_75t_L g5514 ( 
.A1(n_5038),
.A2(n_4114),
.B(n_4313),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_4502),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_4729),
.Y(n_5516)
);

NOR2xp33_ASAP7_75t_L g5517 ( 
.A(n_5018),
.B(n_4083),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_4503),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_4729),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_4730),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_4730),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_4503),
.Y(n_5522)
);

AND2x2_ASAP7_75t_L g5523 ( 
.A(n_4745),
.B(n_4079),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_4647),
.B(n_4313),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_4740),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_4740),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_L g5527 ( 
.A(n_4570),
.B(n_4240),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_4890),
.B(n_4237),
.Y(n_5528)
);

INVx4_ASAP7_75t_L g5529 ( 
.A(n_4514),
.Y(n_5529)
);

INVx3_ASAP7_75t_L g5530 ( 
.A(n_5027),
.Y(n_5530)
);

INVx2_ASAP7_75t_L g5531 ( 
.A(n_4509),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_4742),
.Y(n_5532)
);

BUFx6f_ASAP7_75t_L g5533 ( 
.A(n_4514),
.Y(n_5533)
);

OR2x2_ASAP7_75t_L g5534 ( 
.A(n_5086),
.B(n_4015),
.Y(n_5534)
);

INVx2_ASAP7_75t_L g5535 ( 
.A(n_4509),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_4512),
.Y(n_5536)
);

BUFx3_ASAP7_75t_L g5537 ( 
.A(n_4450),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_4512),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_4745),
.B(n_4787),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_4742),
.Y(n_5540)
);

INVx2_ASAP7_75t_SL g5541 ( 
.A(n_4523),
.Y(n_5541)
);

BUFx2_ASAP7_75t_L g5542 ( 
.A(n_4756),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_4787),
.B(n_4798),
.Y(n_5543)
);

OR2x6_ASAP7_75t_L g5544 ( 
.A(n_4504),
.B(n_4238),
.Y(n_5544)
);

OA21x2_ASAP7_75t_L g5545 ( 
.A1(n_5031),
.A2(n_4098),
.B(n_4094),
.Y(n_5545)
);

HB1xp67_ASAP7_75t_L g5546 ( 
.A(n_4886),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_4750),
.Y(n_5547)
);

INVx2_ASAP7_75t_L g5548 ( 
.A(n_4528),
.Y(n_5548)
);

OAI21x1_ASAP7_75t_L g5549 ( 
.A1(n_5100),
.A2(n_3985),
.B(n_3961),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_4528),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_4798),
.B(n_4079),
.Y(n_5551)
);

BUFx3_ASAP7_75t_L g5552 ( 
.A(n_4508),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_4564),
.Y(n_5553)
);

BUFx2_ASAP7_75t_L g5554 ( 
.A(n_5097),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_4750),
.Y(n_5555)
);

NAND2x1_ASAP7_75t_L g5556 ( 
.A(n_4809),
.B(n_4270),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4752),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_4508),
.Y(n_5558)
);

AND2x2_ASAP7_75t_L g5559 ( 
.A(n_4889),
.B(n_4079),
.Y(n_5559)
);

INVx2_ASAP7_75t_L g5560 ( 
.A(n_4564),
.Y(n_5560)
);

OAI22xp5_ASAP7_75t_L g5561 ( 
.A1(n_4978),
.A2(n_4161),
.B1(n_4399),
.B2(n_4414),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_4752),
.Y(n_5562)
);

INVx4_ASAP7_75t_L g5563 ( 
.A(n_4523),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_4576),
.Y(n_5564)
);

BUFx2_ASAP7_75t_L g5565 ( 
.A(n_5010),
.Y(n_5565)
);

OAI21x1_ASAP7_75t_L g5566 ( 
.A1(n_4749),
.A2(n_3985),
.B(n_3961),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_4753),
.Y(n_5567)
);

INVx4_ASAP7_75t_L g5568 ( 
.A(n_4523),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_4753),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_4758),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_4576),
.Y(n_5571)
);

BUFx12f_ASAP7_75t_L g5572 ( 
.A(n_5075),
.Y(n_5572)
);

INVx3_ASAP7_75t_L g5573 ( 
.A(n_5027),
.Y(n_5573)
);

INVx2_ASAP7_75t_SL g5574 ( 
.A(n_4529),
.Y(n_5574)
);

HB1xp67_ASAP7_75t_L g5575 ( 
.A(n_4904),
.Y(n_5575)
);

AND2x2_ASAP7_75t_L g5576 ( 
.A(n_4889),
.B(n_4086),
.Y(n_5576)
);

NOR2xp33_ASAP7_75t_L g5577 ( 
.A(n_4636),
.B(n_4233),
.Y(n_5577)
);

INVx2_ASAP7_75t_L g5578 ( 
.A(n_4602),
.Y(n_5578)
);

INVx2_ASAP7_75t_SL g5579 ( 
.A(n_4529),
.Y(n_5579)
);

INVx1_ASAP7_75t_SL g5580 ( 
.A(n_4782),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_4758),
.Y(n_5581)
);

INVx3_ASAP7_75t_L g5582 ( 
.A(n_4601),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_4762),
.Y(n_5583)
);

BUFx2_ASAP7_75t_L g5584 ( 
.A(n_5010),
.Y(n_5584)
);

INVx2_ASAP7_75t_L g5585 ( 
.A(n_4602),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_4893),
.B(n_4237),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_4762),
.Y(n_5587)
);

BUFx3_ASAP7_75t_L g5588 ( 
.A(n_4508),
.Y(n_5588)
);

AND2x2_ASAP7_75t_L g5589 ( 
.A(n_4892),
.B(n_4086),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_4764),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_4764),
.Y(n_5591)
);

BUFx2_ASAP7_75t_L g5592 ( 
.A(n_4529),
.Y(n_5592)
);

AOI21x1_ASAP7_75t_L g5593 ( 
.A1(n_4749),
.A2(n_4779),
.B(n_5060),
.Y(n_5593)
);

AND2x4_ASAP7_75t_L g5594 ( 
.A(n_4995),
.B(n_3942),
.Y(n_5594)
);

NOR2xp33_ASAP7_75t_SL g5595 ( 
.A(n_4597),
.B(n_4173),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_4767),
.Y(n_5596)
);

AND2x4_ASAP7_75t_L g5597 ( 
.A(n_4995),
.B(n_3942),
.Y(n_5597)
);

AOI22xp33_ASAP7_75t_L g5598 ( 
.A1(n_5060),
.A2(n_4377),
.B1(n_4349),
.B2(n_4342),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_4619),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_4892),
.B(n_4086),
.Y(n_5600)
);

INVx2_ASAP7_75t_L g5601 ( 
.A(n_4619),
.Y(n_5601)
);

BUFx2_ASAP7_75t_L g5602 ( 
.A(n_4531),
.Y(n_5602)
);

BUFx2_ASAP7_75t_L g5603 ( 
.A(n_4531),
.Y(n_5603)
);

INVx2_ASAP7_75t_L g5604 ( 
.A(n_4619),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_4767),
.Y(n_5605)
);

INVx2_ASAP7_75t_L g5606 ( 
.A(n_4619),
.Y(n_5606)
);

BUFx2_ASAP7_75t_SL g5607 ( 
.A(n_5029),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_4771),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_4542),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_4542),
.Y(n_5610)
);

AND2x2_ASAP7_75t_L g5611 ( 
.A(n_4932),
.B(n_4031),
.Y(n_5611)
);

NOR2xp33_ASAP7_75t_SL g5612 ( 
.A(n_4508),
.B(n_4173),
.Y(n_5612)
);

BUFx12f_ASAP7_75t_L g5613 ( 
.A(n_4799),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_4542),
.Y(n_5614)
);

CKINVDCx6p67_ASAP7_75t_R g5615 ( 
.A(n_5049),
.Y(n_5615)
);

BUFx3_ASAP7_75t_L g5616 ( 
.A(n_4465),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_4771),
.Y(n_5617)
);

BUFx10_ASAP7_75t_L g5618 ( 
.A(n_4465),
.Y(n_5618)
);

AND2x4_ASAP7_75t_L g5619 ( 
.A(n_4995),
.B(n_3945),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_4907),
.B(n_4210),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_4772),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_4772),
.Y(n_5622)
);

HB1xp67_ASAP7_75t_L g5623 ( 
.A(n_4769),
.Y(n_5623)
);

NAND2xp5_ASAP7_75t_L g5624 ( 
.A(n_4732),
.B(n_4210),
.Y(n_5624)
);

INVx2_ASAP7_75t_SL g5625 ( 
.A(n_5052),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_4773),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_4773),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_4786),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_4786),
.Y(n_5629)
);

INVx2_ASAP7_75t_L g5630 ( 
.A(n_4546),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_4791),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_4546),
.Y(n_5632)
);

OR2x6_ASAP7_75t_L g5633 ( 
.A(n_4504),
.B(n_4507),
.Y(n_5633)
);

OAI21x1_ASAP7_75t_L g5634 ( 
.A1(n_4779),
.A2(n_3985),
.B(n_3961),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_4791),
.Y(n_5635)
);

BUFx8_ASAP7_75t_SL g5636 ( 
.A(n_4517),
.Y(n_5636)
);

CKINVDCx5p33_ASAP7_75t_R g5637 ( 
.A(n_4820),
.Y(n_5637)
);

AND2x2_ASAP7_75t_L g5638 ( 
.A(n_4932),
.B(n_4031),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_4546),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_4793),
.Y(n_5640)
);

INVx2_ASAP7_75t_L g5641 ( 
.A(n_4547),
.Y(n_5641)
);

BUFx12f_ASAP7_75t_L g5642 ( 
.A(n_5021),
.Y(n_5642)
);

INVx2_ASAP7_75t_L g5643 ( 
.A(n_4547),
.Y(n_5643)
);

INVx2_ASAP7_75t_L g5644 ( 
.A(n_4547),
.Y(n_5644)
);

OAI21xp33_ASAP7_75t_SL g5645 ( 
.A1(n_5026),
.A2(n_4085),
.B(n_3977),
.Y(n_5645)
);

INVx3_ASAP7_75t_L g5646 ( 
.A(n_4601),
.Y(n_5646)
);

AOI222xp33_ASAP7_75t_L g5647 ( 
.A1(n_4674),
.A2(n_4271),
.B1(n_4375),
.B2(n_4383),
.C1(n_4381),
.C2(n_4220),
.Y(n_5647)
);

INVx1_ASAP7_75t_SL g5648 ( 
.A(n_4705),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_4819),
.B(n_4222),
.Y(n_5649)
);

AND2x4_ASAP7_75t_L g5650 ( 
.A(n_4995),
.B(n_3945),
.Y(n_5650)
);

BUFx2_ASAP7_75t_L g5651 ( 
.A(n_4531),
.Y(n_5651)
);

CKINVDCx14_ASAP7_75t_R g5652 ( 
.A(n_5045),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_4793),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_4552),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_4794),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5026),
.B(n_4031),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_4552),
.Y(n_5657)
);

INVx2_ASAP7_75t_L g5658 ( 
.A(n_4552),
.Y(n_5658)
);

HB1xp67_ASAP7_75t_L g5659 ( 
.A(n_4774),
.Y(n_5659)
);

INVx2_ASAP7_75t_SL g5660 ( 
.A(n_5052),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_4794),
.Y(n_5661)
);

AOI22xp5_ASAP7_75t_L g5662 ( 
.A1(n_4706),
.A2(n_4333),
.B1(n_4244),
.B2(n_4368),
.Y(n_5662)
);

BUFx2_ASAP7_75t_L g5663 ( 
.A(n_4531),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_4795),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_4795),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_4555),
.Y(n_5666)
);

AND2x2_ASAP7_75t_L g5667 ( 
.A(n_5068),
.B(n_4048),
.Y(n_5667)
);

AOI22xp5_ASAP7_75t_L g5668 ( 
.A1(n_4721),
.A2(n_4333),
.B1(n_4368),
.B2(n_4277),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_4555),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_4555),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_4559),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_4801),
.Y(n_5672)
);

AND2x2_ASAP7_75t_L g5673 ( 
.A(n_5068),
.B(n_3974),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_4801),
.Y(n_5674)
);

INVx2_ASAP7_75t_SL g5675 ( 
.A(n_5052),
.Y(n_5675)
);

AND2x2_ASAP7_75t_L g5676 ( 
.A(n_4821),
.B(n_3974),
.Y(n_5676)
);

INVx3_ASAP7_75t_L g5677 ( 
.A(n_4601),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_4803),
.Y(n_5678)
);

AND2x4_ASAP7_75t_L g5679 ( 
.A(n_5074),
.B(n_3945),
.Y(n_5679)
);

INVx2_ASAP7_75t_L g5680 ( 
.A(n_4559),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_4803),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_4559),
.Y(n_5682)
);

OAI21xp5_ASAP7_75t_L g5683 ( 
.A1(n_4817),
.A2(n_4134),
.B(n_4342),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_4805),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_4805),
.Y(n_5685)
);

AO21x2_ASAP7_75t_L g5686 ( 
.A1(n_4723),
.A2(n_3984),
.B(n_4128),
.Y(n_5686)
);

AND2x2_ASAP7_75t_L g5687 ( 
.A(n_4821),
.B(n_4075),
.Y(n_5687)
);

INVx2_ASAP7_75t_L g5688 ( 
.A(n_4569),
.Y(n_5688)
);

AOI22xp33_ASAP7_75t_SL g5689 ( 
.A1(n_4747),
.A2(n_4368),
.B1(n_3984),
.B2(n_4139),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_4569),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_4569),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_4815),
.Y(n_5692)
);

INVx2_ASAP7_75t_SL g5693 ( 
.A(n_5052),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_4815),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_4823),
.Y(n_5695)
);

OR2x6_ASAP7_75t_L g5696 ( 
.A(n_4504),
.B(n_4238),
.Y(n_5696)
);

AND2x2_ASAP7_75t_L g5697 ( 
.A(n_4829),
.B(n_4075),
.Y(n_5697)
);

INVx1_ASAP7_75t_SL g5698 ( 
.A(n_4744),
.Y(n_5698)
);

AO21x1_ASAP7_75t_L g5699 ( 
.A1(n_4958),
.A2(n_4331),
.B(n_4287),
.Y(n_5699)
);

AOI21x1_ASAP7_75t_L g5700 ( 
.A1(n_4452),
.A2(n_4338),
.B(n_3994),
.Y(n_5700)
);

AO21x2_ASAP7_75t_L g5701 ( 
.A1(n_4723),
.A2(n_3984),
.B(n_4128),
.Y(n_5701)
);

AO21x2_ASAP7_75t_L g5702 ( 
.A1(n_4723),
.A2(n_4128),
.B(n_4278),
.Y(n_5702)
);

AND2x2_ASAP7_75t_L g5703 ( 
.A(n_4829),
.B(n_4133),
.Y(n_5703)
);

NAND2x1_ASAP7_75t_L g5704 ( 
.A(n_4809),
.B(n_4270),
.Y(n_5704)
);

OAI21x1_ASAP7_75t_L g5705 ( 
.A1(n_4950),
.A2(n_3985),
.B(n_3961),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_4580),
.Y(n_5706)
);

INVx3_ASAP7_75t_L g5707 ( 
.A(n_4607),
.Y(n_5707)
);

BUFx2_ASAP7_75t_L g5708 ( 
.A(n_4688),
.Y(n_5708)
);

OAI21xp5_ASAP7_75t_L g5709 ( 
.A1(n_4817),
.A2(n_4278),
.B(n_4331),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_4823),
.Y(n_5710)
);

INVx2_ASAP7_75t_L g5711 ( 
.A(n_4580),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_4824),
.Y(n_5712)
);

INVx2_ASAP7_75t_L g5713 ( 
.A(n_4580),
.Y(n_5713)
);

INVx2_ASAP7_75t_L g5714 ( 
.A(n_4582),
.Y(n_5714)
);

OAI21x1_ASAP7_75t_L g5715 ( 
.A1(n_4950),
.A2(n_4092),
.B(n_3997),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_4582),
.Y(n_5716)
);

AOI22xp33_ASAP7_75t_L g5717 ( 
.A1(n_4751),
.A2(n_4389),
.B1(n_4271),
.B2(n_4368),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_4824),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_4825),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_4825),
.Y(n_5720)
);

BUFx6f_ASAP7_75t_L g5721 ( 
.A(n_4465),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_4582),
.Y(n_5722)
);

HB1xp67_ASAP7_75t_L g5723 ( 
.A(n_4777),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_4828),
.Y(n_5724)
);

INVx8_ASAP7_75t_L g5725 ( 
.A(n_4755),
.Y(n_5725)
);

OAI21x1_ASAP7_75t_L g5726 ( 
.A1(n_4950),
.A2(n_4092),
.B(n_3997),
.Y(n_5726)
);

OAI21x1_ASAP7_75t_L g5727 ( 
.A1(n_4962),
.A2(n_4092),
.B(n_3997),
.Y(n_5727)
);

AOI21x1_ASAP7_75t_L g5728 ( 
.A1(n_4452),
.A2(n_4338),
.B(n_3994),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_4828),
.Y(n_5729)
);

AND2x4_ASAP7_75t_L g5730 ( 
.A(n_5074),
.B(n_3945),
.Y(n_5730)
);

AND2x2_ASAP7_75t_L g5731 ( 
.A(n_4834),
.B(n_4133),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_4832),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_4832),
.Y(n_5733)
);

OAI21x1_ASAP7_75t_L g5734 ( 
.A1(n_4962),
.A2(n_4092),
.B(n_3997),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_4587),
.Y(n_5735)
);

HB1xp67_ASAP7_75t_L g5736 ( 
.A(n_4811),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5119),
.Y(n_5737)
);

AO21x2_ASAP7_75t_L g5738 ( 
.A1(n_5189),
.A2(n_4737),
.B(n_4728),
.Y(n_5738)
);

INVx2_ASAP7_75t_L g5739 ( 
.A(n_5119),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5190),
.Y(n_5740)
);

NAND2xp5_ASAP7_75t_L g5741 ( 
.A(n_5158),
.B(n_4915),
.Y(n_5741)
);

INVx4_ASAP7_75t_L g5742 ( 
.A(n_5165),
.Y(n_5742)
);

OAI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5216),
.A2(n_5005),
.B(n_4920),
.Y(n_5743)
);

HB1xp67_ASAP7_75t_L g5744 ( 
.A(n_5155),
.Y(n_5744)
);

INVx2_ASAP7_75t_L g5745 ( 
.A(n_5119),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5159),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5159),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5160),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5160),
.Y(n_5749)
);

OR2x2_ASAP7_75t_L g5750 ( 
.A(n_5225),
.B(n_4684),
.Y(n_5750)
);

OR2x2_ASAP7_75t_L g5751 ( 
.A(n_5225),
.B(n_4850),
.Y(n_5751)
);

INVxp67_ASAP7_75t_L g5752 ( 
.A(n_5421),
.Y(n_5752)
);

INVx1_ASAP7_75t_L g5753 ( 
.A(n_5161),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5161),
.Y(n_5754)
);

BUFx2_ASAP7_75t_L g5755 ( 
.A(n_5572),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5119),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5170),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_5170),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5325),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5325),
.Y(n_5760)
);

AO21x2_ASAP7_75t_L g5761 ( 
.A1(n_5241),
.A2(n_4737),
.B(n_4728),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5119),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5150),
.Y(n_5763)
);

BUFx2_ASAP7_75t_L g5764 ( 
.A(n_5572),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5150),
.Y(n_5765)
);

BUFx3_ASAP7_75t_L g5766 ( 
.A(n_5180),
.Y(n_5766)
);

OR2x2_ASAP7_75t_L g5767 ( 
.A(n_5256),
.B(n_4924),
.Y(n_5767)
);

OR2x2_ASAP7_75t_L g5768 ( 
.A(n_5256),
.B(n_4940),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5539),
.B(n_4714),
.Y(n_5769)
);

AND2x2_ASAP7_75t_L g5770 ( 
.A(n_5539),
.B(n_4714),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5207),
.Y(n_5771)
);

INVx3_ASAP7_75t_L g5772 ( 
.A(n_5216),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5599),
.Y(n_5773)
);

AND2x2_ASAP7_75t_L g5774 ( 
.A(n_5543),
.B(n_4714),
.Y(n_5774)
);

OR2x2_ASAP7_75t_L g5775 ( 
.A(n_5293),
.B(n_4964),
.Y(n_5775)
);

OR2x2_ASAP7_75t_L g5776 ( 
.A(n_5293),
.B(n_4456),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5599),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5601),
.Y(n_5778)
);

AND2x2_ASAP7_75t_L g5779 ( 
.A(n_5543),
.B(n_4802),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5601),
.Y(n_5780)
);

HB1xp67_ASAP7_75t_L g5781 ( 
.A(n_5141),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5152),
.Y(n_5782)
);

INVx3_ASAP7_75t_L g5783 ( 
.A(n_5422),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5152),
.Y(n_5784)
);

BUFx6f_ASAP7_75t_L g5785 ( 
.A(n_5114),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5153),
.Y(n_5786)
);

OR2x2_ASAP7_75t_L g5787 ( 
.A(n_5388),
.B(n_4456),
.Y(n_5787)
);

NAND2xp5_ASAP7_75t_L g5788 ( 
.A(n_5212),
.B(n_4915),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5604),
.Y(n_5789)
);

AO21x2_ASAP7_75t_L g5790 ( 
.A1(n_5350),
.A2(n_4737),
.B(n_4728),
.Y(n_5790)
);

OA21x2_ASAP7_75t_L g5791 ( 
.A1(n_5350),
.A2(n_4761),
.B(n_4746),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5604),
.Y(n_5792)
);

AND2x2_ASAP7_75t_L g5793 ( 
.A(n_5319),
.B(n_5326),
.Y(n_5793)
);

HB1xp67_ASAP7_75t_L g5794 ( 
.A(n_5143),
.Y(n_5794)
);

INVx3_ASAP7_75t_L g5795 ( 
.A(n_5422),
.Y(n_5795)
);

AND2x4_ASAP7_75t_L g5796 ( 
.A(n_5444),
.B(n_4911),
.Y(n_5796)
);

OR2x2_ASAP7_75t_L g5797 ( 
.A(n_5144),
.B(n_4545),
.Y(n_5797)
);

NAND2xp5_ASAP7_75t_L g5798 ( 
.A(n_5527),
.B(n_4915),
.Y(n_5798)
);

AO21x1_ASAP7_75t_SL g5799 ( 
.A1(n_5514),
.A2(n_5059),
.B(n_5040),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5176),
.Y(n_5800)
);

OR2x2_ASAP7_75t_L g5801 ( 
.A(n_5144),
.B(n_4545),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5606),
.Y(n_5802)
);

OR2x6_ASAP7_75t_L g5803 ( 
.A(n_5376),
.B(n_5459),
.Y(n_5803)
);

AND2x2_ASAP7_75t_L g5804 ( 
.A(n_5319),
.B(n_4802),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5326),
.B(n_4802),
.Y(n_5805)
);

AND2x2_ASAP7_75t_L g5806 ( 
.A(n_5377),
.B(n_4913),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5145),
.Y(n_5807)
);

INVx2_ASAP7_75t_L g5808 ( 
.A(n_5606),
.Y(n_5808)
);

HB1xp67_ASAP7_75t_L g5809 ( 
.A(n_5495),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5145),
.Y(n_5810)
);

INVx3_ASAP7_75t_L g5811 ( 
.A(n_5728),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_5423),
.Y(n_5812)
);

HB1xp67_ASAP7_75t_L g5813 ( 
.A(n_5504),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5146),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5146),
.Y(n_5815)
);

NAND2xp5_ASAP7_75t_L g5816 ( 
.A(n_5546),
.B(n_4459),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5214),
.Y(n_5817)
);

NOR2x1_ASAP7_75t_L g5818 ( 
.A(n_5124),
.B(n_4913),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5423),
.Y(n_5819)
);

OAI21x1_ASAP7_75t_L g5820 ( 
.A1(n_5728),
.A2(n_5005),
.B(n_4920),
.Y(n_5820)
);

HB1xp67_ASAP7_75t_L g5821 ( 
.A(n_5575),
.Y(n_5821)
);

INVx2_ASAP7_75t_SL g5822 ( 
.A(n_5175),
.Y(n_5822)
);

AND2x4_ASAP7_75t_L g5823 ( 
.A(n_5444),
.B(n_4623),
.Y(n_5823)
);

OR2x2_ASAP7_75t_L g5824 ( 
.A(n_5408),
.B(n_4627),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5377),
.B(n_4913),
.Y(n_5825)
);

INVx2_ASAP7_75t_L g5826 ( 
.A(n_5427),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_5427),
.Y(n_5827)
);

HB1xp67_ASAP7_75t_L g5828 ( 
.A(n_5201),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5206),
.Y(n_5829)
);

AND2x4_ASAP7_75t_L g5830 ( 
.A(n_5510),
.B(n_4623),
.Y(n_5830)
);

BUFx2_ASAP7_75t_L g5831 ( 
.A(n_5124),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5206),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5431),
.Y(n_5833)
);

BUFx6f_ASAP7_75t_L g5834 ( 
.A(n_5114),
.Y(n_5834)
);

HB1xp67_ASAP7_75t_L g5835 ( 
.A(n_5215),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5207),
.Y(n_5836)
);

NOR2xp33_ASAP7_75t_L g5837 ( 
.A(n_5175),
.B(n_4628),
.Y(n_5837)
);

INVx3_ASAP7_75t_L g5838 ( 
.A(n_5700),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5132),
.B(n_4459),
.Y(n_5839)
);

INVx1_ASAP7_75t_L g5840 ( 
.A(n_5172),
.Y(n_5840)
);

OAI21x1_ASAP7_75t_L g5841 ( 
.A1(n_5700),
.A2(n_5024),
.B(n_5011),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5172),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5210),
.Y(n_5843)
);

AOI21x1_ASAP7_75t_L g5844 ( 
.A1(n_5565),
.A2(n_5584),
.B(n_5592),
.Y(n_5844)
);

AND2x2_ASAP7_75t_L g5845 ( 
.A(n_5395),
.B(n_4921),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5431),
.Y(n_5846)
);

OAI221xp5_ASAP7_75t_L g5847 ( 
.A1(n_5163),
.A2(n_5036),
.B1(n_5066),
.B2(n_4532),
.C(n_5080),
.Y(n_5847)
);

INVx2_ASAP7_75t_SL g5848 ( 
.A(n_5175),
.Y(n_5848)
);

INVx2_ASAP7_75t_L g5849 ( 
.A(n_5433),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5211),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5211),
.Y(n_5851)
);

HB1xp67_ASAP7_75t_L g5852 ( 
.A(n_5235),
.Y(n_5852)
);

AOI21x1_ASAP7_75t_L g5853 ( 
.A1(n_5565),
.A2(n_4583),
.B(n_4516),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5395),
.B(n_4921),
.Y(n_5854)
);

INVx2_ASAP7_75t_L g5855 ( 
.A(n_5433),
.Y(n_5855)
);

OAI21x1_ASAP7_75t_L g5856 ( 
.A1(n_5549),
.A2(n_5024),
.B(n_5011),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5213),
.Y(n_5857)
);

AO21x2_ASAP7_75t_L g5858 ( 
.A1(n_5593),
.A2(n_5117),
.B(n_5365),
.Y(n_5858)
);

BUFx12f_ASAP7_75t_L g5859 ( 
.A(n_5165),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5593),
.Y(n_5860)
);

INVx2_ASAP7_75t_L g5861 ( 
.A(n_5346),
.Y(n_5861)
);

OAI22xp33_ASAP7_75t_L g5862 ( 
.A1(n_5372),
.A2(n_4520),
.B1(n_4844),
.B2(n_4945),
.Y(n_5862)
);

CKINVDCx20_ASAP7_75t_R g5863 ( 
.A(n_5345),
.Y(n_5863)
);

AO21x2_ASAP7_75t_L g5864 ( 
.A1(n_5117),
.A2(n_4761),
.B(n_4746),
.Y(n_5864)
);

OAI221xp5_ASAP7_75t_L g5865 ( 
.A1(n_5475),
.A2(n_5070),
.B1(n_4891),
.B2(n_4855),
.C(n_4845),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5346),
.Y(n_5866)
);

NOR2x1_ASAP7_75t_SL g5867 ( 
.A(n_5633),
.B(n_4982),
.Y(n_5867)
);

HB1xp67_ASAP7_75t_L g5868 ( 
.A(n_5249),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5349),
.Y(n_5869)
);

HB1xp67_ASAP7_75t_L g5870 ( 
.A(n_5270),
.Y(n_5870)
);

INVx3_ASAP7_75t_L g5871 ( 
.A(n_5375),
.Y(n_5871)
);

HB1xp67_ASAP7_75t_L g5872 ( 
.A(n_5273),
.Y(n_5872)
);

BUFx6f_ASAP7_75t_L g5873 ( 
.A(n_5114),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5120),
.Y(n_5874)
);

HB1xp67_ASAP7_75t_L g5875 ( 
.A(n_5275),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5120),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5153),
.Y(n_5877)
);

CKINVDCx8_ASAP7_75t_R g5878 ( 
.A(n_5165),
.Y(n_5878)
);

OA21x2_ASAP7_75t_L g5879 ( 
.A1(n_5484),
.A2(n_4761),
.B(n_4746),
.Y(n_5879)
);

NAND2xp5_ASAP7_75t_L g5880 ( 
.A(n_5414),
.B(n_4475),
.Y(n_5880)
);

NAND2xp5_ASAP7_75t_L g5881 ( 
.A(n_5390),
.B(n_4475),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5274),
.Y(n_5882)
);

AOI21xp5_ASAP7_75t_SL g5883 ( 
.A1(n_5192),
.A2(n_4933),
.B(n_4849),
.Y(n_5883)
);

INVx2_ASAP7_75t_L g5884 ( 
.A(n_5349),
.Y(n_5884)
);

INVx2_ASAP7_75t_SL g5885 ( 
.A(n_5175),
.Y(n_5885)
);

BUFx2_ASAP7_75t_L g5886 ( 
.A(n_5124),
.Y(n_5886)
);

AO21x1_ASAP7_75t_SL g5887 ( 
.A1(n_5372),
.A2(n_5059),
.B(n_5040),
.Y(n_5887)
);

INVx2_ASAP7_75t_L g5888 ( 
.A(n_5353),
.Y(n_5888)
);

OA21x2_ASAP7_75t_L g5889 ( 
.A1(n_5484),
.A2(n_4768),
.B(n_4765),
.Y(n_5889)
);

NAND2xp5_ASAP7_75t_L g5890 ( 
.A(n_5238),
.B(n_4480),
.Y(n_5890)
);

INVx2_ASAP7_75t_L g5891 ( 
.A(n_5353),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5156),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5156),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5190),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5356),
.Y(n_5895)
);

OAI21x1_ASAP7_75t_L g5896 ( 
.A1(n_5549),
.A2(n_4831),
.B(n_4827),
.Y(n_5896)
);

OR2x2_ASAP7_75t_L g5897 ( 
.A(n_5408),
.B(n_4627),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5210),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5213),
.Y(n_5899)
);

AOI21xp5_ASAP7_75t_SL g5900 ( 
.A1(n_5192),
.A2(n_4933),
.B(n_4399),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5254),
.Y(n_5901)
);

BUFx2_ASAP7_75t_L g5902 ( 
.A(n_5187),
.Y(n_5902)
);

OR2x2_ASAP7_75t_L g5903 ( 
.A(n_5110),
.B(n_4668),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5254),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5400),
.B(n_4921),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5400),
.B(n_4980),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5356),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5274),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5284),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5686),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5686),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_L g5912 ( 
.A(n_5246),
.B(n_4480),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5359),
.Y(n_5913)
);

INVx2_ASAP7_75t_L g5914 ( 
.A(n_5686),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5359),
.Y(n_5915)
);

INVx3_ASAP7_75t_L g5916 ( 
.A(n_5375),
.Y(n_5916)
);

OR2x2_ASAP7_75t_L g5917 ( 
.A(n_5110),
.B(n_4813),
.Y(n_5917)
);

NOR2x1_ASAP7_75t_R g5918 ( 
.A(n_5554),
.B(n_4926),
.Y(n_5918)
);

OR2x2_ASAP7_75t_L g5919 ( 
.A(n_5413),
.B(n_4826),
.Y(n_5919)
);

AND2x2_ASAP7_75t_L g5920 ( 
.A(n_5412),
.B(n_4980),
.Y(n_5920)
);

INVxp67_ASAP7_75t_L g5921 ( 
.A(n_5264),
.Y(n_5921)
);

INVx3_ASAP7_75t_L g5922 ( 
.A(n_5375),
.Y(n_5922)
);

INVx2_ASAP7_75t_L g5923 ( 
.A(n_5701),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5227),
.Y(n_5924)
);

BUFx3_ASAP7_75t_L g5925 ( 
.A(n_5554),
.Y(n_5925)
);

OAI21xp5_ASAP7_75t_L g5926 ( 
.A1(n_5296),
.A2(n_5104),
.B(n_5028),
.Y(n_5926)
);

OAI21x1_ASAP7_75t_L g5927 ( 
.A1(n_5705),
.A2(n_4831),
.B(n_4827),
.Y(n_5927)
);

AND2x2_ASAP7_75t_L g5928 ( 
.A(n_5412),
.B(n_4980),
.Y(n_5928)
);

OR2x2_ASAP7_75t_L g5929 ( 
.A(n_5413),
.B(n_4630),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5701),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5227),
.Y(n_5931)
);

INVx2_ASAP7_75t_L g5932 ( 
.A(n_5701),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5248),
.Y(n_5933)
);

HB1xp67_ASAP7_75t_L g5934 ( 
.A(n_5327),
.Y(n_5934)
);

AO21x2_ASAP7_75t_L g5935 ( 
.A1(n_5365),
.A2(n_4768),
.B(n_4765),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5502),
.Y(n_5936)
);

HB1xp67_ASAP7_75t_L g5937 ( 
.A(n_5378),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5502),
.Y(n_5938)
);

OR2x2_ASAP7_75t_L g5939 ( 
.A(n_5220),
.B(n_4630),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5248),
.Y(n_5940)
);

AND2x2_ASAP7_75t_L g5941 ( 
.A(n_5416),
.B(n_4991),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5250),
.Y(n_5942)
);

OR2x6_ASAP7_75t_L g5943 ( 
.A(n_5376),
.B(n_5459),
.Y(n_5943)
);

BUFx6f_ASAP7_75t_L g5944 ( 
.A(n_5165),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5250),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5416),
.B(n_4991),
.Y(n_5946)
);

OAI21x1_ASAP7_75t_L g5947 ( 
.A1(n_5705),
.A2(n_4831),
.B(n_4827),
.Y(n_5947)
);

OR2x2_ASAP7_75t_L g5948 ( 
.A(n_5220),
.B(n_4553),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5112),
.B(n_4991),
.Y(n_5949)
);

HB1xp67_ASAP7_75t_L g5950 ( 
.A(n_5389),
.Y(n_5950)
);

INVx2_ASAP7_75t_L g5951 ( 
.A(n_5505),
.Y(n_5951)
);

OR2x2_ASAP7_75t_L g5952 ( 
.A(n_5142),
.B(n_4451),
.Y(n_5952)
);

AO21x2_ASAP7_75t_L g5953 ( 
.A1(n_5367),
.A2(n_4768),
.B(n_4765),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5194),
.Y(n_5954)
);

BUFx3_ASAP7_75t_L g5955 ( 
.A(n_5264),
.Y(n_5955)
);

HB1xp67_ASAP7_75t_L g5956 ( 
.A(n_5399),
.Y(n_5956)
);

BUFx3_ASAP7_75t_L g5957 ( 
.A(n_5175),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5195),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5505),
.Y(n_5959)
);

INVx2_ASAP7_75t_L g5960 ( 
.A(n_5545),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_L g5961 ( 
.A(n_5255),
.B(n_4747),
.Y(n_5961)
);

HB1xp67_ASAP7_75t_L g5962 ( 
.A(n_5410),
.Y(n_5962)
);

BUFx2_ASAP7_75t_L g5963 ( 
.A(n_5187),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5112),
.B(n_5048),
.Y(n_5964)
);

AO21x2_ASAP7_75t_L g5965 ( 
.A1(n_5367),
.A2(n_4776),
.B(n_4839),
.Y(n_5965)
);

BUFx2_ASAP7_75t_L g5966 ( 
.A(n_5187),
.Y(n_5966)
);

INVx2_ASAP7_75t_L g5967 ( 
.A(n_5545),
.Y(n_5967)
);

AO21x2_ASAP7_75t_L g5968 ( 
.A1(n_5368),
.A2(n_4776),
.B(n_5013),
.Y(n_5968)
);

AO21x1_ASAP7_75t_SL g5969 ( 
.A1(n_5528),
.A2(n_4844),
.B(n_4422),
.Y(n_5969)
);

OR2x6_ASAP7_75t_L g5970 ( 
.A(n_5376),
.B(n_4899),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5118),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5545),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5118),
.Y(n_5973)
);

AO21x2_ASAP7_75t_L g5974 ( 
.A1(n_5368),
.A2(n_5382),
.B(n_5370),
.Y(n_5974)
);

INVx2_ASAP7_75t_SL g5975 ( 
.A(n_5165),
.Y(n_5975)
);

INVx2_ASAP7_75t_L g5976 ( 
.A(n_5545),
.Y(n_5976)
);

AND2x2_ASAP7_75t_L g5977 ( 
.A(n_5115),
.B(n_5048),
.Y(n_5977)
);

AO21x2_ASAP7_75t_L g5978 ( 
.A1(n_5370),
.A2(n_4776),
.B(n_5085),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5109),
.Y(n_5979)
);

NAND2xp5_ASAP7_75t_L g5980 ( 
.A(n_5276),
.B(n_4747),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5128),
.Y(n_5981)
);

INVx2_ASAP7_75t_L g5982 ( 
.A(n_5109),
.Y(n_5982)
);

NOR2xp33_ASAP7_75t_L g5983 ( 
.A(n_5167),
.B(n_4632),
.Y(n_5983)
);

BUFx6f_ASAP7_75t_L g5984 ( 
.A(n_5167),
.Y(n_5984)
);

INVxp67_ASAP7_75t_SL g5985 ( 
.A(n_5138),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5128),
.Y(n_5986)
);

AND2x4_ASAP7_75t_L g5987 ( 
.A(n_5510),
.B(n_4911),
.Y(n_5987)
);

INVx2_ASAP7_75t_L g5988 ( 
.A(n_5113),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5136),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5136),
.Y(n_5990)
);

OA21x2_ASAP7_75t_L g5991 ( 
.A1(n_5566),
.A2(n_4614),
.B(n_4587),
.Y(n_5991)
);

INVx2_ASAP7_75t_L g5992 ( 
.A(n_5113),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5169),
.Y(n_5993)
);

INVx2_ASAP7_75t_L g5994 ( 
.A(n_5122),
.Y(n_5994)
);

BUFx3_ASAP7_75t_L g5995 ( 
.A(n_5167),
.Y(n_5995)
);

OR2x6_ASAP7_75t_L g5996 ( 
.A(n_5459),
.B(n_4842),
.Y(n_5996)
);

BUFx2_ASAP7_75t_L g5997 ( 
.A(n_5265),
.Y(n_5997)
);

OR2x2_ASAP7_75t_L g5998 ( 
.A(n_5419),
.B(n_4451),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5122),
.Y(n_5999)
);

INVx2_ASAP7_75t_L g6000 ( 
.A(n_5125),
.Y(n_6000)
);

OAI21x1_ASAP7_75t_L g6001 ( 
.A1(n_5715),
.A2(n_4857),
.B(n_4836),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5115),
.B(n_5048),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5121),
.B(n_4834),
.Y(n_6003)
);

INVx2_ASAP7_75t_SL g6004 ( 
.A(n_5167),
.Y(n_6004)
);

AO21x2_ASAP7_75t_L g6005 ( 
.A1(n_5382),
.A2(n_4857),
.B(n_4836),
.Y(n_6005)
);

AO21x2_ASAP7_75t_L g6006 ( 
.A1(n_5383),
.A2(n_4857),
.B(n_4836),
.Y(n_6006)
);

CKINVDCx20_ASAP7_75t_R g6007 ( 
.A(n_5311),
.Y(n_6007)
);

OR2x2_ASAP7_75t_L g6008 ( 
.A(n_5419),
.B(n_4533),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5169),
.Y(n_6009)
);

OR2x6_ASAP7_75t_L g6010 ( 
.A(n_5537),
.B(n_5014),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5176),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5125),
.Y(n_6012)
);

NAND2xp5_ASAP7_75t_SL g6013 ( 
.A(n_5612),
.B(n_4465),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5185),
.Y(n_6014)
);

CKINVDCx14_ASAP7_75t_R g6015 ( 
.A(n_5652),
.Y(n_6015)
);

NOR2xp33_ASAP7_75t_L g6016 ( 
.A(n_5167),
.B(n_4960),
.Y(n_6016)
);

BUFx2_ASAP7_75t_L g6017 ( 
.A(n_5265),
.Y(n_6017)
);

OR2x2_ASAP7_75t_L g6018 ( 
.A(n_5452),
.B(n_4533),
.Y(n_6018)
);

INVxp67_ASAP7_75t_L g6019 ( 
.A(n_5111),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5127),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5127),
.Y(n_6021)
);

NOR2xp33_ASAP7_75t_L g6022 ( 
.A(n_5342),
.B(n_4708),
.Y(n_6022)
);

AOI22xp33_ASAP7_75t_L g6023 ( 
.A1(n_5647),
.A2(n_4464),
.B1(n_4520),
.B2(n_4881),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5185),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5194),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5195),
.Y(n_6026)
);

BUFx2_ASAP7_75t_L g6027 ( 
.A(n_5265),
.Y(n_6027)
);

BUFx2_ASAP7_75t_L g6028 ( 
.A(n_5226),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5130),
.Y(n_6029)
);

OA21x2_ASAP7_75t_L g6030 ( 
.A1(n_5566),
.A2(n_4614),
.B(n_4587),
.Y(n_6030)
);

OAI21x1_ASAP7_75t_L g6031 ( 
.A1(n_5715),
.A2(n_4900),
.B(n_4882),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5203),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5203),
.Y(n_6033)
);

INVx3_ASAP7_75t_SL g6034 ( 
.A(n_5221),
.Y(n_6034)
);

AND2x4_ASAP7_75t_L g6035 ( 
.A(n_5512),
.B(n_4623),
.Y(n_6035)
);

INVx2_ASAP7_75t_L g6036 ( 
.A(n_5130),
.Y(n_6036)
);

NOR2xp33_ASAP7_75t_L g6037 ( 
.A(n_5342),
.B(n_5580),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5209),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5121),
.B(n_5166),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5209),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5214),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5223),
.Y(n_6042)
);

OR2x2_ASAP7_75t_L g6043 ( 
.A(n_5452),
.B(n_4535),
.Y(n_6043)
);

INVx2_ASAP7_75t_L g6044 ( 
.A(n_5131),
.Y(n_6044)
);

OA21x2_ASAP7_75t_L g6045 ( 
.A1(n_5634),
.A2(n_4617),
.B(n_4614),
.Y(n_6045)
);

INVx4_ASAP7_75t_L g6046 ( 
.A(n_5200),
.Y(n_6046)
);

INVx2_ASAP7_75t_L g6047 ( 
.A(n_5131),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5134),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5134),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5137),
.Y(n_6050)
);

OAI21xp5_ASAP7_75t_L g6051 ( 
.A1(n_5337),
.A2(n_4727),
.B(n_4583),
.Y(n_6051)
);

OR2x2_ASAP7_75t_L g6052 ( 
.A(n_5507),
.B(n_4535),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5223),
.Y(n_6053)
);

BUFx6f_ASAP7_75t_L g6054 ( 
.A(n_5310),
.Y(n_6054)
);

AO21x2_ASAP7_75t_L g6055 ( 
.A1(n_5383),
.A2(n_4919),
.B(n_4900),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5231),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5231),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5137),
.Y(n_6058)
);

INVxp67_ASAP7_75t_SL g6059 ( 
.A(n_5138),
.Y(n_6059)
);

OAI21xp5_ASAP7_75t_L g6060 ( 
.A1(n_5138),
.A2(n_4727),
.B(n_4693),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5232),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5232),
.Y(n_6062)
);

HB1xp67_ASAP7_75t_L g6063 ( 
.A(n_5417),
.Y(n_6063)
);

INVx3_ASAP7_75t_L g6064 ( 
.A(n_5375),
.Y(n_6064)
);

INVx3_ASAP7_75t_L g6065 ( 
.A(n_5430),
.Y(n_6065)
);

OR2x6_ASAP7_75t_L g6066 ( 
.A(n_5537),
.B(n_4899),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5233),
.Y(n_6067)
);

OA21x2_ASAP7_75t_L g6068 ( 
.A1(n_5634),
.A2(n_4617),
.B(n_4481),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_5166),
.B(n_4856),
.Y(n_6069)
);

NAND2xp5_ASAP7_75t_L g6070 ( 
.A(n_5454),
.B(n_4516),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_5233),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5247),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5247),
.Y(n_6073)
);

AND2x2_ASAP7_75t_L g6074 ( 
.A(n_5173),
.B(n_4856),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_5279),
.Y(n_6075)
);

OR2x2_ASAP7_75t_L g6076 ( 
.A(n_5507),
.B(n_5302),
.Y(n_6076)
);

INVxp67_ASAP7_75t_L g6077 ( 
.A(n_5111),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5279),
.Y(n_6078)
);

INVxp67_ASAP7_75t_R g6079 ( 
.A(n_5129),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5282),
.Y(n_6080)
);

INVx2_ASAP7_75t_L g6081 ( 
.A(n_5139),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5173),
.B(n_4976),
.Y(n_6082)
);

AND2x2_ASAP7_75t_L g6083 ( 
.A(n_5177),
.B(n_4976),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5139),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5282),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5177),
.B(n_4977),
.Y(n_6086)
);

INVxp67_ASAP7_75t_SL g6087 ( 
.A(n_5138),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5283),
.Y(n_6088)
);

INVx3_ASAP7_75t_L g6089 ( 
.A(n_5430),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5283),
.Y(n_6090)
);

AO21x2_ASAP7_75t_L g6091 ( 
.A1(n_5391),
.A2(n_4900),
.B(n_4882),
.Y(n_6091)
);

INVxp67_ASAP7_75t_L g6092 ( 
.A(n_5147),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5284),
.Y(n_6093)
);

INVx1_ASAP7_75t_SL g6094 ( 
.A(n_5474),
.Y(n_6094)
);

BUFx6f_ASAP7_75t_L g6095 ( 
.A(n_5310),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5288),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5288),
.Y(n_6097)
);

OA21x2_ASAP7_75t_L g6098 ( 
.A1(n_5429),
.A2(n_4617),
.B(n_4481),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5140),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5292),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_5292),
.Y(n_6101)
);

INVx6_ASAP7_75t_L g6102 ( 
.A(n_5425),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_5297),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5297),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_5140),
.Y(n_6105)
);

HB1xp67_ASAP7_75t_L g6106 ( 
.A(n_5465),
.Y(n_6106)
);

OR2x2_ASAP7_75t_L g6107 ( 
.A(n_5302),
.B(n_4565),
.Y(n_6107)
);

OAI21x1_ASAP7_75t_L g6108 ( 
.A1(n_5726),
.A2(n_4919),
.B(n_4882),
.Y(n_6108)
);

INVx2_ASAP7_75t_L g6109 ( 
.A(n_5151),
.Y(n_6109)
);

INVx3_ASAP7_75t_L g6110 ( 
.A(n_5430),
.Y(n_6110)
);

BUFx2_ASAP7_75t_L g6111 ( 
.A(n_5492),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_5303),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5303),
.Y(n_6113)
);

INVx2_ASAP7_75t_L g6114 ( 
.A(n_5151),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_5486),
.B(n_4693),
.Y(n_6115)
);

OA21x2_ASAP7_75t_L g6116 ( 
.A1(n_5429),
.A2(n_4482),
.B(n_4479),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5164),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5304),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5304),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_5164),
.Y(n_6120)
);

AND2x2_ASAP7_75t_L g6121 ( 
.A(n_5181),
.B(n_4977),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5305),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5305),
.Y(n_6123)
);

HB1xp67_ASAP7_75t_L g6124 ( 
.A(n_5623),
.Y(n_6124)
);

OA21x2_ASAP7_75t_L g6125 ( 
.A1(n_5224),
.A2(n_4482),
.B(n_4479),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5308),
.Y(n_6126)
);

INVx4_ASAP7_75t_L g6127 ( 
.A(n_5200),
.Y(n_6127)
);

AND2x4_ASAP7_75t_L g6128 ( 
.A(n_5512),
.B(n_4623),
.Y(n_6128)
);

INVx2_ASAP7_75t_L g6129 ( 
.A(n_5178),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5308),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5315),
.Y(n_6131)
);

INVx2_ASAP7_75t_SL g6132 ( 
.A(n_5200),
.Y(n_6132)
);

INVxp67_ASAP7_75t_L g6133 ( 
.A(n_5147),
.Y(n_6133)
);

OAI21x1_ASAP7_75t_L g6134 ( 
.A1(n_5726),
.A2(n_4929),
.B(n_4919),
.Y(n_6134)
);

BUFx2_ASAP7_75t_L g6135 ( 
.A(n_5584),
.Y(n_6135)
);

AO21x2_ASAP7_75t_L g6136 ( 
.A1(n_5391),
.A2(n_4946),
.B(n_4929),
.Y(n_6136)
);

INVx2_ASAP7_75t_L g6137 ( 
.A(n_5178),
.Y(n_6137)
);

INVx3_ASAP7_75t_L g6138 ( 
.A(n_5430),
.Y(n_6138)
);

HB1xp67_ASAP7_75t_L g6139 ( 
.A(n_5659),
.Y(n_6139)
);

BUFx4f_ASAP7_75t_SL g6140 ( 
.A(n_5613),
.Y(n_6140)
);

BUFx2_ASAP7_75t_L g6141 ( 
.A(n_5148),
.Y(n_6141)
);

INVx2_ASAP7_75t_L g6142 ( 
.A(n_5179),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5315),
.Y(n_6143)
);

HB1xp67_ASAP7_75t_L g6144 ( 
.A(n_5723),
.Y(n_6144)
);

AND2x2_ASAP7_75t_L g6145 ( 
.A(n_5181),
.B(n_5025),
.Y(n_6145)
);

OAI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_5709),
.A2(n_4738),
.B(n_4945),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_5179),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5320),
.Y(n_6148)
);

OA21x2_ASAP7_75t_L g6149 ( 
.A1(n_5224),
.A2(n_4486),
.B(n_4618),
.Y(n_6149)
);

OR2x2_ASAP7_75t_L g6150 ( 
.A(n_5396),
.B(n_5405),
.Y(n_6150)
);

AO21x2_ASAP7_75t_L g6151 ( 
.A1(n_5394),
.A2(n_4946),
.B(n_4929),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_5183),
.Y(n_6152)
);

AO21x2_ASAP7_75t_L g6153 ( 
.A1(n_5394),
.A2(n_4946),
.B(n_4653),
.Y(n_6153)
);

OR2x2_ASAP7_75t_L g6154 ( 
.A(n_5396),
.B(n_4565),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_5320),
.Y(n_6155)
);

AND2x4_ASAP7_75t_L g6156 ( 
.A(n_5542),
.B(n_4911),
.Y(n_6156)
);

AO21x2_ASAP7_75t_L g6157 ( 
.A1(n_5397),
.A2(n_4653),
.B(n_4618),
.Y(n_6157)
);

OA21x2_ASAP7_75t_L g6158 ( 
.A1(n_5453),
.A2(n_4486),
.B(n_4618),
.Y(n_6158)
);

NAND2xp5_ASAP7_75t_L g6159 ( 
.A(n_5736),
.B(n_4738),
.Y(n_6159)
);

OR2x2_ASAP7_75t_L g6160 ( 
.A(n_5405),
.B(n_4833),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_5183),
.Y(n_6161)
);

INVx2_ASAP7_75t_SL g6162 ( 
.A(n_5200),
.Y(n_6162)
);

AND2x2_ASAP7_75t_L g6163 ( 
.A(n_5234),
.B(n_5025),
.Y(n_6163)
);

AND2x2_ASAP7_75t_L g6164 ( 
.A(n_5234),
.B(n_4842),
.Y(n_6164)
);

NAND2xp5_ASAP7_75t_SL g6165 ( 
.A(n_5542),
.B(n_4465),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5321),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5321),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5322),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_5322),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_5323),
.Y(n_6170)
);

OA21x2_ASAP7_75t_L g6171 ( 
.A1(n_5453),
.A2(n_4654),
.B(n_4653),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_5524),
.B(n_3981),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5323),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5324),
.Y(n_6174)
);

BUFx3_ASAP7_75t_L g6175 ( 
.A(n_5613),
.Y(n_6175)
);

OA21x2_ASAP7_75t_L g6176 ( 
.A1(n_5482),
.A2(n_4655),
.B(n_4654),
.Y(n_6176)
);

INVx2_ASAP7_75t_L g6177 ( 
.A(n_5184),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5324),
.Y(n_6178)
);

NAND2xp5_ASAP7_75t_L g6179 ( 
.A(n_5624),
.B(n_3981),
.Y(n_6179)
);

INVx2_ASAP7_75t_L g6180 ( 
.A(n_5184),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_5197),
.Y(n_6181)
);

INVx3_ASAP7_75t_SL g6182 ( 
.A(n_5197),
.Y(n_6182)
);

NAND3xp33_ASAP7_75t_L g6183 ( 
.A(n_5668),
.B(n_4797),
.C(n_4707),
.Y(n_6183)
);

BUFx8_ASAP7_75t_SL g6184 ( 
.A(n_5310),
.Y(n_6184)
);

AOI22xp33_ASAP7_75t_L g6185 ( 
.A1(n_5717),
.A2(n_4881),
.B1(n_4982),
.B2(n_4567),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5328),
.Y(n_6186)
);

INVx2_ASAP7_75t_L g6187 ( 
.A(n_5186),
.Y(n_6187)
);

BUFx3_ASAP7_75t_L g6188 ( 
.A(n_5636),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5328),
.Y(n_6189)
);

OA21x2_ASAP7_75t_L g6190 ( 
.A1(n_5482),
.A2(n_4655),
.B(n_4654),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5330),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_L g6192 ( 
.A(n_5649),
.B(n_3981),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5330),
.Y(n_6193)
);

OR2x6_ASAP7_75t_L g6194 ( 
.A(n_5537),
.B(n_5014),
.Y(n_6194)
);

OA21x2_ASAP7_75t_L g6195 ( 
.A1(n_5503),
.A2(n_4662),
.B(n_4655),
.Y(n_6195)
);

INVx2_ASAP7_75t_SL g6196 ( 
.A(n_5200),
.Y(n_6196)
);

AO21x2_ASAP7_75t_L g6197 ( 
.A1(n_5397),
.A2(n_5404),
.B(n_5398),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_5331),
.Y(n_6198)
);

AND2x2_ASAP7_75t_L g6199 ( 
.A(n_5291),
.B(n_5054),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_5291),
.B(n_5054),
.Y(n_6200)
);

OA21x2_ASAP7_75t_L g6201 ( 
.A1(n_5503),
.A2(n_4669),
.B(n_4662),
.Y(n_6201)
);

AO21x2_ASAP7_75t_L g6202 ( 
.A1(n_5398),
.A2(n_4669),
.B(n_4662),
.Y(n_6202)
);

AO21x2_ASAP7_75t_L g6203 ( 
.A1(n_5404),
.A2(n_4698),
.B(n_4669),
.Y(n_6203)
);

AO21x2_ASAP7_75t_L g6204 ( 
.A1(n_5418),
.A2(n_5485),
.B(n_5472),
.Y(n_6204)
);

INVx2_ASAP7_75t_L g6205 ( 
.A(n_5186),
.Y(n_6205)
);

INVx2_ASAP7_75t_L g6206 ( 
.A(n_5191),
.Y(n_6206)
);

OA21x2_ASAP7_75t_L g6207 ( 
.A1(n_5244),
.A2(n_4711),
.B(n_4698),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_5331),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5338),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_5191),
.Y(n_6210)
);

INVx1_ASAP7_75t_SL g6211 ( 
.A(n_5243),
.Y(n_6211)
);

INVx2_ASAP7_75t_L g6212 ( 
.A(n_5199),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_5338),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_5307),
.B(n_4608),
.Y(n_6214)
);

INVx2_ASAP7_75t_L g6215 ( 
.A(n_5199),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5341),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_5341),
.Y(n_6217)
);

AND2x2_ASAP7_75t_L g6218 ( 
.A(n_5307),
.B(n_5697),
.Y(n_6218)
);

OA21x2_ASAP7_75t_L g6219 ( 
.A1(n_5244),
.A2(n_4711),
.B(n_4698),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_5344),
.Y(n_6220)
);

INVx2_ASAP7_75t_L g6221 ( 
.A(n_5202),
.Y(n_6221)
);

NOR2xp33_ASAP7_75t_L g6222 ( 
.A(n_5339),
.B(n_4784),
.Y(n_6222)
);

INVx2_ASAP7_75t_L g6223 ( 
.A(n_5202),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_5204),
.Y(n_6224)
);

INVx3_ASAP7_75t_L g6225 ( 
.A(n_5464),
.Y(n_6225)
);

INVx3_ASAP7_75t_L g6226 ( 
.A(n_5464),
.Y(n_6226)
);

OR2x2_ASAP7_75t_L g6227 ( 
.A(n_5174),
.B(n_4833),
.Y(n_6227)
);

INVx1_ASAP7_75t_L g6228 ( 
.A(n_5344),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_5204),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5348),
.Y(n_6230)
);

OAI21xp5_ASAP7_75t_L g6231 ( 
.A1(n_5668),
.A2(n_4591),
.B(n_4843),
.Y(n_6231)
);

INVx2_ASAP7_75t_L g6232 ( 
.A(n_5217),
.Y(n_6232)
);

NAND2xp5_ASAP7_75t_L g6233 ( 
.A(n_5592),
.B(n_3981),
.Y(n_6233)
);

AND2x2_ASAP7_75t_L g6234 ( 
.A(n_5697),
.B(n_5703),
.Y(n_6234)
);

OAI21x1_ASAP7_75t_L g6235 ( 
.A1(n_5727),
.A2(n_5043),
.B(n_4962),
.Y(n_6235)
);

OR2x6_ASAP7_75t_L g6236 ( 
.A(n_5552),
.B(n_5558),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_5348),
.Y(n_6237)
);

HB1xp67_ASAP7_75t_L g6238 ( 
.A(n_5586),
.Y(n_6238)
);

AO21x2_ASAP7_75t_L g6239 ( 
.A1(n_5418),
.A2(n_4711),
.B(n_4881),
.Y(n_6239)
);

AO21x2_ASAP7_75t_L g6240 ( 
.A1(n_5472),
.A2(n_4990),
.B(n_4951),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5351),
.Y(n_6241)
);

OAI21xp5_ASAP7_75t_L g6242 ( 
.A1(n_5278),
.A2(n_4843),
.B(n_4858),
.Y(n_6242)
);

INVx1_ASAP7_75t_SL g6243 ( 
.A(n_5243),
.Y(n_6243)
);

HB1xp67_ASAP7_75t_L g6244 ( 
.A(n_5351),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5354),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_5354),
.Y(n_6246)
);

AOI21x1_ASAP7_75t_L g6247 ( 
.A1(n_5271),
.A2(n_4736),
.B(n_4608),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5217),
.Y(n_6248)
);

INVx2_ASAP7_75t_L g6249 ( 
.A(n_5222),
.Y(n_6249)
);

AO21x2_ASAP7_75t_L g6250 ( 
.A1(n_5485),
.A2(n_4990),
.B(n_4951),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5355),
.Y(n_6251)
);

AND2x2_ASAP7_75t_L g6252 ( 
.A(n_5703),
.B(n_4736),
.Y(n_6252)
);

NAND2x1p5_ASAP7_75t_L g6253 ( 
.A(n_5200),
.B(n_4688),
.Y(n_6253)
);

AO21x2_ASAP7_75t_L g6254 ( 
.A1(n_5489),
.A2(n_4990),
.B(n_4951),
.Y(n_6254)
);

INVx3_ASAP7_75t_L g6255 ( 
.A(n_5464),
.Y(n_6255)
);

INVx2_ASAP7_75t_L g6256 ( 
.A(n_5222),
.Y(n_6256)
);

BUFx2_ASAP7_75t_L g6257 ( 
.A(n_5148),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5355),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_5228),
.Y(n_6259)
);

AND2x4_ASAP7_75t_L g6260 ( 
.A(n_5803),
.B(n_5425),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_5921),
.B(n_5741),
.Y(n_6261)
);

CKINVDCx5p33_ASAP7_75t_R g6262 ( 
.A(n_5863),
.Y(n_6262)
);

INVx1_ASAP7_75t_SL g6263 ( 
.A(n_5863),
.Y(n_6263)
);

AND2x2_ASAP7_75t_L g6264 ( 
.A(n_5769),
.B(n_5529),
.Y(n_6264)
);

AND2x2_ASAP7_75t_L g6265 ( 
.A(n_5769),
.B(n_5529),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_6244),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5744),
.Y(n_6267)
);

AO21x2_ASAP7_75t_L g6268 ( 
.A1(n_5985),
.A2(n_5699),
.B(n_5445),
.Y(n_6268)
);

NAND2xp5_ASAP7_75t_L g6269 ( 
.A(n_6019),
.B(n_5541),
.Y(n_6269)
);

NOR2xp33_ASAP7_75t_SL g6270 ( 
.A(n_5766),
.B(n_5317),
.Y(n_6270)
);

AND2x2_ASAP7_75t_L g6271 ( 
.A(n_5770),
.B(n_5529),
.Y(n_6271)
);

HB1xp67_ASAP7_75t_L g6272 ( 
.A(n_6077),
.Y(n_6272)
);

INVx2_ASAP7_75t_L g6273 ( 
.A(n_5790),
.Y(n_6273)
);

NAND2xp5_ASAP7_75t_L g6274 ( 
.A(n_6092),
.B(n_5541),
.Y(n_6274)
);

INVx2_ASAP7_75t_SL g6275 ( 
.A(n_6102),
.Y(n_6275)
);

AND2x2_ASAP7_75t_L g6276 ( 
.A(n_6111),
.B(n_5126),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_5790),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_5790),
.Y(n_6278)
);

AND2x2_ASAP7_75t_L g6279 ( 
.A(n_6111),
.B(n_5126),
.Y(n_6279)
);

BUFx3_ASAP7_75t_L g6280 ( 
.A(n_5766),
.Y(n_6280)
);

OR2x2_ASAP7_75t_L g6281 ( 
.A(n_6076),
.B(n_6150),
.Y(n_6281)
);

AND2x2_ASAP7_75t_L g6282 ( 
.A(n_5770),
.B(n_5774),
.Y(n_6282)
);

NAND2x1_ASAP7_75t_L g6283 ( 
.A(n_6065),
.B(n_5582),
.Y(n_6283)
);

AND2x2_ASAP7_75t_L g6284 ( 
.A(n_5774),
.B(n_5126),
.Y(n_6284)
);

AND2x2_ASAP7_75t_L g6285 ( 
.A(n_5779),
.B(n_5126),
.Y(n_6285)
);

BUFx6f_ASAP7_75t_L g6286 ( 
.A(n_6175),
.Y(n_6286)
);

BUFx3_ASAP7_75t_L g6287 ( 
.A(n_6188),
.Y(n_6287)
);

INVxp67_ASAP7_75t_SL g6288 ( 
.A(n_6059),
.Y(n_6288)
);

BUFx2_ASAP7_75t_L g6289 ( 
.A(n_6015),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_5791),
.Y(n_6290)
);

NAND2xp5_ASAP7_75t_L g6291 ( 
.A(n_6133),
.B(n_5574),
.Y(n_6291)
);

AND2x2_ASAP7_75t_SL g6292 ( 
.A(n_6028),
.B(n_5373),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_5740),
.Y(n_6293)
);

AND2x4_ASAP7_75t_L g6294 ( 
.A(n_5803),
.B(n_5425),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_5779),
.B(n_5126),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_6234),
.B(n_5129),
.Y(n_6296)
);

OR2x2_ASAP7_75t_L g6297 ( 
.A(n_6076),
.B(n_5620),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6234),
.B(n_5129),
.Y(n_6298)
);

AND2x2_ASAP7_75t_L g6299 ( 
.A(n_5955),
.B(n_6252),
.Y(n_6299)
);

AND2x4_ASAP7_75t_SL g6300 ( 
.A(n_5944),
.B(n_5615),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5746),
.Y(n_6301)
);

INVx3_ASAP7_75t_L g6302 ( 
.A(n_5772),
.Y(n_6302)
);

OR2x2_ASAP7_75t_L g6303 ( 
.A(n_6150),
.B(n_5534),
.Y(n_6303)
);

NAND2xp5_ASAP7_75t_L g6304 ( 
.A(n_5955),
.B(n_5781),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_5791),
.Y(n_6305)
);

BUFx3_ASAP7_75t_L g6306 ( 
.A(n_6188),
.Y(n_6306)
);

NAND2xp5_ASAP7_75t_L g6307 ( 
.A(n_5794),
.B(n_5574),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5747),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5748),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_6252),
.B(n_5129),
.Y(n_6310)
);

AND2x4_ASAP7_75t_L g6311 ( 
.A(n_5803),
.B(n_5425),
.Y(n_6311)
);

AND2x2_ASAP7_75t_L g6312 ( 
.A(n_5949),
.B(n_5437),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5749),
.Y(n_6313)
);

AND2x2_ASAP7_75t_L g6314 ( 
.A(n_5949),
.B(n_5437),
.Y(n_6314)
);

HB1xp67_ASAP7_75t_L g6315 ( 
.A(n_5809),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_5753),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_5754),
.Y(n_6317)
);

OR2x2_ASAP7_75t_L g6318 ( 
.A(n_5787),
.B(n_5775),
.Y(n_6318)
);

AND2x4_ASAP7_75t_L g6319 ( 
.A(n_5803),
.B(n_5552),
.Y(n_6319)
);

INVx2_ASAP7_75t_SL g6320 ( 
.A(n_6102),
.Y(n_6320)
);

AND2x2_ASAP7_75t_L g6321 ( 
.A(n_5964),
.B(n_5449),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_5791),
.Y(n_6322)
);

INVx2_ASAP7_75t_R g6323 ( 
.A(n_5925),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_5757),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5758),
.Y(n_6325)
);

INVxp67_ASAP7_75t_SL g6326 ( 
.A(n_6087),
.Y(n_6326)
);

INVx2_ASAP7_75t_L g6327 ( 
.A(n_5858),
.Y(n_6327)
);

AND2x2_ASAP7_75t_L g6328 ( 
.A(n_5964),
.B(n_5449),
.Y(n_6328)
);

AND2x2_ASAP7_75t_L g6329 ( 
.A(n_5977),
.B(n_5508),
.Y(n_6329)
);

INVx2_ASAP7_75t_R g6330 ( 
.A(n_5925),
.Y(n_6330)
);

NOR2xp67_ASAP7_75t_L g6331 ( 
.A(n_5752),
.B(n_5645),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_5759),
.Y(n_6332)
);

AND2x2_ASAP7_75t_L g6333 ( 
.A(n_5977),
.B(n_5508),
.Y(n_6333)
);

INVx2_ASAP7_75t_L g6334 ( 
.A(n_5858),
.Y(n_6334)
);

BUFx3_ASAP7_75t_L g6335 ( 
.A(n_6007),
.Y(n_6335)
);

OR2x6_ASAP7_75t_L g6336 ( 
.A(n_6102),
.B(n_5552),
.Y(n_6336)
);

AND2x4_ASAP7_75t_L g6337 ( 
.A(n_5943),
.B(n_5558),
.Y(n_6337)
);

AOI21xp5_ASAP7_75t_L g6338 ( 
.A1(n_5883),
.A2(n_5699),
.B(n_5561),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_5858),
.Y(n_6339)
);

AND2x2_ASAP7_75t_L g6340 ( 
.A(n_6002),
.B(n_5529),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_5760),
.Y(n_6341)
);

AOI22xp33_ASAP7_75t_L g6342 ( 
.A1(n_6023),
.A2(n_5689),
.B1(n_5133),
.B2(n_5229),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_5763),
.Y(n_6343)
);

INVx3_ASAP7_75t_L g6344 ( 
.A(n_5772),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_6002),
.B(n_5563),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_5765),
.Y(n_6346)
);

AND2x2_ASAP7_75t_L g6347 ( 
.A(n_5804),
.B(n_5563),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_5771),
.Y(n_6348)
);

AND2x4_ASAP7_75t_L g6349 ( 
.A(n_5943),
.B(n_5558),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_5738),
.Y(n_6350)
);

OAI22xp5_ASAP7_75t_L g6351 ( 
.A1(n_6183),
.A2(n_5281),
.B1(n_5219),
.B2(n_5205),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_5782),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_5738),
.Y(n_6353)
);

OR2x2_ASAP7_75t_L g6354 ( 
.A(n_5787),
.B(n_5775),
.Y(n_6354)
);

AND2x2_ASAP7_75t_L g6355 ( 
.A(n_5804),
.B(n_5805),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_5805),
.B(n_5373),
.Y(n_6356)
);

AND2x2_ASAP7_75t_L g6357 ( 
.A(n_5806),
.B(n_5373),
.Y(n_6357)
);

OR2x2_ASAP7_75t_L g6358 ( 
.A(n_5776),
.B(n_5534),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_5738),
.Y(n_6359)
);

INVx4_ASAP7_75t_L g6360 ( 
.A(n_6140),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5784),
.Y(n_6361)
);

INVx2_ASAP7_75t_L g6362 ( 
.A(n_5761),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_5806),
.B(n_5373),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_5786),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_5800),
.Y(n_6365)
);

AND2x2_ASAP7_75t_L g6366 ( 
.A(n_5825),
.B(n_5208),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_5761),
.Y(n_6367)
);

NOR2xp33_ASAP7_75t_L g6368 ( 
.A(n_6015),
.B(n_5339),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_5761),
.Y(n_6369)
);

INVx2_ASAP7_75t_L g6370 ( 
.A(n_5864),
.Y(n_6370)
);

AND2x2_ASAP7_75t_L g6371 ( 
.A(n_5825),
.B(n_5208),
.Y(n_6371)
);

HB1xp67_ASAP7_75t_L g6372 ( 
.A(n_5813),
.Y(n_6372)
);

BUFx3_ASAP7_75t_L g6373 ( 
.A(n_6007),
.Y(n_6373)
);

HB1xp67_ASAP7_75t_L g6374 ( 
.A(n_5821),
.Y(n_6374)
);

AND2x2_ASAP7_75t_L g6375 ( 
.A(n_5845),
.B(n_5615),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_5807),
.Y(n_6376)
);

AND2x4_ASAP7_75t_L g6377 ( 
.A(n_5943),
.B(n_5588),
.Y(n_6377)
);

AND2x2_ASAP7_75t_L g6378 ( 
.A(n_5845),
.B(n_5148),
.Y(n_6378)
);

AND2x2_ASAP7_75t_L g6379 ( 
.A(n_5854),
.B(n_5148),
.Y(n_6379)
);

NOR2xp33_ASAP7_75t_L g6380 ( 
.A(n_6034),
.B(n_5339),
.Y(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_5854),
.B(n_5148),
.Y(n_6381)
);

NAND2xp5_ASAP7_75t_L g6382 ( 
.A(n_5828),
.B(n_5579),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_5810),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_5905),
.B(n_5154),
.Y(n_6384)
);

OR2x2_ASAP7_75t_L g6385 ( 
.A(n_5776),
.B(n_5174),
.Y(n_6385)
);

INVx2_ASAP7_75t_L g6386 ( 
.A(n_5864),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_5814),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5815),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_5864),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_5817),
.Y(n_6390)
);

INVx2_ASAP7_75t_L g6391 ( 
.A(n_6240),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_6240),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_5835),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_5829),
.Y(n_6394)
);

HB1xp67_ASAP7_75t_L g6395 ( 
.A(n_5852),
.Y(n_6395)
);

BUFx3_ASAP7_75t_L g6396 ( 
.A(n_5755),
.Y(n_6396)
);

INVx2_ASAP7_75t_SL g6397 ( 
.A(n_6102),
.Y(n_6397)
);

INVx2_ASAP7_75t_L g6398 ( 
.A(n_6240),
.Y(n_6398)
);

INVx2_ASAP7_75t_L g6399 ( 
.A(n_6250),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_5832),
.Y(n_6400)
);

AND2x4_ASAP7_75t_L g6401 ( 
.A(n_5943),
.B(n_5588),
.Y(n_6401)
);

BUFx2_ASAP7_75t_L g6402 ( 
.A(n_6028),
.Y(n_6402)
);

INVxp67_ASAP7_75t_SL g6403 ( 
.A(n_5811),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_5868),
.B(n_5579),
.Y(n_6404)
);

INVx2_ASAP7_75t_L g6405 ( 
.A(n_6250),
.Y(n_6405)
);

INVx2_ASAP7_75t_L g6406 ( 
.A(n_6250),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_5905),
.B(n_5154),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5836),
.Y(n_6408)
);

AND2x2_ASAP7_75t_L g6409 ( 
.A(n_5906),
.B(n_5563),
.Y(n_6409)
);

INVx2_ASAP7_75t_L g6410 ( 
.A(n_6254),
.Y(n_6410)
);

AOI22xp33_ASAP7_75t_L g6411 ( 
.A1(n_5788),
.A2(n_5133),
.B1(n_5229),
.B2(n_4368),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_6254),
.Y(n_6412)
);

INVx1_ASAP7_75t_SL g6413 ( 
.A(n_6182),
.Y(n_6413)
);

AND2x2_ASAP7_75t_L g6414 ( 
.A(n_5906),
.B(n_5563),
.Y(n_6414)
);

AND2x2_ASAP7_75t_L g6415 ( 
.A(n_5920),
.B(n_5568),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5840),
.Y(n_6416)
);

INVx2_ASAP7_75t_SL g6417 ( 
.A(n_5944),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6254),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_5870),
.B(n_5154),
.Y(n_6419)
);

AOI22xp33_ASAP7_75t_L g6420 ( 
.A1(n_5737),
.A2(n_5133),
.B1(n_5229),
.B2(n_5588),
.Y(n_6420)
);

INVx2_ASAP7_75t_L g6421 ( 
.A(n_5974),
.Y(n_6421)
);

AND2x2_ASAP7_75t_L g6422 ( 
.A(n_5920),
.B(n_5568),
.Y(n_6422)
);

NOR2xp33_ASAP7_75t_L g6423 ( 
.A(n_6034),
.B(n_6182),
.Y(n_6423)
);

INVx2_ASAP7_75t_L g6424 ( 
.A(n_5974),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_5928),
.B(n_5568),
.Y(n_6425)
);

BUFx2_ASAP7_75t_L g6426 ( 
.A(n_5755),
.Y(n_6426)
);

BUFx2_ASAP7_75t_L g6427 ( 
.A(n_5764),
.Y(n_6427)
);

BUFx2_ASAP7_75t_L g6428 ( 
.A(n_5764),
.Y(n_6428)
);

INVx3_ASAP7_75t_L g6429 ( 
.A(n_5772),
.Y(n_6429)
);

AOI22xp33_ASAP7_75t_SL g6430 ( 
.A1(n_5847),
.A2(n_5300),
.B1(n_5358),
.B2(n_5352),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_5842),
.Y(n_6431)
);

NAND3xp33_ASAP7_75t_L g6432 ( 
.A(n_5890),
.B(n_5568),
.C(n_5384),
.Y(n_6432)
);

AND2x2_ASAP7_75t_L g6433 ( 
.A(n_5928),
.B(n_5602),
.Y(n_6433)
);

AND2x2_ASAP7_75t_L g6434 ( 
.A(n_5941),
.B(n_5602),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_5974),
.Y(n_6435)
);

AND2x2_ASAP7_75t_L g6436 ( 
.A(n_5941),
.B(n_5603),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_5946),
.B(n_5603),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_6197),
.Y(n_6438)
);

OR2x2_ASAP7_75t_L g6439 ( 
.A(n_5751),
.B(n_5196),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6197),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_6197),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_L g6442 ( 
.A(n_5872),
.B(n_5154),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5843),
.Y(n_6443)
);

INVxp67_ASAP7_75t_SL g6444 ( 
.A(n_5811),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_5850),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_5851),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_5946),
.B(n_5651),
.Y(n_6447)
);

BUFx3_ASAP7_75t_L g6448 ( 
.A(n_6184),
.Y(n_6448)
);

AOI22xp33_ASAP7_75t_SL g6449 ( 
.A1(n_5865),
.A2(n_5300),
.B1(n_5358),
.B2(n_5352),
.Y(n_6449)
);

HB1xp67_ASAP7_75t_L g6450 ( 
.A(n_5875),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_5857),
.Y(n_6451)
);

INVx2_ASAP7_75t_L g6452 ( 
.A(n_6204),
.Y(n_6452)
);

BUFx4f_ASAP7_75t_L g6453 ( 
.A(n_5944),
.Y(n_6453)
);

AND2x2_ASAP7_75t_L g6454 ( 
.A(n_6039),
.B(n_5651),
.Y(n_6454)
);

BUFx2_ASAP7_75t_L g6455 ( 
.A(n_5859),
.Y(n_6455)
);

AND2x2_ASAP7_75t_L g6456 ( 
.A(n_5831),
.B(n_5154),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_5874),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_5876),
.Y(n_6458)
);

OR2x2_ASAP7_75t_L g6459 ( 
.A(n_5751),
.B(n_5196),
.Y(n_6459)
);

INVx2_ASAP7_75t_L g6460 ( 
.A(n_6204),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_6204),
.Y(n_6461)
);

NOR2xp33_ASAP7_75t_R g6462 ( 
.A(n_6181),
.B(n_5257),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5877),
.Y(n_6463)
);

NAND2xp5_ASAP7_75t_L g6464 ( 
.A(n_5934),
.B(n_5290),
.Y(n_6464)
);

INVx3_ASAP7_75t_L g6465 ( 
.A(n_5783),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_5937),
.B(n_5290),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_5882),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_5831),
.B(n_5259),
.Y(n_6468)
);

AND2x2_ASAP7_75t_L g6469 ( 
.A(n_5886),
.B(n_5259),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_5950),
.B(n_5290),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_5886),
.B(n_5259),
.Y(n_6471)
);

INVx2_ASAP7_75t_L g6472 ( 
.A(n_5968),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_5892),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_5893),
.Y(n_6474)
);

AND2x2_ASAP7_75t_L g6475 ( 
.A(n_5902),
.B(n_5259),
.Y(n_6475)
);

AND2x2_ASAP7_75t_L g6476 ( 
.A(n_5902),
.B(n_5188),
.Y(n_6476)
);

INVx2_ASAP7_75t_L g6477 ( 
.A(n_5968),
.Y(n_6477)
);

INVx2_ASAP7_75t_SL g6478 ( 
.A(n_5944),
.Y(n_6478)
);

AND2x2_ASAP7_75t_L g6479 ( 
.A(n_5963),
.B(n_5188),
.Y(n_6479)
);

OR2x2_ASAP7_75t_L g6480 ( 
.A(n_5767),
.B(n_5648),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_5894),
.Y(n_6481)
);

NAND2xp5_ASAP7_75t_L g6482 ( 
.A(n_5956),
.B(n_5962),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_5898),
.Y(n_6483)
);

AOI22xp33_ASAP7_75t_L g6484 ( 
.A1(n_5737),
.A2(n_5598),
.B1(n_5476),
.B2(n_5318),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_5899),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_5968),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_5901),
.Y(n_6487)
);

AND2x2_ASAP7_75t_L g6488 ( 
.A(n_5963),
.B(n_5230),
.Y(n_6488)
);

INVx2_ASAP7_75t_R g6489 ( 
.A(n_5957),
.Y(n_6489)
);

AND2x2_ASAP7_75t_L g6490 ( 
.A(n_5966),
.B(n_5997),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_5904),
.Y(n_6491)
);

HB1xp67_ASAP7_75t_L g6492 ( 
.A(n_6063),
.Y(n_6492)
);

BUFx2_ASAP7_75t_L g6493 ( 
.A(n_5859),
.Y(n_6493)
);

HB1xp67_ASAP7_75t_L g6494 ( 
.A(n_6106),
.Y(n_6494)
);

NOR2xp33_ASAP7_75t_L g6495 ( 
.A(n_6184),
.B(n_5428),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_5908),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_5966),
.B(n_5997),
.Y(n_6497)
);

INVx2_ASAP7_75t_L g6498 ( 
.A(n_5978),
.Y(n_6498)
);

INVx2_ASAP7_75t_L g6499 ( 
.A(n_5978),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_5978),
.Y(n_6500)
);

AND2x4_ASAP7_75t_L g6501 ( 
.A(n_6236),
.B(n_5290),
.Y(n_6501)
);

AND2x2_ASAP7_75t_L g6502 ( 
.A(n_6017),
.B(n_5230),
.Y(n_6502)
);

AOI33xp33_ASAP7_75t_L g6503 ( 
.A1(n_6185),
.A2(n_5698),
.A3(n_5198),
.B1(n_4865),
.B2(n_5228),
.B3(n_5237),
.Y(n_6503)
);

AND2x2_ASAP7_75t_L g6504 ( 
.A(n_6017),
.B(n_5251),
.Y(n_6504)
);

NAND2xp5_ASAP7_75t_L g6505 ( 
.A(n_6124),
.B(n_5290),
.Y(n_6505)
);

AND2x4_ASAP7_75t_L g6506 ( 
.A(n_6236),
.B(n_5332),
.Y(n_6506)
);

AND2x4_ASAP7_75t_L g6507 ( 
.A(n_6236),
.B(n_5332),
.Y(n_6507)
);

OA21x2_ASAP7_75t_L g6508 ( 
.A1(n_6060),
.A2(n_5491),
.B(n_5489),
.Y(n_6508)
);

INVx1_ASAP7_75t_L g6509 ( 
.A(n_5909),
.Y(n_6509)
);

BUFx6f_ASAP7_75t_L g6510 ( 
.A(n_6175),
.Y(n_6510)
);

NAND2xp5_ASAP7_75t_L g6511 ( 
.A(n_6139),
.B(n_6144),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_5811),
.Y(n_6512)
);

AND2x2_ASAP7_75t_L g6513 ( 
.A(n_6027),
.B(n_5251),
.Y(n_6513)
);

INVx2_ASAP7_75t_SL g6514 ( 
.A(n_5984),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_6238),
.B(n_5332),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_5838),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6027),
.B(n_5261),
.Y(n_6517)
);

OR2x2_ASAP7_75t_L g6518 ( 
.A(n_5767),
.B(n_5625),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_5913),
.Y(n_6519)
);

OR2x2_ASAP7_75t_L g6520 ( 
.A(n_5768),
.B(n_5625),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_5915),
.Y(n_6521)
);

INVx3_ASAP7_75t_SL g6522 ( 
.A(n_6181),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_5924),
.Y(n_6523)
);

INVx3_ASAP7_75t_L g6524 ( 
.A(n_5783),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_5931),
.Y(n_6525)
);

AND2x2_ASAP7_75t_L g6526 ( 
.A(n_5871),
.B(n_5261),
.Y(n_6526)
);

OR2x2_ASAP7_75t_L g6527 ( 
.A(n_5768),
.B(n_5660),
.Y(n_6527)
);

INVx3_ASAP7_75t_L g6528 ( 
.A(n_5783),
.Y(n_6528)
);

AND2x4_ASAP7_75t_L g6529 ( 
.A(n_6236),
.B(n_5332),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6135),
.B(n_5332),
.Y(n_6530)
);

INVx2_ASAP7_75t_L g6531 ( 
.A(n_5838),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_5933),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_5838),
.Y(n_6533)
);

AND2x2_ASAP7_75t_L g6534 ( 
.A(n_5871),
.B(n_5333),
.Y(n_6534)
);

OR2x2_ASAP7_75t_L g6535 ( 
.A(n_5903),
.B(n_5660),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_5940),
.Y(n_6536)
);

BUFx3_ASAP7_75t_L g6537 ( 
.A(n_5878),
.Y(n_6537)
);

OR2x2_ASAP7_75t_L g6538 ( 
.A(n_5903),
.B(n_5675),
.Y(n_6538)
);

AND2x4_ASAP7_75t_L g6539 ( 
.A(n_5818),
.B(n_5357),
.Y(n_6539)
);

BUFx2_ASAP7_75t_L g6540 ( 
.A(n_5957),
.Y(n_6540)
);

AND2x2_ASAP7_75t_L g6541 ( 
.A(n_6039),
.B(n_6218),
.Y(n_6541)
);

INVxp67_ASAP7_75t_SL g6542 ( 
.A(n_5860),
.Y(n_6542)
);

INVx2_ASAP7_75t_L g6543 ( 
.A(n_5879),
.Y(n_6543)
);

INVx3_ASAP7_75t_L g6544 ( 
.A(n_5795),
.Y(n_6544)
);

AO31x2_ASAP7_75t_L g6545 ( 
.A1(n_5860),
.A2(n_5745),
.A3(n_5756),
.B(n_5739),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6135),
.B(n_5357),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_5879),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_5879),
.Y(n_6548)
);

AND2x2_ASAP7_75t_L g6549 ( 
.A(n_6218),
.B(n_5871),
.Y(n_6549)
);

INVx2_ASAP7_75t_L g6550 ( 
.A(n_5889),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_5942),
.Y(n_6551)
);

BUFx2_ASAP7_75t_L g6552 ( 
.A(n_5995),
.Y(n_6552)
);

BUFx3_ASAP7_75t_L g6553 ( 
.A(n_5878),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_5945),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_5916),
.B(n_5663),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_5954),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_6163),
.B(n_5357),
.Y(n_6557)
);

INVx4_ASAP7_75t_L g6558 ( 
.A(n_5785),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_5889),
.Y(n_6559)
);

NAND2xp5_ASAP7_75t_L g6560 ( 
.A(n_6163),
.B(n_5357),
.Y(n_6560)
);

INVx1_ASAP7_75t_L g6561 ( 
.A(n_5958),
.Y(n_6561)
);

AND2x2_ASAP7_75t_L g6562 ( 
.A(n_5916),
.B(n_5922),
.Y(n_6562)
);

INVx2_ASAP7_75t_L g6563 ( 
.A(n_5889),
.Y(n_6563)
);

BUFx3_ASAP7_75t_L g6564 ( 
.A(n_5785),
.Y(n_6564)
);

INVxp67_ASAP7_75t_SL g6565 ( 
.A(n_5795),
.Y(n_6565)
);

INVx4_ASAP7_75t_SL g6566 ( 
.A(n_5984),
.Y(n_6566)
);

AND2x2_ASAP7_75t_L g6567 ( 
.A(n_5916),
.B(n_5333),
.Y(n_6567)
);

AND2x2_ASAP7_75t_L g6568 ( 
.A(n_5922),
.B(n_5407),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_5971),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_5973),
.Y(n_6570)
);

AOI21x1_ASAP7_75t_L g6571 ( 
.A1(n_5844),
.A2(n_5384),
.B(n_5271),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_5981),
.Y(n_6572)
);

AOI22xp33_ASAP7_75t_L g6573 ( 
.A1(n_5739),
.A2(n_5476),
.B1(n_5318),
.B2(n_5662),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_5922),
.B(n_5407),
.Y(n_6574)
);

INVx3_ASAP7_75t_L g6575 ( 
.A(n_5795),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6064),
.B(n_5411),
.Y(n_6576)
);

NOR2x1_ASAP7_75t_R g6577 ( 
.A(n_5742),
.B(n_5428),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_6064),
.B(n_5411),
.Y(n_6578)
);

INVxp67_ASAP7_75t_L g6579 ( 
.A(n_6016),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_5986),
.Y(n_6580)
);

NAND2xp5_ASAP7_75t_L g6581 ( 
.A(n_5880),
.B(n_5357),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_5989),
.Y(n_6582)
);

AND2x4_ASAP7_75t_L g6583 ( 
.A(n_6064),
.B(n_5796),
.Y(n_6583)
);

OA21x2_ASAP7_75t_L g6584 ( 
.A1(n_6051),
.A2(n_5499),
.B(n_5491),
.Y(n_6584)
);

INVx5_ASAP7_75t_L g6585 ( 
.A(n_5785),
.Y(n_6585)
);

BUFx6f_ASAP7_75t_L g6586 ( 
.A(n_5785),
.Y(n_6586)
);

NAND2xp5_ASAP7_75t_L g6587 ( 
.A(n_6172),
.B(n_5533),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_5990),
.Y(n_6588)
);

OR2x2_ASAP7_75t_L g6589 ( 
.A(n_5797),
.B(n_5675),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_5993),
.Y(n_6590)
);

INVxp67_ASAP7_75t_SL g6591 ( 
.A(n_6233),
.Y(n_6591)
);

AND2x2_ASAP7_75t_L g6592 ( 
.A(n_6079),
.B(n_5533),
.Y(n_6592)
);

BUFx2_ASAP7_75t_L g6593 ( 
.A(n_5995),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6009),
.Y(n_6594)
);

AND2x2_ASAP7_75t_L g6595 ( 
.A(n_6079),
.B(n_5533),
.Y(n_6595)
);

AND2x2_ASAP7_75t_L g6596 ( 
.A(n_6164),
.B(n_5533),
.Y(n_6596)
);

INVx2_ASAP7_75t_L g6597 ( 
.A(n_6239),
.Y(n_6597)
);

INVx4_ASAP7_75t_L g6598 ( 
.A(n_5834),
.Y(n_6598)
);

AND2x2_ASAP7_75t_L g6599 ( 
.A(n_6164),
.B(n_5533),
.Y(n_6599)
);

NAND2xp5_ASAP7_75t_L g6600 ( 
.A(n_5798),
.B(n_5467),
.Y(n_6600)
);

NOR2xp67_ASAP7_75t_L g6601 ( 
.A(n_6065),
.B(n_5645),
.Y(n_6601)
);

BUFx3_ASAP7_75t_L g6602 ( 
.A(n_5834),
.Y(n_6602)
);

INVxp67_ASAP7_75t_L g6603 ( 
.A(n_5837),
.Y(n_6603)
);

BUFx2_ASAP7_75t_L g6604 ( 
.A(n_5984),
.Y(n_6604)
);

NAND3xp33_ASAP7_75t_L g6605 ( 
.A(n_5745),
.B(n_5440),
.C(n_5420),
.Y(n_6605)
);

NAND2xp5_ASAP7_75t_SL g6606 ( 
.A(n_6013),
.B(n_5595),
.Y(n_6606)
);

AND2x2_ASAP7_75t_L g6607 ( 
.A(n_5796),
.B(n_5693),
.Y(n_6607)
);

AOI221xp5_ASAP7_75t_L g6608 ( 
.A1(n_6179),
.A2(n_5300),
.B1(n_5379),
.B2(n_5358),
.C(n_5352),
.Y(n_6608)
);

INVx2_ASAP7_75t_L g6609 ( 
.A(n_6239),
.Y(n_6609)
);

INVx2_ASAP7_75t_L g6610 ( 
.A(n_6239),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_6011),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_5796),
.B(n_5693),
.Y(n_6612)
);

INVx3_ASAP7_75t_L g6613 ( 
.A(n_5743),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6014),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_5960),
.Y(n_6615)
);

BUFx2_ASAP7_75t_L g6616 ( 
.A(n_5984),
.Y(n_6616)
);

NOR2xp67_ASAP7_75t_L g6617 ( 
.A(n_6065),
.B(n_5582),
.Y(n_6617)
);

OAI22xp5_ASAP7_75t_SL g6618 ( 
.A1(n_5983),
.A2(n_5438),
.B1(n_5517),
.B2(n_5116),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_5823),
.B(n_5663),
.Y(n_6619)
);

OAI21xp5_ASAP7_75t_SL g6620 ( 
.A1(n_6146),
.A2(n_5347),
.B(n_5463),
.Y(n_6620)
);

HB1xp67_ASAP7_75t_L g6621 ( 
.A(n_6024),
.Y(n_6621)
);

NOR2x1p5_ASAP7_75t_L g6622 ( 
.A(n_5834),
.B(n_5257),
.Y(n_6622)
);

AO21x2_ASAP7_75t_L g6623 ( 
.A1(n_5756),
.A2(n_5445),
.B(n_5442),
.Y(n_6623)
);

HB1xp67_ASAP7_75t_L g6624 ( 
.A(n_6025),
.Y(n_6624)
);

BUFx2_ASAP7_75t_L g6625 ( 
.A(n_5834),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_6026),
.Y(n_6626)
);

HB1xp67_ASAP7_75t_L g6627 ( 
.A(n_6032),
.Y(n_6627)
);

INVx2_ASAP7_75t_L g6628 ( 
.A(n_5960),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6033),
.Y(n_6629)
);

INVx2_ASAP7_75t_L g6630 ( 
.A(n_5967),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_5917),
.B(n_5218),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_5967),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6038),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_5823),
.B(n_5708),
.Y(n_6634)
);

INVx2_ASAP7_75t_L g6635 ( 
.A(n_5972),
.Y(n_6635)
);

AND2x4_ASAP7_75t_L g6636 ( 
.A(n_5823),
.B(n_5420),
.Y(n_6636)
);

INVx2_ASAP7_75t_L g6637 ( 
.A(n_5972),
.Y(n_6637)
);

NOR2xp33_ASAP7_75t_L g6638 ( 
.A(n_6211),
.B(n_5607),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6040),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6041),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_5830),
.B(n_5708),
.Y(n_6641)
);

HB1xp67_ASAP7_75t_L g6642 ( 
.A(n_6042),
.Y(n_6642)
);

AND2x2_ASAP7_75t_L g6643 ( 
.A(n_5830),
.B(n_5607),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_5976),
.Y(n_6644)
);

INVx2_ASAP7_75t_L g6645 ( 
.A(n_5976),
.Y(n_6645)
);

AND2x2_ASAP7_75t_L g6646 ( 
.A(n_5830),
.B(n_5731),
.Y(n_6646)
);

HB1xp67_ASAP7_75t_L g6647 ( 
.A(n_6053),
.Y(n_6647)
);

BUFx3_ASAP7_75t_L g6648 ( 
.A(n_5873),
.Y(n_6648)
);

INVx2_ASAP7_75t_L g6649 ( 
.A(n_5965),
.Y(n_6649)
);

INVx3_ASAP7_75t_L g6650 ( 
.A(n_5743),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_5965),
.Y(n_6651)
);

AND2x2_ASAP7_75t_L g6652 ( 
.A(n_5987),
.B(n_6035),
.Y(n_6652)
);

AND2x2_ASAP7_75t_L g6653 ( 
.A(n_5987),
.B(n_5731),
.Y(n_6653)
);

INVx2_ASAP7_75t_SL g6654 ( 
.A(n_5873),
.Y(n_6654)
);

INVx2_ASAP7_75t_L g6655 ( 
.A(n_5965),
.Y(n_6655)
);

INVx2_ASAP7_75t_L g6656 ( 
.A(n_5797),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_5917),
.B(n_5218),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6056),
.Y(n_6658)
);

NAND3xp33_ASAP7_75t_L g6659 ( 
.A(n_5762),
.B(n_5440),
.C(n_5662),
.Y(n_6659)
);

INVx2_ASAP7_75t_L g6660 ( 
.A(n_5801),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_5987),
.B(n_5049),
.Y(n_6661)
);

HB1xp67_ASAP7_75t_L g6662 ( 
.A(n_6057),
.Y(n_6662)
);

HB1xp67_ASAP7_75t_L g6663 ( 
.A(n_6061),
.Y(n_6663)
);

HB1xp67_ASAP7_75t_L g6664 ( 
.A(n_6062),
.Y(n_6664)
);

NAND2xp5_ASAP7_75t_L g6665 ( 
.A(n_5824),
.B(n_5897),
.Y(n_6665)
);

OR2x2_ASAP7_75t_L g6666 ( 
.A(n_5801),
.B(n_5718),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6067),
.Y(n_6667)
);

AND2x2_ASAP7_75t_L g6668 ( 
.A(n_6035),
.B(n_5239),
.Y(n_6668)
);

BUFx6f_ASAP7_75t_L g6669 ( 
.A(n_5873),
.Y(n_6669)
);

OR2x2_ASAP7_75t_L g6670 ( 
.A(n_5824),
.B(n_5718),
.Y(n_6670)
);

AND2x2_ASAP7_75t_L g6671 ( 
.A(n_5867),
.B(n_5616),
.Y(n_6671)
);

AND2x2_ASAP7_75t_L g6672 ( 
.A(n_5793),
.B(n_5616),
.Y(n_6672)
);

INVx3_ASAP7_75t_L g6673 ( 
.A(n_5873),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6071),
.Y(n_6674)
);

OAI211xp5_ASAP7_75t_SL g6675 ( 
.A1(n_5883),
.A2(n_5900),
.B(n_6165),
.C(n_6013),
.Y(n_6675)
);

BUFx8_ASAP7_75t_L g6676 ( 
.A(n_6095),
.Y(n_6676)
);

HB1xp67_ASAP7_75t_L g6677 ( 
.A(n_6072),
.Y(n_6677)
);

HB1xp67_ASAP7_75t_L g6678 ( 
.A(n_6073),
.Y(n_6678)
);

AND2x2_ASAP7_75t_L g6679 ( 
.A(n_5793),
.B(n_5616),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6003),
.B(n_5721),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6003),
.B(n_5721),
.Y(n_6681)
);

AND2x2_ASAP7_75t_L g6682 ( 
.A(n_6069),
.B(n_5721),
.Y(n_6682)
);

INVx2_ASAP7_75t_L g6683 ( 
.A(n_6005),
.Y(n_6683)
);

HB1xp67_ASAP7_75t_L g6684 ( 
.A(n_6075),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_6078),
.Y(n_6685)
);

INVx2_ASAP7_75t_L g6686 ( 
.A(n_6005),
.Y(n_6686)
);

OR2x2_ASAP7_75t_L g6687 ( 
.A(n_5897),
.B(n_5720),
.Y(n_6687)
);

OR2x2_ASAP7_75t_L g6688 ( 
.A(n_5948),
.B(n_5750),
.Y(n_6688)
);

BUFx2_ASAP7_75t_L g6689 ( 
.A(n_5742),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6080),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6085),
.Y(n_6691)
);

AND2x2_ASAP7_75t_L g6692 ( 
.A(n_6069),
.B(n_5721),
.Y(n_6692)
);

INVx1_ASAP7_75t_SL g6693 ( 
.A(n_6094),
.Y(n_6693)
);

INVxp67_ASAP7_75t_L g6694 ( 
.A(n_6037),
.Y(n_6694)
);

INVx2_ASAP7_75t_L g6695 ( 
.A(n_6005),
.Y(n_6695)
);

INVx2_ASAP7_75t_L g6696 ( 
.A(n_6006),
.Y(n_6696)
);

AND2x4_ASAP7_75t_L g6697 ( 
.A(n_6035),
.B(n_5679),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6088),
.Y(n_6698)
);

AND2x2_ASAP7_75t_L g6699 ( 
.A(n_6074),
.B(n_5721),
.Y(n_6699)
);

HB1xp67_ASAP7_75t_L g6700 ( 
.A(n_6288),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6281),
.Y(n_6701)
);

OAI22xp5_ASAP7_75t_L g6702 ( 
.A1(n_6338),
.A2(n_6242),
.B1(n_5900),
.B2(n_5862),
.Y(n_6702)
);

INVx3_ASAP7_75t_L g6703 ( 
.A(n_6335),
.Y(n_6703)
);

AND2x2_ASAP7_75t_L g6704 ( 
.A(n_6289),
.B(n_5822),
.Y(n_6704)
);

AND2x2_ASAP7_75t_L g6705 ( 
.A(n_6541),
.B(n_5822),
.Y(n_6705)
);

AND2x2_ASAP7_75t_L g6706 ( 
.A(n_6541),
.B(n_5848),
.Y(n_6706)
);

INVx2_ASAP7_75t_SL g6707 ( 
.A(n_6262),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_6280),
.Y(n_6708)
);

AND2x2_ASAP7_75t_L g6709 ( 
.A(n_6282),
.B(n_5848),
.Y(n_6709)
);

BUFx2_ASAP7_75t_L g6710 ( 
.A(n_6280),
.Y(n_6710)
);

AND2x4_ASAP7_75t_L g6711 ( 
.A(n_6643),
.B(n_5885),
.Y(n_6711)
);

AND2x2_ASAP7_75t_L g6712 ( 
.A(n_6355),
.B(n_5885),
.Y(n_6712)
);

AND2x2_ASAP7_75t_L g6713 ( 
.A(n_6276),
.B(n_5975),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6621),
.Y(n_6714)
);

OR2x2_ASAP7_75t_L g6715 ( 
.A(n_6303),
.B(n_5948),
.Y(n_6715)
);

INVx2_ASAP7_75t_SL g6716 ( 
.A(n_6262),
.Y(n_6716)
);

INVxp67_ASAP7_75t_SL g6717 ( 
.A(n_6288),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6396),
.Y(n_6718)
);

NAND2xp5_ASAP7_75t_L g6719 ( 
.A(n_6326),
.B(n_6090),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6621),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6624),
.Y(n_6721)
);

AND2x2_ASAP7_75t_L g6722 ( 
.A(n_6279),
.B(n_5975),
.Y(n_6722)
);

AND2x2_ASAP7_75t_L g6723 ( 
.A(n_6549),
.B(n_6004),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6624),
.Y(n_6724)
);

NAND2xp5_ASAP7_75t_L g6725 ( 
.A(n_6326),
.B(n_6093),
.Y(n_6725)
);

INVxp67_ASAP7_75t_L g6726 ( 
.A(n_6335),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6627),
.Y(n_6727)
);

BUFx6f_ASAP7_75t_L g6728 ( 
.A(n_6373),
.Y(n_6728)
);

OR2x2_ASAP7_75t_L g6729 ( 
.A(n_6318),
.B(n_5919),
.Y(n_6729)
);

BUFx6f_ASAP7_75t_L g6730 ( 
.A(n_6373),
.Y(n_6730)
);

BUFx3_ASAP7_75t_L g6731 ( 
.A(n_6448),
.Y(n_6731)
);

INVx2_ASAP7_75t_L g6732 ( 
.A(n_6268),
.Y(n_6732)
);

AND2x2_ASAP7_75t_L g6733 ( 
.A(n_6549),
.B(n_6004),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6627),
.Y(n_6734)
);

AND2x2_ASAP7_75t_L g6735 ( 
.A(n_6402),
.B(n_5742),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6299),
.B(n_6095),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6642),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6642),
.Y(n_6738)
);

AND2x2_ASAP7_75t_L g6739 ( 
.A(n_6378),
.B(n_6379),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6396),
.Y(n_6740)
);

AND2x2_ASAP7_75t_L g6741 ( 
.A(n_6381),
.B(n_6095),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6384),
.B(n_6095),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_6656),
.B(n_6096),
.Y(n_6743)
);

INVxp67_ASAP7_75t_L g6744 ( 
.A(n_6426),
.Y(n_6744)
);

BUFx3_ASAP7_75t_L g6745 ( 
.A(n_6448),
.Y(n_6745)
);

AND2x2_ASAP7_75t_L g6746 ( 
.A(n_6407),
.B(n_6054),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6652),
.B(n_6054),
.Y(n_6747)
);

AND2x2_ASAP7_75t_L g6748 ( 
.A(n_6284),
.B(n_6054),
.Y(n_6748)
);

OR2x6_ASAP7_75t_L g6749 ( 
.A(n_6336),
.B(n_6054),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6656),
.B(n_6097),
.Y(n_6750)
);

NOR2xp33_ASAP7_75t_L g6751 ( 
.A(n_6360),
.B(n_6054),
.Y(n_6751)
);

HB1xp67_ASAP7_75t_L g6752 ( 
.A(n_6272),
.Y(n_6752)
);

AND2x4_ASAP7_75t_L g6753 ( 
.A(n_6490),
.B(n_6128),
.Y(n_6753)
);

BUFx2_ASAP7_75t_SL g6754 ( 
.A(n_6287),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_SL g6755 ( 
.A(n_6263),
.B(n_6693),
.Y(n_6755)
);

AND2x2_ASAP7_75t_L g6756 ( 
.A(n_6285),
.B(n_6222),
.Y(n_6756)
);

NOR2xp33_ASAP7_75t_L g6757 ( 
.A(n_6360),
.B(n_6270),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6660),
.B(n_6100),
.Y(n_6758)
);

BUFx2_ASAP7_75t_L g6759 ( 
.A(n_6676),
.Y(n_6759)
);

BUFx3_ASAP7_75t_L g6760 ( 
.A(n_6287),
.Y(n_6760)
);

BUFx2_ASAP7_75t_SL g6761 ( 
.A(n_6306),
.Y(n_6761)
);

HB1xp67_ASAP7_75t_L g6762 ( 
.A(n_6272),
.Y(n_6762)
);

OR2x6_ASAP7_75t_L g6763 ( 
.A(n_6336),
.B(n_5301),
.Y(n_6763)
);

AND2x4_ASAP7_75t_L g6764 ( 
.A(n_6497),
.B(n_6128),
.Y(n_6764)
);

OR2x2_ASAP7_75t_L g6765 ( 
.A(n_6354),
.B(n_5919),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_6586),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6660),
.B(n_6101),
.Y(n_6767)
);

AND2x4_ASAP7_75t_L g6768 ( 
.A(n_6375),
.B(n_6128),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6295),
.B(n_6156),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6296),
.B(n_6156),
.Y(n_6770)
);

INVx2_ASAP7_75t_L g6771 ( 
.A(n_6586),
.Y(n_6771)
);

NAND2xp5_ASAP7_75t_L g6772 ( 
.A(n_6315),
.B(n_6103),
.Y(n_6772)
);

BUFx2_ASAP7_75t_L g6773 ( 
.A(n_6676),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_L g6774 ( 
.A(n_6315),
.B(n_6104),
.Y(n_6774)
);

HB1xp67_ASAP7_75t_L g6775 ( 
.A(n_6290),
.Y(n_6775)
);

HB1xp67_ASAP7_75t_L g6776 ( 
.A(n_6290),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6647),
.Y(n_6777)
);

NAND2xp5_ASAP7_75t_L g6778 ( 
.A(n_6372),
.B(n_6112),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6647),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6298),
.B(n_6156),
.Y(n_6780)
);

NAND2xp5_ASAP7_75t_L g6781 ( 
.A(n_6372),
.B(n_6113),
.Y(n_6781)
);

AND2x2_ASAP7_75t_L g6782 ( 
.A(n_6427),
.B(n_6214),
.Y(n_6782)
);

OR2x2_ASAP7_75t_L g6783 ( 
.A(n_6665),
.B(n_5750),
.Y(n_6783)
);

AND2x2_ASAP7_75t_L g6784 ( 
.A(n_6428),
.B(n_6214),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6662),
.Y(n_6785)
);

OR2x2_ASAP7_75t_L g6786 ( 
.A(n_6688),
.B(n_5929),
.Y(n_6786)
);

AND2x2_ASAP7_75t_L g6787 ( 
.A(n_6646),
.B(n_6074),
.Y(n_6787)
);

AND2x2_ASAP7_75t_L g6788 ( 
.A(n_6653),
.B(n_6082),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6662),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6663),
.Y(n_6790)
);

AND2x2_ASAP7_75t_L g6791 ( 
.A(n_6454),
.B(n_6082),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6454),
.B(n_6583),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6663),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6664),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6664),
.Y(n_6795)
);

AND2x2_ASAP7_75t_L g6796 ( 
.A(n_6583),
.B(n_6083),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_L g6797 ( 
.A(n_6374),
.B(n_6118),
.Y(n_6797)
);

AND2x2_ASAP7_75t_L g6798 ( 
.A(n_6583),
.B(n_6433),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6677),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6433),
.B(n_6083),
.Y(n_6800)
);

AND2x2_ASAP7_75t_L g6801 ( 
.A(n_6434),
.B(n_6086),
.Y(n_6801)
);

INVx2_ASAP7_75t_L g6802 ( 
.A(n_6268),
.Y(n_6802)
);

INVx3_ASAP7_75t_L g6803 ( 
.A(n_6306),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6305),
.Y(n_6804)
);

INVx2_ASAP7_75t_L g6805 ( 
.A(n_6305),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6677),
.Y(n_6806)
);

INVx1_ASAP7_75t_L g6807 ( 
.A(n_6678),
.Y(n_6807)
);

AND2x2_ASAP7_75t_L g6808 ( 
.A(n_6434),
.B(n_6086),
.Y(n_6808)
);

OR2x2_ASAP7_75t_L g6809 ( 
.A(n_6358),
.B(n_5929),
.Y(n_6809)
);

AND2x2_ASAP7_75t_L g6810 ( 
.A(n_6436),
.B(n_6121),
.Y(n_6810)
);

AND2x2_ASAP7_75t_L g6811 ( 
.A(n_6436),
.B(n_6121),
.Y(n_6811)
);

OR2x2_ASAP7_75t_L g6812 ( 
.A(n_6480),
.B(n_5939),
.Y(n_6812)
);

AND2x2_ASAP7_75t_L g6813 ( 
.A(n_6437),
.B(n_6145),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6678),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6586),
.Y(n_6815)
);

AND2x2_ASAP7_75t_SL g6816 ( 
.A(n_6292),
.B(n_6046),
.Y(n_6816)
);

AND2x4_ASAP7_75t_L g6817 ( 
.A(n_6300),
.B(n_5844),
.Y(n_6817)
);

OR2x2_ASAP7_75t_L g6818 ( 
.A(n_6297),
.B(n_5939),
.Y(n_6818)
);

AND2x2_ASAP7_75t_L g6819 ( 
.A(n_6437),
.B(n_6145),
.Y(n_6819)
);

OR2x2_ASAP7_75t_L g6820 ( 
.A(n_6482),
.B(n_6511),
.Y(n_6820)
);

AND2x4_ASAP7_75t_SL g6821 ( 
.A(n_6319),
.B(n_6337),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_L g6822 ( 
.A(n_6374),
.B(n_6119),
.Y(n_6822)
);

INVxp67_ASAP7_75t_L g6823 ( 
.A(n_6638),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6684),
.Y(n_6824)
);

AND2x2_ASAP7_75t_L g6825 ( 
.A(n_6447),
.B(n_6243),
.Y(n_6825)
);

HB1xp67_ASAP7_75t_L g6826 ( 
.A(n_6322),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6586),
.Y(n_6827)
);

INVx1_ASAP7_75t_SL g6828 ( 
.A(n_6522),
.Y(n_6828)
);

OR2x2_ASAP7_75t_L g6829 ( 
.A(n_6267),
.B(n_5998),
.Y(n_6829)
);

AND2x4_ASAP7_75t_L g6830 ( 
.A(n_6300),
.B(n_6089),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6684),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6393),
.Y(n_6832)
);

INVxp67_ASAP7_75t_L g6833 ( 
.A(n_6638),
.Y(n_6833)
);

HB1xp67_ASAP7_75t_L g6834 ( 
.A(n_6322),
.Y(n_6834)
);

INVx2_ASAP7_75t_L g6835 ( 
.A(n_6669),
.Y(n_6835)
);

AND2x2_ASAP7_75t_L g6836 ( 
.A(n_6447),
.B(n_6199),
.Y(n_6836)
);

OR2x2_ASAP7_75t_L g6837 ( 
.A(n_6304),
.B(n_5998),
.Y(n_6837)
);

INVxp67_ASAP7_75t_SL g6838 ( 
.A(n_6565),
.Y(n_6838)
);

AND2x4_ASAP7_75t_L g6839 ( 
.A(n_6260),
.B(n_6089),
.Y(n_6839)
);

NOR2x1_ASAP7_75t_L g6840 ( 
.A(n_6558),
.B(n_6598),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6596),
.B(n_6199),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6599),
.B(n_6310),
.Y(n_6842)
);

BUFx2_ASAP7_75t_L g6843 ( 
.A(n_6676),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6393),
.Y(n_6844)
);

AND2x2_ASAP7_75t_L g6845 ( 
.A(n_6495),
.B(n_6200),
.Y(n_6845)
);

INVx1_ASAP7_75t_SL g6846 ( 
.A(n_6522),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6395),
.Y(n_6847)
);

NAND2xp5_ASAP7_75t_L g6848 ( 
.A(n_6395),
.B(n_6122),
.Y(n_6848)
);

AND2x2_ASAP7_75t_L g6849 ( 
.A(n_6495),
.B(n_6200),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6450),
.B(n_6123),
.Y(n_6850)
);

OR2x2_ASAP7_75t_L g6851 ( 
.A(n_6631),
.B(n_6008),
.Y(n_6851)
);

OR2x2_ASAP7_75t_L g6852 ( 
.A(n_6657),
.B(n_6261),
.Y(n_6852)
);

INVxp67_ASAP7_75t_SL g6853 ( 
.A(n_6565),
.Y(n_6853)
);

INVx4_ASAP7_75t_L g6854 ( 
.A(n_6360),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6312),
.B(n_5970),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6450),
.Y(n_6856)
);

INVx3_ASAP7_75t_L g6857 ( 
.A(n_6697),
.Y(n_6857)
);

INVxp67_ASAP7_75t_L g6858 ( 
.A(n_6540),
.Y(n_6858)
);

INVx1_ASAP7_75t_L g6859 ( 
.A(n_6492),
.Y(n_6859)
);

OR2x2_ASAP7_75t_L g6860 ( 
.A(n_6492),
.B(n_6008),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_6494),
.B(n_6126),
.Y(n_6861)
);

HB1xp67_ASAP7_75t_L g6862 ( 
.A(n_6494),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6293),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_6669),
.Y(n_6864)
);

OR2x2_ASAP7_75t_L g6865 ( 
.A(n_6518),
.B(n_6018),
.Y(n_6865)
);

AND2x2_ASAP7_75t_L g6866 ( 
.A(n_6314),
.B(n_5970),
.Y(n_6866)
);

AND2x4_ASAP7_75t_L g6867 ( 
.A(n_6260),
.B(n_6294),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_6266),
.B(n_6130),
.Y(n_6868)
);

AOI22xp33_ASAP7_75t_L g6869 ( 
.A1(n_6342),
.A2(n_5762),
.B1(n_6231),
.B2(n_5799),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6301),
.Y(n_6870)
);

INVx1_ASAP7_75t_SL g6871 ( 
.A(n_6462),
.Y(n_6871)
);

INVx2_ASAP7_75t_L g6872 ( 
.A(n_6669),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6308),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6309),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6321),
.B(n_5970),
.Y(n_6875)
);

AND2x4_ASAP7_75t_L g6876 ( 
.A(n_6260),
.B(n_6089),
.Y(n_6876)
);

INVx1_ASAP7_75t_L g6877 ( 
.A(n_6313),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6316),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6317),
.Y(n_6879)
);

INVx3_ASAP7_75t_L g6880 ( 
.A(n_6697),
.Y(n_6880)
);

AND2x2_ASAP7_75t_L g6881 ( 
.A(n_6328),
.B(n_5970),
.Y(n_6881)
);

AND2x4_ASAP7_75t_L g6882 ( 
.A(n_6294),
.B(n_6110),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6324),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_6325),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6329),
.B(n_5996),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6333),
.B(n_5996),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6332),
.Y(n_6887)
);

AND2x2_ASAP7_75t_L g6888 ( 
.A(n_6264),
.B(n_5996),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_6669),
.Y(n_6889)
);

INVx2_ASAP7_75t_L g6890 ( 
.A(n_6564),
.Y(n_6890)
);

NOR2xp33_ASAP7_75t_L g6891 ( 
.A(n_6368),
.B(n_6022),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6564),
.Y(n_6892)
);

INVx4_ASAP7_75t_L g6893 ( 
.A(n_6286),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6341),
.Y(n_6894)
);

BUFx3_ASAP7_75t_L g6895 ( 
.A(n_6286),
.Y(n_6895)
);

AND2x4_ASAP7_75t_L g6896 ( 
.A(n_6294),
.B(n_6110),
.Y(n_6896)
);

INVx2_ASAP7_75t_L g6897 ( 
.A(n_6273),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6343),
.Y(n_6898)
);

AND2x4_ASAP7_75t_L g6899 ( 
.A(n_6311),
.B(n_6110),
.Y(n_6899)
);

AND2x2_ASAP7_75t_L g6900 ( 
.A(n_6264),
.B(n_6265),
.Y(n_6900)
);

BUFx2_ASAP7_75t_L g6901 ( 
.A(n_6462),
.Y(n_6901)
);

NAND2xp5_ASAP7_75t_L g6902 ( 
.A(n_6591),
.B(n_6131),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6346),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_6591),
.B(n_6143),
.Y(n_6904)
);

NAND2x1_ASAP7_75t_L g6905 ( 
.A(n_6311),
.B(n_6138),
.Y(n_6905)
);

AND2x2_ASAP7_75t_L g6906 ( 
.A(n_6265),
.B(n_5996),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6273),
.Y(n_6907)
);

AND2x2_ASAP7_75t_L g6908 ( 
.A(n_6271),
.B(n_6010),
.Y(n_6908)
);

INVx2_ASAP7_75t_L g6909 ( 
.A(n_6277),
.Y(n_6909)
);

AND2x2_ASAP7_75t_L g6910 ( 
.A(n_6271),
.B(n_6010),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6348),
.Y(n_6911)
);

AND2x4_ASAP7_75t_L g6912 ( 
.A(n_6311),
.B(n_6138),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6352),
.Y(n_6913)
);

AND2x2_ASAP7_75t_L g6914 ( 
.A(n_6340),
.B(n_6010),
.Y(n_6914)
);

AND2x2_ASAP7_75t_L g6915 ( 
.A(n_6340),
.B(n_6010),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6361),
.Y(n_6916)
);

NAND2x1p5_ASAP7_75t_SL g6917 ( 
.A(n_6654),
.B(n_6132),
.Y(n_6917)
);

INVx2_ASAP7_75t_SL g6918 ( 
.A(n_6622),
.Y(n_6918)
);

AND2x4_ASAP7_75t_L g6919 ( 
.A(n_6319),
.B(n_6138),
.Y(n_6919)
);

OR2x2_ASAP7_75t_L g6920 ( 
.A(n_6520),
.B(n_6018),
.Y(n_6920)
);

OR2x2_ASAP7_75t_L g6921 ( 
.A(n_6527),
.B(n_6043),
.Y(n_6921)
);

INVxp67_ASAP7_75t_SL g6922 ( 
.A(n_6403),
.Y(n_6922)
);

NAND2xp5_ASAP7_75t_L g6923 ( 
.A(n_6364),
.B(n_6148),
.Y(n_6923)
);

NAND2xp5_ASAP7_75t_L g6924 ( 
.A(n_6365),
.B(n_6155),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6602),
.Y(n_6925)
);

INVx2_ASAP7_75t_L g6926 ( 
.A(n_6602),
.Y(n_6926)
);

INVx2_ASAP7_75t_L g6927 ( 
.A(n_6648),
.Y(n_6927)
);

INVx2_ASAP7_75t_L g6928 ( 
.A(n_6648),
.Y(n_6928)
);

OAI21xp5_ASAP7_75t_L g6929 ( 
.A1(n_6606),
.A2(n_5853),
.B(n_5926),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6345),
.B(n_6066),
.Y(n_6930)
);

AND2x4_ASAP7_75t_SL g6931 ( 
.A(n_6319),
.B(n_4926),
.Y(n_6931)
);

NAND2xp5_ASAP7_75t_L g6932 ( 
.A(n_6376),
.B(n_6166),
.Y(n_6932)
);

NAND2xp5_ASAP7_75t_L g6933 ( 
.A(n_6383),
.B(n_6167),
.Y(n_6933)
);

OR2x6_ASAP7_75t_L g6934 ( 
.A(n_6336),
.B(n_5301),
.Y(n_6934)
);

INVx1_ASAP7_75t_L g6935 ( 
.A(n_6387),
.Y(n_6935)
);

INVxp67_ASAP7_75t_L g6936 ( 
.A(n_6552),
.Y(n_6936)
);

AND2x2_ASAP7_75t_L g6937 ( 
.A(n_6345),
.B(n_6066),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6388),
.Y(n_6938)
);

AND2x2_ASAP7_75t_L g6939 ( 
.A(n_6347),
.B(n_6066),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_6347),
.B(n_6066),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6390),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_6394),
.B(n_6168),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6400),
.Y(n_6943)
);

INVx2_ASAP7_75t_L g6944 ( 
.A(n_6673),
.Y(n_6944)
);

INVx4_ASAP7_75t_L g6945 ( 
.A(n_6286),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6408),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_6409),
.B(n_6194),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6416),
.Y(n_6948)
);

NAND2xp5_ASAP7_75t_L g6949 ( 
.A(n_6431),
.B(n_6169),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6443),
.Y(n_6950)
);

AOI22xp33_ASAP7_75t_L g6951 ( 
.A1(n_6342),
.A2(n_5799),
.B1(n_5887),
.B2(n_5969),
.Y(n_6951)
);

AND2x4_ASAP7_75t_L g6952 ( 
.A(n_6337),
.B(n_6225),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_6409),
.B(n_6194),
.Y(n_6953)
);

AND2x2_ASAP7_75t_L g6954 ( 
.A(n_6414),
.B(n_6194),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6673),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6445),
.Y(n_6956)
);

BUFx2_ASAP7_75t_L g6957 ( 
.A(n_6337),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_6446),
.Y(n_6958)
);

HB1xp67_ASAP7_75t_L g6959 ( 
.A(n_6327),
.Y(n_6959)
);

AND2x2_ASAP7_75t_SL g6960 ( 
.A(n_6292),
.B(n_6046),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6451),
.Y(n_6961)
);

AND2x2_ASAP7_75t_L g6962 ( 
.A(n_6414),
.B(n_6194),
.Y(n_6962)
);

AND2x2_ASAP7_75t_L g6963 ( 
.A(n_6415),
.B(n_6422),
.Y(n_6963)
);

INVx3_ASAP7_75t_L g6964 ( 
.A(n_6697),
.Y(n_6964)
);

AND2x2_ASAP7_75t_L g6965 ( 
.A(n_6415),
.B(n_6422),
.Y(n_6965)
);

AND2x2_ASAP7_75t_L g6966 ( 
.A(n_6425),
.B(n_6141),
.Y(n_6966)
);

OR2x2_ASAP7_75t_L g6967 ( 
.A(n_6666),
.B(n_6043),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6425),
.B(n_6141),
.Y(n_6968)
);

BUFx6f_ASAP7_75t_L g6969 ( 
.A(n_6286),
.Y(n_6969)
);

AND2x2_ASAP7_75t_L g6970 ( 
.A(n_6356),
.B(n_6257),
.Y(n_6970)
);

OR2x2_ASAP7_75t_L g6971 ( 
.A(n_6535),
.B(n_6052),
.Y(n_6971)
);

INVx2_ASAP7_75t_L g6972 ( 
.A(n_6673),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6457),
.Y(n_6973)
);

HB1xp67_ASAP7_75t_L g6974 ( 
.A(n_6327),
.Y(n_6974)
);

HB1xp67_ASAP7_75t_L g6975 ( 
.A(n_6334),
.Y(n_6975)
);

NAND2xp5_ASAP7_75t_L g6976 ( 
.A(n_6458),
.B(n_6463),
.Y(n_6976)
);

BUFx2_ASAP7_75t_L g6977 ( 
.A(n_6349),
.Y(n_6977)
);

AND2x2_ASAP7_75t_L g6978 ( 
.A(n_6357),
.B(n_6257),
.Y(n_6978)
);

AND2x4_ASAP7_75t_SL g6979 ( 
.A(n_6349),
.B(n_4926),
.Y(n_6979)
);

NAND2x1p5_ASAP7_75t_SL g6980 ( 
.A(n_6654),
.B(n_6132),
.Y(n_6980)
);

AND2x4_ASAP7_75t_L g6981 ( 
.A(n_6349),
.B(n_6225),
.Y(n_6981)
);

BUFx3_ASAP7_75t_L g6982 ( 
.A(n_6510),
.Y(n_6982)
);

INVxp67_ASAP7_75t_L g6983 ( 
.A(n_6593),
.Y(n_6983)
);

INVx3_ASAP7_75t_L g6984 ( 
.A(n_6501),
.Y(n_6984)
);

INVx2_ASAP7_75t_L g6985 ( 
.A(n_6672),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6467),
.Y(n_6986)
);

NOR2x1_ASAP7_75t_SL g6987 ( 
.A(n_6606),
.B(n_5887),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_6672),
.Y(n_6988)
);

OR2x2_ASAP7_75t_L g6989 ( 
.A(n_6538),
.B(n_6052),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6473),
.Y(n_6990)
);

AND2x2_ASAP7_75t_L g6991 ( 
.A(n_6363),
.B(n_6225),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_6474),
.B(n_6170),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6481),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_6483),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6485),
.Y(n_6995)
);

AND2x4_ASAP7_75t_L g6996 ( 
.A(n_6377),
.B(n_6226),
.Y(n_6996)
);

NAND2x1_ASAP7_75t_L g6997 ( 
.A(n_6601),
.B(n_6226),
.Y(n_6997)
);

INVx2_ASAP7_75t_L g6998 ( 
.A(n_6277),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6487),
.B(n_6173),
.Y(n_6999)
);

BUFx3_ASAP7_75t_L g7000 ( 
.A(n_6510),
.Y(n_7000)
);

INVx4_ASAP7_75t_L g7001 ( 
.A(n_6510),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6537),
.B(n_6226),
.Y(n_7002)
);

AND2x2_ASAP7_75t_L g7003 ( 
.A(n_6537),
.B(n_6255),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6278),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6491),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6553),
.B(n_6255),
.Y(n_7006)
);

BUFx2_ASAP7_75t_L g7007 ( 
.A(n_6377),
.Y(n_7007)
);

HB1xp67_ASAP7_75t_L g7008 ( 
.A(n_6334),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6496),
.Y(n_7009)
);

NOR2xp33_ASAP7_75t_L g7010 ( 
.A(n_6368),
.B(n_5123),
.Y(n_7010)
);

AND2x2_ASAP7_75t_L g7011 ( 
.A(n_6553),
.B(n_6255),
.Y(n_7011)
);

AND2x6_ASAP7_75t_L g7012 ( 
.A(n_6510),
.B(n_6423),
.Y(n_7012)
);

AND2x2_ASAP7_75t_L g7013 ( 
.A(n_6661),
.B(n_6455),
.Y(n_7013)
);

AND2x2_ASAP7_75t_L g7014 ( 
.A(n_6493),
.B(n_6162),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6679),
.Y(n_7015)
);

AND2x2_ASAP7_75t_L g7016 ( 
.A(n_6526),
.B(n_6162),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6509),
.B(n_6174),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6534),
.B(n_6196),
.Y(n_7018)
);

INVx2_ASAP7_75t_L g7019 ( 
.A(n_6679),
.Y(n_7019)
);

NAND2xp5_ASAP7_75t_L g7020 ( 
.A(n_6519),
.B(n_6178),
.Y(n_7020)
);

INVxp67_ASAP7_75t_L g7021 ( 
.A(n_6380),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6558),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6521),
.Y(n_7023)
);

INVx2_ASAP7_75t_L g7024 ( 
.A(n_6558),
.Y(n_7024)
);

AND2x2_ASAP7_75t_L g7025 ( 
.A(n_6567),
.B(n_6196),
.Y(n_7025)
);

AND2x4_ASAP7_75t_L g7026 ( 
.A(n_6377),
.B(n_6046),
.Y(n_7026)
);

AND2x2_ASAP7_75t_L g7027 ( 
.A(n_6568),
.B(n_6253),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6523),
.Y(n_7028)
);

NAND2xp5_ASAP7_75t_L g7029 ( 
.A(n_6525),
.B(n_6186),
.Y(n_7029)
);

INVx2_ASAP7_75t_L g7030 ( 
.A(n_6278),
.Y(n_7030)
);

AND2x2_ASAP7_75t_L g7031 ( 
.A(n_6574),
.B(n_6253),
.Y(n_7031)
);

INVx1_ASAP7_75t_L g7032 ( 
.A(n_6532),
.Y(n_7032)
);

NOR2xp33_ASAP7_75t_L g7033 ( 
.A(n_6413),
.B(n_6423),
.Y(n_7033)
);

BUFx2_ASAP7_75t_L g7034 ( 
.A(n_6401),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6536),
.Y(n_7035)
);

OR2x2_ASAP7_75t_L g7036 ( 
.A(n_6670),
.B(n_6687),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6350),
.Y(n_7037)
);

BUFx2_ASAP7_75t_L g7038 ( 
.A(n_6401),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6551),
.Y(n_7039)
);

INVx2_ASAP7_75t_L g7040 ( 
.A(n_6598),
.Y(n_7040)
);

AND2x2_ASAP7_75t_L g7041 ( 
.A(n_6576),
.B(n_6253),
.Y(n_7041)
);

INVxp67_ASAP7_75t_SL g7042 ( 
.A(n_6403),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6554),
.Y(n_7043)
);

AND2x2_ASAP7_75t_L g7044 ( 
.A(n_6578),
.B(n_4816),
.Y(n_7044)
);

AND2x2_ASAP7_75t_L g7045 ( 
.A(n_6668),
.B(n_4816),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_6366),
.B(n_4974),
.Y(n_7046)
);

OR2x2_ASAP7_75t_L g7047 ( 
.A(n_6589),
.B(n_6107),
.Y(n_7047)
);

AND2x2_ASAP7_75t_L g7048 ( 
.A(n_6371),
.B(n_6607),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6556),
.Y(n_7049)
);

BUFx3_ASAP7_75t_L g7050 ( 
.A(n_6380),
.Y(n_7050)
);

NOR2x1_ASAP7_75t_L g7051 ( 
.A(n_6598),
.B(n_6675),
.Y(n_7051)
);

AND2x2_ASAP7_75t_L g7052 ( 
.A(n_6612),
.B(n_4974),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6561),
.Y(n_7053)
);

INVx2_ASAP7_75t_L g7054 ( 
.A(n_6350),
.Y(n_7054)
);

OR2x2_ASAP7_75t_L g7055 ( 
.A(n_6600),
.B(n_6107),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_6592),
.B(n_4987),
.Y(n_7056)
);

HB1xp67_ASAP7_75t_L g7057 ( 
.A(n_6339),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6569),
.Y(n_7058)
);

INVxp33_ASAP7_75t_L g7059 ( 
.A(n_6577),
.Y(n_7059)
);

INVx2_ASAP7_75t_L g7060 ( 
.A(n_6302),
.Y(n_7060)
);

HB1xp67_ASAP7_75t_L g7061 ( 
.A(n_6339),
.Y(n_7061)
);

AND2x4_ASAP7_75t_L g7062 ( 
.A(n_6401),
.B(n_6127),
.Y(n_7062)
);

INVx6_ASAP7_75t_L g7063 ( 
.A(n_6585),
.Y(n_7063)
);

AND2x2_ASAP7_75t_L g7064 ( 
.A(n_6595),
.B(n_4987),
.Y(n_7064)
);

AND2x4_ASAP7_75t_L g7065 ( 
.A(n_6275),
.B(n_6127),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_6476),
.B(n_6127),
.Y(n_7066)
);

INVxp67_ASAP7_75t_SL g7067 ( 
.A(n_6444),
.Y(n_7067)
);

AND2x2_ASAP7_75t_L g7068 ( 
.A(n_6479),
.B(n_4688),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6302),
.Y(n_7069)
);

INVx2_ASAP7_75t_L g7070 ( 
.A(n_6302),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6488),
.B(n_4688),
.Y(n_7071)
);

AOI22xp33_ASAP7_75t_L g7072 ( 
.A1(n_6430),
.A2(n_5969),
.B1(n_6192),
.B2(n_5938),
.Y(n_7072)
);

HB1xp67_ASAP7_75t_L g7073 ( 
.A(n_6323),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6570),
.Y(n_7074)
);

NOR2xp33_ASAP7_75t_L g7075 ( 
.A(n_6694),
.B(n_5123),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_6572),
.B(n_6580),
.Y(n_7076)
);

AND2x2_ASAP7_75t_L g7077 ( 
.A(n_6502),
.B(n_4699),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6504),
.B(n_6513),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6582),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6588),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_6344),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6590),
.B(n_6189),
.Y(n_7082)
);

AND2x2_ASAP7_75t_L g7083 ( 
.A(n_6517),
.B(n_4699),
.Y(n_7083)
);

INVx2_ASAP7_75t_L g7084 ( 
.A(n_6344),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6594),
.Y(n_7085)
);

OAI22xp33_ASAP7_75t_L g7086 ( 
.A1(n_6620),
.A2(n_5476),
.B1(n_5683),
.B2(n_5352),
.Y(n_7086)
);

AND2x4_ASAP7_75t_L g7087 ( 
.A(n_6275),
.B(n_6165),
.Y(n_7087)
);

OR2x2_ASAP7_75t_L g7088 ( 
.A(n_6269),
.B(n_6154),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6611),
.Y(n_7089)
);

AO21x2_ASAP7_75t_L g7090 ( 
.A1(n_6542),
.A2(n_5938),
.B(n_5936),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_L g7091 ( 
.A(n_6614),
.B(n_6191),
.Y(n_7091)
);

INVx2_ASAP7_75t_L g7092 ( 
.A(n_6344),
.Y(n_7092)
);

NAND2xp5_ASAP7_75t_L g7093 ( 
.A(n_6626),
.B(n_6193),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6562),
.B(n_4699),
.Y(n_7094)
);

BUFx3_ASAP7_75t_L g7095 ( 
.A(n_6625),
.Y(n_7095)
);

INVx2_ASAP7_75t_L g7096 ( 
.A(n_6353),
.Y(n_7096)
);

BUFx2_ASAP7_75t_SL g7097 ( 
.A(n_6585),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6629),
.Y(n_7098)
);

AND2x2_ASAP7_75t_L g7099 ( 
.A(n_6619),
.B(n_4699),
.Y(n_7099)
);

AND2x2_ASAP7_75t_L g7100 ( 
.A(n_6634),
.B(n_5611),
.Y(n_7100)
);

BUFx3_ASAP7_75t_L g7101 ( 
.A(n_6585),
.Y(n_7101)
);

AND2x2_ASAP7_75t_L g7102 ( 
.A(n_6641),
.B(n_5611),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6633),
.Y(n_7103)
);

INVx2_ASAP7_75t_L g7104 ( 
.A(n_6429),
.Y(n_7104)
);

OR2x2_ASAP7_75t_L g7105 ( 
.A(n_6274),
.B(n_6154),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6639),
.Y(n_7106)
);

INVx3_ASAP7_75t_L g7107 ( 
.A(n_6501),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6640),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6658),
.Y(n_7109)
);

OR2x2_ASAP7_75t_L g7110 ( 
.A(n_6291),
.B(n_5881),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6667),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_6456),
.B(n_5638),
.Y(n_7112)
);

AND2x2_ASAP7_75t_L g7113 ( 
.A(n_6501),
.B(n_6506),
.Y(n_7113)
);

INVx2_ASAP7_75t_L g7114 ( 
.A(n_6429),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_L g7115 ( 
.A(n_6674),
.B(n_6198),
.Y(n_7115)
);

AND2x4_ASAP7_75t_L g7116 ( 
.A(n_6320),
.B(n_4926),
.Y(n_7116)
);

BUFx2_ASAP7_75t_L g7117 ( 
.A(n_6506),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6685),
.Y(n_7118)
);

NOR2xp33_ASAP7_75t_SL g7119 ( 
.A(n_6585),
.B(n_6453),
.Y(n_7119)
);

NOR2x1p5_ASAP7_75t_L g7120 ( 
.A(n_6557),
.B(n_5642),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6690),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6775),
.Y(n_7122)
);

OAI21xp5_ASAP7_75t_L g7123 ( 
.A1(n_6929),
.A2(n_6702),
.B(n_6951),
.Y(n_7123)
);

AOI21xp5_ASAP7_75t_L g7124 ( 
.A1(n_6987),
.A2(n_6449),
.B(n_6331),
.Y(n_7124)
);

NAND2xp5_ASAP7_75t_L g7125 ( 
.A(n_6755),
.B(n_6603),
.Y(n_7125)
);

INVx3_ASAP7_75t_L g7126 ( 
.A(n_6728),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6700),
.Y(n_7127)
);

AND2x2_ASAP7_75t_L g7128 ( 
.A(n_6754),
.B(n_6323),
.Y(n_7128)
);

AOI21xp5_ASAP7_75t_L g7129 ( 
.A1(n_6951),
.A2(n_6659),
.B(n_6351),
.Y(n_7129)
);

INVx4_ASAP7_75t_SL g7130 ( 
.A(n_7012),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6700),
.Y(n_7131)
);

INVx2_ASAP7_75t_L g7132 ( 
.A(n_6728),
.Y(n_7132)
);

NOR2xp67_ASAP7_75t_L g7133 ( 
.A(n_6703),
.B(n_6707),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6717),
.Y(n_7134)
);

OAI21xp5_ASAP7_75t_L g7135 ( 
.A1(n_6929),
.A2(n_6432),
.B(n_6584),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_6717),
.Y(n_7136)
);

OAI21xp5_ASAP7_75t_L g7137 ( 
.A1(n_6702),
.A2(n_6584),
.B(n_6420),
.Y(n_7137)
);

OAI21x1_ASAP7_75t_L g7138 ( 
.A1(n_6997),
.A2(n_6571),
.B(n_5853),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_6838),
.Y(n_7139)
);

AOI21xp5_ASAP7_75t_L g7140 ( 
.A1(n_7086),
.A2(n_6755),
.B(n_6869),
.Y(n_7140)
);

AOI21xp5_ASAP7_75t_L g7141 ( 
.A1(n_7086),
.A2(n_6508),
.B(n_6584),
.Y(n_7141)
);

OAI21xp33_ASAP7_75t_L g7142 ( 
.A1(n_7033),
.A2(n_6503),
.B(n_6560),
.Y(n_7142)
);

AOI21xp5_ASAP7_75t_L g7143 ( 
.A1(n_6869),
.A2(n_6508),
.B(n_6444),
.Y(n_7143)
);

OA21x2_ASAP7_75t_L g7144 ( 
.A1(n_6732),
.A2(n_6655),
.B(n_6649),
.Y(n_7144)
);

OAI21xp33_ASAP7_75t_L g7145 ( 
.A1(n_7033),
.A2(n_6503),
.B(n_6726),
.Y(n_7145)
);

INVx2_ASAP7_75t_L g7146 ( 
.A(n_6728),
.Y(n_7146)
);

OR2x2_ASAP7_75t_L g7147 ( 
.A(n_6786),
.B(n_6330),
.Y(n_7147)
);

BUFx3_ASAP7_75t_L g7148 ( 
.A(n_6730),
.Y(n_7148)
);

INVx3_ASAP7_75t_L g7149 ( 
.A(n_6730),
.Y(n_7149)
);

AND2x2_ASAP7_75t_L g7150 ( 
.A(n_6761),
.B(n_6330),
.Y(n_7150)
);

OA21x2_ASAP7_75t_L g7151 ( 
.A1(n_6732),
.A2(n_6651),
.B(n_6649),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_L g7152 ( 
.A(n_6726),
.B(n_6579),
.Y(n_7152)
);

OAI21xp5_ASAP7_75t_L g7153 ( 
.A1(n_7072),
.A2(n_7073),
.B(n_7051),
.Y(n_7153)
);

NOR2xp33_ASAP7_75t_R g7154 ( 
.A(n_6703),
.B(n_5393),
.Y(n_7154)
);

INVx2_ASAP7_75t_L g7155 ( 
.A(n_6730),
.Y(n_7155)
);

INVx2_ASAP7_75t_L g7156 ( 
.A(n_6760),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_6710),
.B(n_6307),
.Y(n_7157)
);

HB1xp67_ASAP7_75t_L g7158 ( 
.A(n_7073),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6858),
.B(n_6936),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6775),
.Y(n_7160)
);

INVx4_ASAP7_75t_L g7161 ( 
.A(n_6854),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6776),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_6858),
.B(n_6382),
.Y(n_7163)
);

INVx4_ASAP7_75t_L g7164 ( 
.A(n_6854),
.Y(n_7164)
);

AND2x4_ASAP7_75t_L g7165 ( 
.A(n_6760),
.B(n_6320),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_6776),
.Y(n_7166)
);

INVx2_ASAP7_75t_SL g7167 ( 
.A(n_6821),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6826),
.Y(n_7168)
);

NOR3xp33_ASAP7_75t_L g7169 ( 
.A(n_6871),
.B(n_6397),
.C(n_6542),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_6936),
.B(n_6404),
.Y(n_7170)
);

OA21x2_ASAP7_75t_L g7171 ( 
.A1(n_6802),
.A2(n_6651),
.B(n_6655),
.Y(n_7171)
);

OAI21xp33_ASAP7_75t_L g7172 ( 
.A1(n_7072),
.A2(n_6581),
.B(n_6546),
.Y(n_7172)
);

INVx2_ASAP7_75t_L g7173 ( 
.A(n_6731),
.Y(n_7173)
);

INVx2_ASAP7_75t_L g7174 ( 
.A(n_6731),
.Y(n_7174)
);

AND2x2_ASAP7_75t_L g7175 ( 
.A(n_6825),
.B(n_6468),
.Y(n_7175)
);

NAND2xp5_ASAP7_75t_SL g7176 ( 
.A(n_6768),
.B(n_6506),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6826),
.Y(n_7177)
);

INVx1_ASAP7_75t_SL g7178 ( 
.A(n_6871),
.Y(n_7178)
);

CKINVDCx14_ASAP7_75t_R g7179 ( 
.A(n_6757),
.Y(n_7179)
);

INVxp67_ASAP7_75t_L g7180 ( 
.A(n_6757),
.Y(n_7180)
);

INVx2_ASAP7_75t_L g7181 ( 
.A(n_6745),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6745),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6834),
.Y(n_7183)
);

AND2x2_ASAP7_75t_L g7184 ( 
.A(n_6792),
.B(n_6469),
.Y(n_7184)
);

AO21x2_ASAP7_75t_L g7185 ( 
.A1(n_6802),
.A2(n_6359),
.B(n_6353),
.Y(n_7185)
);

AOI21xp5_ASAP7_75t_L g7186 ( 
.A1(n_6838),
.A2(n_6508),
.B(n_6411),
.Y(n_7186)
);

AND2x2_ASAP7_75t_L g7187 ( 
.A(n_6803),
.B(n_6471),
.Y(n_7187)
);

A2O1A1Ixp33_ASAP7_75t_L g7188 ( 
.A1(n_6834),
.A2(n_6573),
.B(n_6411),
.C(n_6484),
.Y(n_7188)
);

OAI21x1_ASAP7_75t_L g7189 ( 
.A1(n_6984),
.A2(n_6465),
.B(n_6429),
.Y(n_7189)
);

HB1xp67_ASAP7_75t_L g7190 ( 
.A(n_6716),
.Y(n_7190)
);

INVx2_ASAP7_75t_L g7191 ( 
.A(n_6803),
.Y(n_7191)
);

AOI21xp33_ASAP7_75t_L g7192 ( 
.A1(n_7090),
.A2(n_7055),
.B(n_6852),
.Y(n_7192)
);

AOI211x1_ASAP7_75t_SL g7193 ( 
.A1(n_6718),
.A2(n_6605),
.B(n_6530),
.C(n_6464),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_6959),
.Y(n_7194)
);

CKINVDCx5p33_ASAP7_75t_R g7195 ( 
.A(n_6901),
.Y(n_7195)
);

AOI21xp33_ASAP7_75t_L g7196 ( 
.A1(n_7090),
.A2(n_6420),
.B(n_6397),
.Y(n_7196)
);

INVx2_ASAP7_75t_L g7197 ( 
.A(n_6857),
.Y(n_7197)
);

OA21x2_ASAP7_75t_L g7198 ( 
.A1(n_6853),
.A2(n_6362),
.B(n_6359),
.Y(n_7198)
);

NAND2xp5_ASAP7_75t_L g7199 ( 
.A(n_6983),
.B(n_6744),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_6983),
.B(n_6475),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6959),
.Y(n_7201)
);

INVx3_ASAP7_75t_L g7202 ( 
.A(n_6969),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_6798),
.B(n_6821),
.Y(n_7203)
);

AOI21xp33_ASAP7_75t_L g7204 ( 
.A1(n_6719),
.A2(n_6516),
.B(n_6512),
.Y(n_7204)
);

INVx1_ASAP7_75t_L g7205 ( 
.A(n_6974),
.Y(n_7205)
);

AND2x2_ASAP7_75t_L g7206 ( 
.A(n_6791),
.B(n_6800),
.Y(n_7206)
);

A2O1A1Ixp33_ASAP7_75t_L g7207 ( 
.A1(n_6853),
.A2(n_6573),
.B(n_6484),
.C(n_6608),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6974),
.Y(n_7208)
);

INVx4_ASAP7_75t_SL g7209 ( 
.A(n_7012),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6744),
.B(n_6689),
.Y(n_7210)
);

INVx2_ASAP7_75t_L g7211 ( 
.A(n_6857),
.Y(n_7211)
);

OR2x2_ASAP7_75t_L g7212 ( 
.A(n_6809),
.B(n_6419),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6975),
.Y(n_7213)
);

INVx2_ASAP7_75t_L g7214 ( 
.A(n_6880),
.Y(n_7214)
);

BUFx3_ASAP7_75t_L g7215 ( 
.A(n_7050),
.Y(n_7215)
);

AND2x2_ASAP7_75t_L g7216 ( 
.A(n_6801),
.B(n_6507),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6975),
.Y(n_7217)
);

INVx1_ASAP7_75t_L g7218 ( 
.A(n_7008),
.Y(n_7218)
);

OAI21x1_ASAP7_75t_L g7219 ( 
.A1(n_6984),
.A2(n_6524),
.B(n_6465),
.Y(n_7219)
);

AOI21xp5_ASAP7_75t_L g7220 ( 
.A1(n_6922),
.A2(n_6453),
.B(n_5918),
.Y(n_7220)
);

INVx5_ASAP7_75t_L g7221 ( 
.A(n_7012),
.Y(n_7221)
);

AOI21xp5_ASAP7_75t_L g7222 ( 
.A1(n_6922),
.A2(n_6453),
.B(n_6618),
.Y(n_7222)
);

NAND2xp5_ASAP7_75t_L g7223 ( 
.A(n_6823),
.B(n_6514),
.Y(n_7223)
);

HB1xp67_ASAP7_75t_L g7224 ( 
.A(n_6708),
.Y(n_7224)
);

AND2x4_ASAP7_75t_L g7225 ( 
.A(n_6895),
.B(n_6982),
.Y(n_7225)
);

INVx3_ASAP7_75t_L g7226 ( 
.A(n_6969),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_7008),
.Y(n_7227)
);

OAI211xp5_ASAP7_75t_L g7228 ( 
.A1(n_7042),
.A2(n_6283),
.B(n_6617),
.C(n_6616),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_7057),
.Y(n_7229)
);

AND2x2_ASAP7_75t_L g7230 ( 
.A(n_6808),
.B(n_6507),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7057),
.Y(n_7231)
);

INVx2_ASAP7_75t_L g7232 ( 
.A(n_6880),
.Y(n_7232)
);

AND2x2_ASAP7_75t_L g7233 ( 
.A(n_6810),
.B(n_6811),
.Y(n_7233)
);

INVx2_ASAP7_75t_SL g7234 ( 
.A(n_6796),
.Y(n_7234)
);

OR2x6_ASAP7_75t_L g7235 ( 
.A(n_7050),
.B(n_5642),
.Y(n_7235)
);

INVx2_ASAP7_75t_L g7236 ( 
.A(n_6964),
.Y(n_7236)
);

HB1xp67_ASAP7_75t_L g7237 ( 
.A(n_7021),
.Y(n_7237)
);

OAI21x1_ASAP7_75t_L g7238 ( 
.A1(n_7107),
.A2(n_6524),
.B(n_6465),
.Y(n_7238)
);

AND2x4_ASAP7_75t_L g7239 ( 
.A(n_6895),
.B(n_6566),
.Y(n_7239)
);

AOI21xp5_ASAP7_75t_L g7240 ( 
.A1(n_7042),
.A2(n_6529),
.B(n_6507),
.Y(n_7240)
);

INVx4_ASAP7_75t_SL g7241 ( 
.A(n_7012),
.Y(n_7241)
);

OAI21xp5_ASAP7_75t_SL g7242 ( 
.A1(n_7059),
.A2(n_6671),
.B(n_6529),
.Y(n_7242)
);

NAND3xp33_ASAP7_75t_L g7243 ( 
.A(n_6752),
.B(n_6604),
.C(n_6466),
.Y(n_7243)
);

AND2x2_ASAP7_75t_L g7244 ( 
.A(n_6813),
.B(n_6529),
.Y(n_7244)
);

INVx3_ASAP7_75t_L g7245 ( 
.A(n_6969),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_7061),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_6823),
.B(n_6417),
.Y(n_7247)
);

NAND3xp33_ASAP7_75t_SL g7248 ( 
.A(n_7119),
.B(n_6515),
.C(n_6470),
.Y(n_7248)
);

INVx2_ASAP7_75t_L g7249 ( 
.A(n_6964),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_6819),
.B(n_6692),
.Y(n_7250)
);

AND2x2_ASAP7_75t_L g7251 ( 
.A(n_6787),
.B(n_6692),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_7061),
.Y(n_7252)
);

HB1xp67_ASAP7_75t_L g7253 ( 
.A(n_7021),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_6862),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_6833),
.B(n_6782),
.Y(n_7255)
);

INVx2_ASAP7_75t_L g7256 ( 
.A(n_7107),
.Y(n_7256)
);

A2O1A1Ixp33_ASAP7_75t_L g7257 ( 
.A1(n_7067),
.A2(n_5980),
.B(n_6650),
.C(n_6613),
.Y(n_7257)
);

NAND2xp5_ASAP7_75t_L g7258 ( 
.A(n_6833),
.B(n_6417),
.Y(n_7258)
);

INVx2_ASAP7_75t_L g7259 ( 
.A(n_6982),
.Y(n_7259)
);

OR2x6_ASAP7_75t_L g7260 ( 
.A(n_7000),
.B(n_5301),
.Y(n_7260)
);

AND2x2_ASAP7_75t_L g7261 ( 
.A(n_6788),
.B(n_6699),
.Y(n_7261)
);

A2O1A1Ixp33_ASAP7_75t_L g7262 ( 
.A1(n_7067),
.A2(n_6613),
.B(n_6650),
.C(n_5961),
.Y(n_7262)
);

BUFx3_ASAP7_75t_L g7263 ( 
.A(n_6759),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_6862),
.Y(n_7264)
);

A2O1A1Ixp33_ASAP7_75t_L g7265 ( 
.A1(n_6804),
.A2(n_6650),
.B(n_6613),
.C(n_6547),
.Y(n_7265)
);

AND2x2_ASAP7_75t_L g7266 ( 
.A(n_6845),
.B(n_6680),
.Y(n_7266)
);

AND2x2_ASAP7_75t_L g7267 ( 
.A(n_6849),
.B(n_6680),
.Y(n_7267)
);

INVx2_ASAP7_75t_SL g7268 ( 
.A(n_6749),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_6784),
.B(n_6478),
.Y(n_7269)
);

INVx2_ASAP7_75t_SL g7270 ( 
.A(n_6749),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_7000),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6752),
.Y(n_7272)
);

NOR3xp33_ASAP7_75t_L g7273 ( 
.A(n_6828),
.B(n_6528),
.C(n_6524),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_6762),
.Y(n_7274)
);

HB1xp67_ASAP7_75t_L g7275 ( 
.A(n_6762),
.Y(n_7275)
);

AND2x2_ASAP7_75t_L g7276 ( 
.A(n_6704),
.B(n_6682),
.Y(n_7276)
);

AND2x2_ASAP7_75t_L g7277 ( 
.A(n_6736),
.B(n_6682),
.Y(n_7277)
);

NAND2xp5_ASAP7_75t_L g7278 ( 
.A(n_6985),
.B(n_6478),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_6804),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_6739),
.B(n_6681),
.Y(n_7280)
);

OAI21x1_ASAP7_75t_L g7281 ( 
.A1(n_6905),
.A2(n_6544),
.B(n_6528),
.Y(n_7281)
);

OAI21xp33_ASAP7_75t_L g7282 ( 
.A1(n_6828),
.A2(n_6505),
.B(n_6442),
.Y(n_7282)
);

AND2x4_ASAP7_75t_L g7283 ( 
.A(n_6867),
.B(n_6566),
.Y(n_7283)
);

BUFx2_ASAP7_75t_L g7284 ( 
.A(n_6749),
.Y(n_7284)
);

OAI21xp5_ASAP7_75t_L g7285 ( 
.A1(n_7117),
.A2(n_6539),
.B(n_6514),
.Y(n_7285)
);

OAI21xp5_ASAP7_75t_L g7286 ( 
.A1(n_6957),
.A2(n_6539),
.B(n_6555),
.Y(n_7286)
);

INVxp67_ASAP7_75t_L g7287 ( 
.A(n_6891),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_6836),
.B(n_6681),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_6867),
.B(n_6699),
.Y(n_7289)
);

AOI21xp5_ASAP7_75t_L g7290 ( 
.A1(n_6891),
.A2(n_6539),
.B(n_6543),
.Y(n_7290)
);

AOI21x1_ASAP7_75t_L g7291 ( 
.A1(n_6840),
.A2(n_6516),
.B(n_6512),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_6805),
.Y(n_7292)
);

NOR2xp33_ASAP7_75t_L g7293 ( 
.A(n_6893),
.B(n_5123),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_6805),
.Y(n_7294)
);

CKINVDCx20_ASAP7_75t_R g7295 ( 
.A(n_6773),
.Y(n_7295)
);

INVx1_ASAP7_75t_L g7296 ( 
.A(n_6818),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_6715),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6719),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6725),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_6725),
.Y(n_7300)
);

AND2x4_ASAP7_75t_L g7301 ( 
.A(n_6977),
.B(n_6566),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7037),
.Y(n_7302)
);

CKINVDCx14_ASAP7_75t_R g7303 ( 
.A(n_6843),
.Y(n_7303)
);

AND2x4_ASAP7_75t_L g7304 ( 
.A(n_7007),
.B(n_6636),
.Y(n_7304)
);

INVx2_ASAP7_75t_L g7305 ( 
.A(n_6893),
.Y(n_7305)
);

OR2x2_ASAP7_75t_L g7306 ( 
.A(n_6729),
.B(n_6385),
.Y(n_7306)
);

AO21x2_ASAP7_75t_L g7307 ( 
.A1(n_6917),
.A2(n_6369),
.B(n_6367),
.Y(n_7307)
);

INVx1_ASAP7_75t_L g7308 ( 
.A(n_7037),
.Y(n_7308)
);

NOR2xp33_ASAP7_75t_L g7309 ( 
.A(n_6945),
.B(n_7001),
.Y(n_7309)
);

CKINVDCx5p33_ASAP7_75t_R g7310 ( 
.A(n_6846),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_SL g7311 ( 
.A(n_6768),
.B(n_6636),
.Y(n_7311)
);

OA21x2_ASAP7_75t_L g7312 ( 
.A1(n_6714),
.A2(n_6367),
.B(n_6362),
.Y(n_7312)
);

OA21x2_ASAP7_75t_L g7313 ( 
.A1(n_6720),
.A2(n_6369),
.B(n_6370),
.Y(n_7313)
);

AND2x2_ASAP7_75t_L g7314 ( 
.A(n_6769),
.B(n_6746),
.Y(n_7314)
);

NAND2xp5_ASAP7_75t_L g7315 ( 
.A(n_6988),
.B(n_6691),
.Y(n_7315)
);

NAND2xp5_ASAP7_75t_L g7316 ( 
.A(n_7015),
.B(n_6698),
.Y(n_7316)
);

AOI21xp5_ASAP7_75t_L g7317 ( 
.A1(n_7059),
.A2(n_6547),
.B(n_6543),
.Y(n_7317)
);

INVx4_ASAP7_75t_L g7318 ( 
.A(n_7012),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_7054),
.Y(n_7319)
);

AND2x2_ASAP7_75t_L g7320 ( 
.A(n_6741),
.B(n_6636),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_7054),
.Y(n_7321)
);

AND2x4_ASAP7_75t_L g7322 ( 
.A(n_7034),
.B(n_7038),
.Y(n_7322)
);

OA21x2_ASAP7_75t_L g7323 ( 
.A1(n_6721),
.A2(n_6386),
.B(n_6370),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7096),
.Y(n_7324)
);

AND2x4_ASAP7_75t_L g7325 ( 
.A(n_6945),
.B(n_6555),
.Y(n_7325)
);

OAI21x1_ASAP7_75t_L g7326 ( 
.A1(n_7060),
.A2(n_6544),
.B(n_6528),
.Y(n_7326)
);

AO21x2_ASAP7_75t_L g7327 ( 
.A1(n_6917),
.A2(n_6389),
.B(n_6386),
.Y(n_7327)
);

NAND2xp5_ASAP7_75t_L g7328 ( 
.A(n_7019),
.B(n_6545),
.Y(n_7328)
);

INVx2_ASAP7_75t_L g7329 ( 
.A(n_7001),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_6742),
.B(n_6489),
.Y(n_7330)
);

INVx2_ASAP7_75t_L g7331 ( 
.A(n_7101),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_7096),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_6812),
.B(n_6545),
.Y(n_7333)
);

NAND4xp25_ASAP7_75t_L g7334 ( 
.A(n_6751),
.B(n_6671),
.C(n_6575),
.D(n_6544),
.Y(n_7334)
);

OA21x2_ASAP7_75t_L g7335 ( 
.A1(n_6724),
.A2(n_6389),
.B(n_6472),
.Y(n_7335)
);

NAND2xp5_ASAP7_75t_L g7336 ( 
.A(n_6765),
.B(n_6545),
.Y(n_7336)
);

AOI21xp5_ASAP7_75t_L g7337 ( 
.A1(n_6902),
.A2(n_6550),
.B(n_6548),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_7101),
.Y(n_7338)
);

AOI21xp5_ASAP7_75t_L g7339 ( 
.A1(n_6902),
.A2(n_6550),
.B(n_6548),
.Y(n_7339)
);

INVxp67_ASAP7_75t_SL g7340 ( 
.A(n_6751),
.Y(n_7340)
);

INVx3_ASAP7_75t_L g7341 ( 
.A(n_7063),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_6832),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6844),
.Y(n_7343)
);

BUFx2_ASAP7_75t_L g7344 ( 
.A(n_6980),
.Y(n_7344)
);

NOR2x1_ASAP7_75t_L g7345 ( 
.A(n_7095),
.B(n_6575),
.Y(n_7345)
);

NAND2xp5_ASAP7_75t_L g7346 ( 
.A(n_6701),
.B(n_6545),
.Y(n_7346)
);

AND2x4_ASAP7_75t_L g7347 ( 
.A(n_6756),
.B(n_5393),
.Y(n_7347)
);

AO21x2_ASAP7_75t_L g7348 ( 
.A1(n_6980),
.A2(n_6856),
.B(n_6847),
.Y(n_7348)
);

NOR2xp33_ASAP7_75t_L g7349 ( 
.A(n_6846),
.B(n_5637),
.Y(n_7349)
);

OAI21x1_ASAP7_75t_L g7350 ( 
.A1(n_7069),
.A2(n_6575),
.B(n_6247),
.Y(n_7350)
);

INVx3_ASAP7_75t_L g7351 ( 
.A(n_7063),
.Y(n_7351)
);

AOI21xp5_ASAP7_75t_L g7352 ( 
.A1(n_6904),
.A2(n_6563),
.B(n_6559),
.Y(n_7352)
);

AND2x2_ASAP7_75t_L g7353 ( 
.A(n_6748),
.B(n_6489),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_6859),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_SL g7355 ( 
.A(n_6753),
.B(n_6070),
.Y(n_7355)
);

AND2x2_ASAP7_75t_L g7356 ( 
.A(n_7078),
.B(n_5582),
.Y(n_7356)
);

INVx2_ASAP7_75t_L g7357 ( 
.A(n_7095),
.Y(n_7357)
);

OR2x2_ASAP7_75t_L g7358 ( 
.A(n_6783),
.B(n_5816),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_6860),
.Y(n_7359)
);

INVx2_ASAP7_75t_L g7360 ( 
.A(n_6753),
.Y(n_7360)
);

BUFx2_ASAP7_75t_L g7361 ( 
.A(n_6764),
.Y(n_7361)
);

AOI21xp5_ASAP7_75t_L g7362 ( 
.A1(n_6904),
.A2(n_6563),
.B(n_6559),
.Y(n_7362)
);

INVx2_ASAP7_75t_L g7363 ( 
.A(n_6764),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6897),
.Y(n_7364)
);

HB1xp67_ASAP7_75t_L g7365 ( 
.A(n_6740),
.Y(n_7365)
);

AOI21xp5_ASAP7_75t_L g7366 ( 
.A1(n_7119),
.A2(n_6587),
.B(n_6615),
.Y(n_7366)
);

AND2x2_ASAP7_75t_L g7367 ( 
.A(n_7113),
.B(n_5582),
.Y(n_7367)
);

INVx2_ASAP7_75t_L g7368 ( 
.A(n_6919),
.Y(n_7368)
);

AO21x2_ASAP7_75t_L g7369 ( 
.A1(n_6897),
.A2(n_6533),
.B(n_6531),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_6907),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_6907),
.Y(n_7371)
);

BUFx2_ASAP7_75t_L g7372 ( 
.A(n_6763),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6919),
.Y(n_7373)
);

INVx3_ASAP7_75t_L g7374 ( 
.A(n_7063),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_6842),
.B(n_5646),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6909),
.Y(n_7376)
);

INVxp67_ASAP7_75t_L g7377 ( 
.A(n_7013),
.Y(n_7377)
);

OR2x2_ASAP7_75t_L g7378 ( 
.A(n_7036),
.B(n_6115),
.Y(n_7378)
);

INVx2_ASAP7_75t_L g7379 ( 
.A(n_6952),
.Y(n_7379)
);

AND2x2_ASAP7_75t_L g7380 ( 
.A(n_6747),
.B(n_6770),
.Y(n_7380)
);

AND2x6_ASAP7_75t_SL g7381 ( 
.A(n_7010),
.B(n_5577),
.Y(n_7381)
);

OA21x2_ASAP7_75t_L g7382 ( 
.A1(n_6727),
.A2(n_6477),
.B(n_6472),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6909),
.Y(n_7383)
);

AND2x2_ASAP7_75t_L g7384 ( 
.A(n_6780),
.B(n_5646),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_6998),
.Y(n_7385)
);

NAND4xp25_ASAP7_75t_L g7386 ( 
.A(n_7010),
.B(n_6531),
.C(n_6533),
.D(n_4936),
.Y(n_7386)
);

OA21x2_ASAP7_75t_L g7387 ( 
.A1(n_6734),
.A2(n_6486),
.B(n_6477),
.Y(n_7387)
);

INVx1_ASAP7_75t_SL g7388 ( 
.A(n_6723),
.Y(n_7388)
);

NOR2xp33_ASAP7_75t_L g7389 ( 
.A(n_6918),
.B(n_5637),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_6998),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_7004),
.Y(n_7391)
);

INVx3_ASAP7_75t_L g7392 ( 
.A(n_6952),
.Y(n_7392)
);

NAND3xp33_ASAP7_75t_L g7393 ( 
.A(n_7075),
.B(n_6628),
.C(n_6615),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_6705),
.B(n_6628),
.Y(n_7394)
);

HB1xp67_ASAP7_75t_L g7395 ( 
.A(n_6706),
.Y(n_7395)
);

BUFx8_ASAP7_75t_L g7396 ( 
.A(n_6890),
.Y(n_7396)
);

AND3x2_ASAP7_75t_L g7397 ( 
.A(n_7075),
.B(n_6632),
.C(n_6630),
.Y(n_7397)
);

AND2x2_ASAP7_75t_L g7398 ( 
.A(n_6900),
.B(n_5646),
.Y(n_7398)
);

INVxp67_ASAP7_75t_SL g7399 ( 
.A(n_6817),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_7004),
.Y(n_7400)
);

BUFx3_ASAP7_75t_L g7401 ( 
.A(n_6735),
.Y(n_7401)
);

INVx1_ASAP7_75t_L g7402 ( 
.A(n_7030),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_7030),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_6772),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_6981),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_6772),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_6774),
.Y(n_7407)
);

AO21x2_ASAP7_75t_L g7408 ( 
.A1(n_6737),
.A2(n_6424),
.B(n_6421),
.Y(n_7408)
);

OAI21x1_ASAP7_75t_L g7409 ( 
.A1(n_7070),
.A2(n_6247),
.B(n_6630),
.Y(n_7409)
);

AO21x2_ASAP7_75t_L g7410 ( 
.A1(n_6738),
.A2(n_6424),
.B(n_6421),
.Y(n_7410)
);

OAI21xp5_ASAP7_75t_SL g7411 ( 
.A1(n_6931),
.A2(n_5358),
.B(n_5300),
.Y(n_7411)
);

OAI21x1_ASAP7_75t_L g7412 ( 
.A1(n_7081),
.A2(n_6635),
.B(n_6632),
.Y(n_7412)
);

INVx1_ASAP7_75t_L g7413 ( 
.A(n_6774),
.Y(n_7413)
);

INVx2_ASAP7_75t_L g7414 ( 
.A(n_6981),
.Y(n_7414)
);

OR2x6_ASAP7_75t_L g7415 ( 
.A(n_6892),
.B(n_5301),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_6778),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_6778),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6781),
.Y(n_7418)
);

AND2x2_ASAP7_75t_L g7419 ( 
.A(n_6963),
.B(n_5646),
.Y(n_7419)
);

AOI21xp5_ASAP7_75t_L g7420 ( 
.A1(n_6817),
.A2(n_6637),
.B(n_6635),
.Y(n_7420)
);

AO21x2_ASAP7_75t_L g7421 ( 
.A1(n_6777),
.A2(n_6438),
.B(n_6435),
.Y(n_7421)
);

BUFx3_ASAP7_75t_L g7422 ( 
.A(n_7002),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6781),
.Y(n_7423)
);

NOR2xp33_ASAP7_75t_L g7424 ( 
.A(n_6925),
.B(n_5374),
.Y(n_7424)
);

INVx4_ASAP7_75t_R g7425 ( 
.A(n_7003),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_6797),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6797),
.Y(n_7427)
);

OR2x2_ASAP7_75t_L g7428 ( 
.A(n_6967),
.B(n_6159),
.Y(n_7428)
);

AND2x2_ASAP7_75t_L g7429 ( 
.A(n_6965),
.B(n_5677),
.Y(n_7429)
);

NOR2xp33_ASAP7_75t_L g7430 ( 
.A(n_6926),
.B(n_5374),
.Y(n_7430)
);

NAND2xp5_ASAP7_75t_L g7431 ( 
.A(n_6927),
.B(n_6637),
.Y(n_7431)
);

INVx2_ASAP7_75t_L g7432 ( 
.A(n_6996),
.Y(n_7432)
);

INVxp67_ASAP7_75t_SL g7433 ( 
.A(n_7006),
.Y(n_7433)
);

OAI31xp33_ASAP7_75t_SL g7434 ( 
.A1(n_6839),
.A2(n_6882),
.A3(n_6896),
.B(n_6876),
.Y(n_7434)
);

BUFx3_ASAP7_75t_L g7435 ( 
.A(n_7011),
.Y(n_7435)
);

INVx2_ASAP7_75t_SL g7436 ( 
.A(n_6996),
.Y(n_7436)
);

INVx2_ASAP7_75t_L g7437 ( 
.A(n_7087),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_6822),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_6822),
.Y(n_7439)
);

HB1xp67_ASAP7_75t_L g7440 ( 
.A(n_6928),
.Y(n_7440)
);

NOR2x1p5_ASAP7_75t_L g7441 ( 
.A(n_6837),
.B(n_4936),
.Y(n_7441)
);

OAI21xp5_ASAP7_75t_L g7442 ( 
.A1(n_6733),
.A2(n_6645),
.B(n_6644),
.Y(n_7442)
);

NAND2xp5_ASAP7_75t_L g7443 ( 
.A(n_6865),
.B(n_6644),
.Y(n_7443)
);

INVx3_ASAP7_75t_L g7444 ( 
.A(n_6839),
.Y(n_7444)
);

INVx4_ASAP7_75t_L g7445 ( 
.A(n_6763),
.Y(n_7445)
);

A2O1A1Ixp33_ASAP7_75t_L g7446 ( 
.A1(n_6743),
.A2(n_6645),
.B(n_5379),
.C(n_5415),
.Y(n_7446)
);

NAND2xp5_ASAP7_75t_L g7447 ( 
.A(n_6920),
.B(n_6439),
.Y(n_7447)
);

INVx5_ASAP7_75t_L g7448 ( 
.A(n_6763),
.Y(n_7448)
);

AND2x2_ASAP7_75t_L g7449 ( 
.A(n_6709),
.B(n_5677),
.Y(n_7449)
);

OA21x2_ASAP7_75t_L g7450 ( 
.A1(n_6779),
.A2(n_6498),
.B(n_6486),
.Y(n_7450)
);

AOI22xp5_ASAP7_75t_L g7451 ( 
.A1(n_6712),
.A2(n_5476),
.B1(n_5951),
.B2(n_5936),
.Y(n_7451)
);

INVx2_ASAP7_75t_L g7452 ( 
.A(n_7087),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_L g7453 ( 
.A(n_6921),
.B(n_6459),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_6711),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_6848),
.Y(n_7455)
);

INVx4_ASAP7_75t_SL g7456 ( 
.A(n_6934),
.Y(n_7456)
);

INVx5_ASAP7_75t_L g7457 ( 
.A(n_6934),
.Y(n_7457)
);

INVx2_ASAP7_75t_L g7458 ( 
.A(n_6711),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_6970),
.B(n_5677),
.Y(n_7459)
);

AND2x2_ASAP7_75t_L g7460 ( 
.A(n_6978),
.B(n_5677),
.Y(n_7460)
);

INVx2_ASAP7_75t_L g7461 ( 
.A(n_6966),
.Y(n_7461)
);

AND2x2_ASAP7_75t_L g7462 ( 
.A(n_6934),
.B(n_5707),
.Y(n_7462)
);

BUFx2_ASAP7_75t_L g7463 ( 
.A(n_6876),
.Y(n_7463)
);

INVx2_ASAP7_75t_L g7464 ( 
.A(n_6968),
.Y(n_7464)
);

OA21x2_ASAP7_75t_L g7465 ( 
.A1(n_6785),
.A2(n_6499),
.B(n_6498),
.Y(n_7465)
);

BUFx2_ASAP7_75t_L g7466 ( 
.A(n_6882),
.Y(n_7466)
);

INVx2_ASAP7_75t_L g7467 ( 
.A(n_6841),
.Y(n_7467)
);

INVxp67_ASAP7_75t_L g7468 ( 
.A(n_6713),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_6848),
.Y(n_7469)
);

HB1xp67_ASAP7_75t_L g7470 ( 
.A(n_7084),
.Y(n_7470)
);

A2O1A1Ixp33_ASAP7_75t_L g7471 ( 
.A1(n_6743),
.A2(n_5379),
.B(n_5415),
.C(n_5402),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_6789),
.Y(n_7472)
);

NAND2xp5_ASAP7_75t_SL g7473 ( 
.A(n_6830),
.B(n_5618),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6790),
.Y(n_7474)
);

INVxp67_ASAP7_75t_SL g7475 ( 
.A(n_7120),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_6793),
.Y(n_7476)
);

INVxp67_ASAP7_75t_L g7477 ( 
.A(n_6722),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_6794),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_6795),
.Y(n_7479)
);

INVx2_ASAP7_75t_L g7480 ( 
.A(n_6896),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_6971),
.B(n_6160),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_6799),
.Y(n_7482)
);

INVx1_ASAP7_75t_L g7483 ( 
.A(n_6806),
.Y(n_7483)
);

OA211x2_ASAP7_75t_L g7484 ( 
.A1(n_7153),
.A2(n_6861),
.B(n_6850),
.C(n_6758),
.Y(n_7484)
);

AND2x2_ASAP7_75t_L g7485 ( 
.A(n_7347),
.B(n_7048),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7158),
.Y(n_7486)
);

AND2x2_ASAP7_75t_L g7487 ( 
.A(n_7347),
.B(n_6855),
.Y(n_7487)
);

NOR2xp33_ASAP7_75t_L g7488 ( 
.A(n_7179),
.B(n_7026),
.Y(n_7488)
);

INVx2_ASAP7_75t_L g7489 ( 
.A(n_7295),
.Y(n_7489)
);

INVx2_ASAP7_75t_SL g7490 ( 
.A(n_7396),
.Y(n_7490)
);

NOR3xp33_ASAP7_75t_L g7491 ( 
.A(n_7145),
.B(n_6771),
.C(n_6766),
.Y(n_7491)
);

AOI21xp5_ASAP7_75t_L g7492 ( 
.A1(n_7141),
.A2(n_6861),
.B(n_6850),
.Y(n_7492)
);

HB1xp67_ASAP7_75t_L g7493 ( 
.A(n_7348),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_7287),
.B(n_6807),
.Y(n_7494)
);

OAI211xp5_ASAP7_75t_SL g7495 ( 
.A1(n_7193),
.A2(n_6820),
.B(n_6824),
.C(n_6814),
.Y(n_7495)
);

NAND3xp33_ASAP7_75t_L g7496 ( 
.A(n_7192),
.B(n_6831),
.C(n_6976),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_7178),
.B(n_7088),
.Y(n_7497)
);

NAND3xp33_ASAP7_75t_L g7498 ( 
.A(n_7123),
.B(n_7076),
.C(n_6976),
.Y(n_7498)
);

NAND2xp5_ASAP7_75t_L g7499 ( 
.A(n_7377),
.B(n_7105),
.Y(n_7499)
);

INVx2_ASAP7_75t_L g7500 ( 
.A(n_7444),
.Y(n_7500)
);

NAND3xp33_ASAP7_75t_L g7501 ( 
.A(n_7143),
.B(n_7076),
.C(n_6870),
.Y(n_7501)
);

AOI211xp5_ASAP7_75t_L g7502 ( 
.A1(n_7140),
.A2(n_7124),
.B(n_7135),
.C(n_7222),
.Y(n_7502)
);

AND2x2_ASAP7_75t_L g7503 ( 
.A(n_7206),
.B(n_6866),
.Y(n_7503)
);

AND2x2_ASAP7_75t_L g7504 ( 
.A(n_7233),
.B(n_6875),
.Y(n_7504)
);

AND2x2_ASAP7_75t_L g7505 ( 
.A(n_7361),
.B(n_6881),
.Y(n_7505)
);

NOR3xp33_ASAP7_75t_L g7506 ( 
.A(n_7125),
.B(n_7137),
.C(n_7196),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_7275),
.Y(n_7507)
);

OR2x2_ASAP7_75t_L g7508 ( 
.A(n_7296),
.B(n_6851),
.Y(n_7508)
);

AND2x4_ASAP7_75t_L g7509 ( 
.A(n_7133),
.B(n_6899),
.Y(n_7509)
);

AOI22xp5_ASAP7_75t_L g7510 ( 
.A1(n_7348),
.A2(n_6758),
.B1(n_6767),
.B2(n_6750),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7237),
.Y(n_7511)
);

AOI22xp5_ASAP7_75t_L g7512 ( 
.A1(n_7142),
.A2(n_6767),
.B1(n_6750),
.B2(n_6863),
.Y(n_7512)
);

NOR2xp33_ASAP7_75t_L g7513 ( 
.A(n_7126),
.B(n_7026),
.Y(n_7513)
);

AOI22xp33_ASAP7_75t_L g7514 ( 
.A1(n_7186),
.A2(n_6438),
.B1(n_6440),
.B2(n_6435),
.Y(n_7514)
);

INVx2_ASAP7_75t_L g7515 ( 
.A(n_7444),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_7148),
.Y(n_7516)
);

NAND4xp75_ASAP7_75t_L g7517 ( 
.A(n_7129),
.B(n_6816),
.C(n_6960),
.D(n_6827),
.Y(n_7517)
);

OAI21xp5_ASAP7_75t_L g7518 ( 
.A1(n_7207),
.A2(n_6960),
.B(n_6816),
.Y(n_7518)
);

AND2x2_ASAP7_75t_L g7519 ( 
.A(n_7203),
.B(n_6885),
.Y(n_7519)
);

AO21x2_ASAP7_75t_L g7520 ( 
.A1(n_7134),
.A2(n_7136),
.B(n_7139),
.Y(n_7520)
);

NOR3xp33_ASAP7_75t_L g7521 ( 
.A(n_7169),
.B(n_6835),
.C(n_6815),
.Y(n_7521)
);

NAND4xp75_ASAP7_75t_L g7522 ( 
.A(n_7128),
.B(n_6872),
.C(n_6889),
.D(n_6864),
.Y(n_7522)
);

OR2x2_ASAP7_75t_L g7523 ( 
.A(n_7296),
.B(n_6829),
.Y(n_7523)
);

NAND3xp33_ASAP7_75t_L g7524 ( 
.A(n_7397),
.B(n_7024),
.C(n_7022),
.Y(n_7524)
);

INVx2_ASAP7_75t_L g7525 ( 
.A(n_7392),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_7310),
.B(n_7322),
.Y(n_7526)
);

AO21x2_ASAP7_75t_L g7527 ( 
.A1(n_7134),
.A2(n_7136),
.B(n_7139),
.Y(n_7527)
);

AND2x2_ASAP7_75t_L g7528 ( 
.A(n_7216),
.B(n_6886),
.Y(n_7528)
);

AND2x2_ASAP7_75t_L g7529 ( 
.A(n_7230),
.B(n_7244),
.Y(n_7529)
);

AND2x2_ASAP7_75t_L g7530 ( 
.A(n_7380),
.B(n_6899),
.Y(n_7530)
);

NAND2xp5_ASAP7_75t_L g7531 ( 
.A(n_7322),
.B(n_6989),
.Y(n_7531)
);

AND2x2_ASAP7_75t_L g7532 ( 
.A(n_7280),
.B(n_6912),
.Y(n_7532)
);

NOR2xp33_ASAP7_75t_L g7533 ( 
.A(n_7126),
.B(n_7062),
.Y(n_7533)
);

AND2x2_ASAP7_75t_L g7534 ( 
.A(n_7314),
.B(n_6912),
.Y(n_7534)
);

NAND4xp25_ASAP7_75t_L g7535 ( 
.A(n_7434),
.B(n_7014),
.C(n_7062),
.D(n_7040),
.Y(n_7535)
);

OAI211xp5_ASAP7_75t_SL g7536 ( 
.A1(n_7242),
.A2(n_7104),
.B(n_7114),
.C(n_7092),
.Y(n_7536)
);

INVxp67_ASAP7_75t_SL g7537 ( 
.A(n_7396),
.Y(n_7537)
);

AND2x2_ASAP7_75t_L g7538 ( 
.A(n_7235),
.B(n_6931),
.Y(n_7538)
);

INVxp67_ASAP7_75t_SL g7539 ( 
.A(n_7149),
.Y(n_7539)
);

INVx3_ASAP7_75t_L g7540 ( 
.A(n_7283),
.Y(n_7540)
);

HB1xp67_ASAP7_75t_L g7541 ( 
.A(n_7395),
.Y(n_7541)
);

NAND2xp5_ASAP7_75t_L g7542 ( 
.A(n_7433),
.B(n_7047),
.Y(n_7542)
);

OR2x2_ASAP7_75t_L g7543 ( 
.A(n_7297),
.B(n_7110),
.Y(n_7543)
);

AND2x2_ASAP7_75t_SL g7544 ( 
.A(n_7344),
.B(n_6979),
.Y(n_7544)
);

NAND2xp5_ASAP7_75t_L g7545 ( 
.A(n_7149),
.B(n_6873),
.Y(n_7545)
);

NAND3xp33_ASAP7_75t_L g7546 ( 
.A(n_7273),
.B(n_6955),
.C(n_6944),
.Y(n_7546)
);

BUFx3_ASAP7_75t_L g7547 ( 
.A(n_7215),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7235),
.B(n_6979),
.Y(n_7548)
);

AOI22xp33_ASAP7_75t_L g7549 ( 
.A1(n_7292),
.A2(n_6441),
.B1(n_6452),
.B2(n_6440),
.Y(n_7549)
);

OAI22xp5_ASAP7_75t_L g7550 ( 
.A1(n_7388),
.A2(n_5839),
.B1(n_7097),
.B2(n_7031),
.Y(n_7550)
);

NAND3xp33_ASAP7_75t_L g7551 ( 
.A(n_7195),
.B(n_6972),
.C(n_7065),
.Y(n_7551)
);

NOR2xp33_ASAP7_75t_L g7552 ( 
.A(n_7303),
.B(n_6830),
.Y(n_7552)
);

AO21x2_ASAP7_75t_L g7553 ( 
.A1(n_7127),
.A2(n_6868),
.B(n_6923),
.Y(n_7553)
);

INVxp67_ASAP7_75t_L g7554 ( 
.A(n_7349),
.Y(n_7554)
);

OR2x2_ASAP7_75t_L g7555 ( 
.A(n_7297),
.B(n_6868),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_7288),
.B(n_7016),
.Y(n_7556)
);

NOR3xp33_ASAP7_75t_L g7557 ( 
.A(n_7202),
.B(n_6877),
.C(n_6874),
.Y(n_7557)
);

AOI221xp5_ASAP7_75t_L g7558 ( 
.A1(n_7188),
.A2(n_7106),
.B1(n_7108),
.B2(n_7103),
.C(n_7098),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_7253),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_7440),
.B(n_6878),
.Y(n_7560)
);

AOI221xp5_ASAP7_75t_L g7561 ( 
.A1(n_7317),
.A2(n_7118),
.B1(n_7121),
.B2(n_7111),
.C(n_7109),
.Y(n_7561)
);

OAI221xp5_ASAP7_75t_SL g7562 ( 
.A1(n_7147),
.A2(n_6906),
.B1(n_6914),
.B2(n_6910),
.C(n_6888),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_7122),
.Y(n_7563)
);

NAND2xp5_ASAP7_75t_L g7564 ( 
.A(n_7224),
.B(n_6879),
.Y(n_7564)
);

AO21x2_ASAP7_75t_L g7565 ( 
.A1(n_7127),
.A2(n_6924),
.B(n_6923),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7266),
.B(n_7018),
.Y(n_7566)
);

AOI22xp33_ASAP7_75t_L g7567 ( 
.A1(n_7292),
.A2(n_6452),
.B1(n_6460),
.B2(n_6441),
.Y(n_7567)
);

NOR3xp33_ASAP7_75t_L g7568 ( 
.A(n_7202),
.B(n_7089),
.C(n_7085),
.Y(n_7568)
);

OAI21xp5_ASAP7_75t_L g7569 ( 
.A1(n_7290),
.A2(n_7065),
.B(n_7066),
.Y(n_7569)
);

NAND2xp5_ASAP7_75t_L g7570 ( 
.A(n_7467),
.B(n_6883),
.Y(n_7570)
);

OR2x2_ASAP7_75t_L g7571 ( 
.A(n_7306),
.B(n_7115),
.Y(n_7571)
);

NOR2xp33_ASAP7_75t_L g7572 ( 
.A(n_7283),
.B(n_7116),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7160),
.Y(n_7573)
);

NOR2x1_ASAP7_75t_L g7574 ( 
.A(n_7318),
.B(n_7341),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7162),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7166),
.Y(n_7576)
);

AOI22xp33_ASAP7_75t_L g7577 ( 
.A1(n_7294),
.A2(n_7279),
.B1(n_7198),
.B2(n_7302),
.Y(n_7577)
);

NAND4xp75_ASAP7_75t_L g7578 ( 
.A(n_7150),
.B(n_6915),
.C(n_6930),
.D(n_6908),
.Y(n_7578)
);

AOI22xp33_ASAP7_75t_L g7579 ( 
.A1(n_7294),
.A2(n_6461),
.B1(n_6460),
.B2(n_5959),
.Y(n_7579)
);

AND2x2_ASAP7_75t_L g7580 ( 
.A(n_7267),
.B(n_7025),
.Y(n_7580)
);

NOR3xp33_ASAP7_75t_L g7581 ( 
.A(n_7226),
.B(n_6887),
.C(n_6884),
.Y(n_7581)
);

AO21x2_ASAP7_75t_L g7582 ( 
.A1(n_7131),
.A2(n_6932),
.B(n_6924),
.Y(n_7582)
);

OAI211xp5_ASAP7_75t_L g7583 ( 
.A1(n_7220),
.A2(n_6939),
.B(n_6940),
.C(n_6937),
.Y(n_7583)
);

NAND3xp33_ASAP7_75t_L g7584 ( 
.A(n_7243),
.B(n_7080),
.C(n_6898),
.Y(n_7584)
);

NAND3xp33_ASAP7_75t_L g7585 ( 
.A(n_7393),
.B(n_6903),
.C(n_6894),
.Y(n_7585)
);

OA211x2_ASAP7_75t_L g7586 ( 
.A1(n_7180),
.A2(n_6933),
.B(n_6942),
.C(n_6932),
.Y(n_7586)
);

AND2x2_ASAP7_75t_L g7587 ( 
.A(n_7250),
.B(n_6947),
.Y(n_7587)
);

INVxp33_ASAP7_75t_L g7588 ( 
.A(n_7154),
.Y(n_7588)
);

INVx3_ASAP7_75t_L g7589 ( 
.A(n_7301),
.Y(n_7589)
);

AND2x2_ASAP7_75t_L g7590 ( 
.A(n_7289),
.B(n_6953),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7168),
.Y(n_7591)
);

NAND4xp75_ASAP7_75t_L g7592 ( 
.A(n_7345),
.B(n_6954),
.C(n_6962),
.D(n_7027),
.Y(n_7592)
);

INVx2_ASAP7_75t_L g7593 ( 
.A(n_7392),
.Y(n_7593)
);

NAND3xp33_ASAP7_75t_SL g7594 ( 
.A(n_7240),
.B(n_7041),
.C(n_6991),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_7177),
.Y(n_7595)
);

OR2x2_ASAP7_75t_L g7596 ( 
.A(n_7255),
.B(n_6933),
.Y(n_7596)
);

NAND2xp5_ASAP7_75t_L g7597 ( 
.A(n_7173),
.B(n_7174),
.Y(n_7597)
);

OR2x2_ASAP7_75t_L g7598 ( 
.A(n_7152),
.B(n_7082),
.Y(n_7598)
);

NOR3xp33_ASAP7_75t_L g7599 ( 
.A(n_7226),
.B(n_7079),
.C(n_7074),
.Y(n_7599)
);

BUFx3_ASAP7_75t_L g7600 ( 
.A(n_7422),
.Y(n_7600)
);

OAI221xp5_ASAP7_75t_L g7601 ( 
.A1(n_7265),
.A2(n_5379),
.B1(n_5979),
.B2(n_5959),
.C(n_5951),
.Y(n_7601)
);

NAND3xp33_ASAP7_75t_L g7602 ( 
.A(n_7131),
.B(n_6913),
.C(n_6911),
.Y(n_7602)
);

AOI22xp5_ASAP7_75t_L g7603 ( 
.A1(n_7183),
.A2(n_6916),
.B1(n_6938),
.B2(n_6935),
.Y(n_7603)
);

AND2x2_ASAP7_75t_L g7604 ( 
.A(n_7251),
.B(n_7046),
.Y(n_7604)
);

NAND4xp75_ASAP7_75t_L g7605 ( 
.A(n_7268),
.B(n_6461),
.C(n_6943),
.D(n_6941),
.Y(n_7605)
);

AND2x2_ASAP7_75t_L g7606 ( 
.A(n_7261),
.B(n_7068),
.Y(n_7606)
);

AND2x2_ASAP7_75t_L g7607 ( 
.A(n_7175),
.B(n_7071),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_7312),
.Y(n_7608)
);

NOR3xp33_ASAP7_75t_L g7609 ( 
.A(n_7245),
.B(n_7058),
.C(n_6948),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_7312),
.Y(n_7610)
);

AND2x4_ASAP7_75t_L g7611 ( 
.A(n_7165),
.B(n_7116),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_7313),
.Y(n_7612)
);

NAND4xp75_ASAP7_75t_L g7613 ( 
.A(n_7270),
.B(n_6950),
.C(n_6956),
.D(n_6946),
.Y(n_7613)
);

NOR2xp33_ASAP7_75t_L g7614 ( 
.A(n_7448),
.B(n_7083),
.Y(n_7614)
);

NOR3xp33_ASAP7_75t_L g7615 ( 
.A(n_7245),
.B(n_7318),
.C(n_7248),
.Y(n_7615)
);

NAND2xp5_ASAP7_75t_L g7616 ( 
.A(n_7181),
.B(n_6958),
.Y(n_7616)
);

AND2x2_ASAP7_75t_L g7617 ( 
.A(n_7276),
.B(n_7077),
.Y(n_7617)
);

OAI221xp5_ASAP7_75t_SL g7618 ( 
.A1(n_7172),
.A2(n_5436),
.B1(n_5468),
.B2(n_5415),
.C(n_5402),
.Y(n_7618)
);

OA211x2_ASAP7_75t_L g7619 ( 
.A1(n_7424),
.A2(n_7430),
.B(n_7293),
.C(n_7389),
.Y(n_7619)
);

CKINVDCx5p33_ASAP7_75t_R g7620 ( 
.A(n_7381),
.Y(n_7620)
);

NOR3xp33_ASAP7_75t_L g7621 ( 
.A(n_7284),
.B(n_6973),
.C(n_6961),
.Y(n_7621)
);

AND2x2_ASAP7_75t_L g7622 ( 
.A(n_7277),
.B(n_7099),
.Y(n_7622)
);

AOI22xp33_ASAP7_75t_L g7623 ( 
.A1(n_7198),
.A2(n_5982),
.B1(n_5988),
.B2(n_5979),
.Y(n_7623)
);

NAND3xp33_ASAP7_75t_SL g7624 ( 
.A(n_7228),
.B(n_7286),
.C(n_7285),
.Y(n_7624)
);

OR2x2_ASAP7_75t_L g7625 ( 
.A(n_7359),
.B(n_7115),
.Y(n_7625)
);

NOR2x1_ASAP7_75t_L g7626 ( 
.A(n_7341),
.B(n_7351),
.Y(n_7626)
);

INVx2_ASAP7_75t_L g7627 ( 
.A(n_7463),
.Y(n_7627)
);

INVx2_ASAP7_75t_L g7628 ( 
.A(n_7466),
.Y(n_7628)
);

OA211x2_ASAP7_75t_L g7629 ( 
.A1(n_7309),
.A2(n_6949),
.B(n_6992),
.C(n_6942),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_7320),
.B(n_7045),
.Y(n_7630)
);

AND2x2_ASAP7_75t_L g7631 ( 
.A(n_7184),
.B(n_7052),
.Y(n_7631)
);

AND2x2_ASAP7_75t_L g7632 ( 
.A(n_7330),
.B(n_7435),
.Y(n_7632)
);

NAND4xp75_ASAP7_75t_L g7633 ( 
.A(n_7353),
.B(n_6990),
.C(n_6993),
.D(n_6986),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7313),
.Y(n_7634)
);

NAND3xp33_ASAP7_75t_SL g7635 ( 
.A(n_7437),
.B(n_7094),
.C(n_7064),
.Y(n_7635)
);

HB1xp67_ASAP7_75t_L g7636 ( 
.A(n_7263),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7323),
.Y(n_7637)
);

NOR2x1_ASAP7_75t_SL g7638 ( 
.A(n_7448),
.B(n_5401),
.Y(n_7638)
);

NAND3xp33_ASAP7_75t_L g7639 ( 
.A(n_7272),
.B(n_6995),
.C(n_6994),
.Y(n_7639)
);

AND2x2_ASAP7_75t_L g7640 ( 
.A(n_7167),
.B(n_7056),
.Y(n_7640)
);

INVx1_ASAP7_75t_L g7641 ( 
.A(n_7323),
.Y(n_7641)
);

INVx2_ASAP7_75t_L g7642 ( 
.A(n_7304),
.Y(n_7642)
);

NAND3xp33_ASAP7_75t_L g7643 ( 
.A(n_7365),
.B(n_7009),
.C(n_7005),
.Y(n_7643)
);

NAND3xp33_ASAP7_75t_L g7644 ( 
.A(n_7448),
.B(n_7028),
.C(n_7023),
.Y(n_7644)
);

NAND2xp5_ASAP7_75t_L g7645 ( 
.A(n_7182),
.B(n_7032),
.Y(n_7645)
);

AND2x4_ASAP7_75t_L g7646 ( 
.A(n_7165),
.B(n_7044),
.Y(n_7646)
);

AND2x2_ASAP7_75t_L g7647 ( 
.A(n_7187),
.B(n_7100),
.Y(n_7647)
);

NAND2xp5_ASAP7_75t_L g7648 ( 
.A(n_7190),
.B(n_7035),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7335),
.Y(n_7649)
);

NOR3xp33_ASAP7_75t_SL g7650 ( 
.A(n_7386),
.B(n_7043),
.C(n_7039),
.Y(n_7650)
);

AOI22xp5_ASAP7_75t_L g7651 ( 
.A1(n_7327),
.A2(n_7053),
.B1(n_7049),
.B2(n_5982),
.Y(n_7651)
);

NOR3xp33_ASAP7_75t_L g7652 ( 
.A(n_7445),
.B(n_6992),
.C(n_6949),
.Y(n_7652)
);

NAND3xp33_ASAP7_75t_L g7653 ( 
.A(n_7457),
.B(n_7017),
.C(n_6999),
.Y(n_7653)
);

NOR3xp33_ASAP7_75t_L g7654 ( 
.A(n_7445),
.B(n_7017),
.C(n_6999),
.Y(n_7654)
);

OAI22xp5_ASAP7_75t_L g7655 ( 
.A1(n_7468),
.A2(n_7477),
.B1(n_7461),
.B2(n_7464),
.Y(n_7655)
);

NAND4xp75_ASAP7_75t_L g7656 ( 
.A(n_7366),
.B(n_6500),
.C(n_6499),
.D(n_6683),
.Y(n_7656)
);

NAND3xp33_ASAP7_75t_L g7657 ( 
.A(n_7457),
.B(n_7029),
.C(n_7020),
.Y(n_7657)
);

AND2x2_ASAP7_75t_L g7658 ( 
.A(n_7452),
.B(n_7304),
.Y(n_7658)
);

INVx1_ASAP7_75t_SL g7659 ( 
.A(n_7301),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7335),
.Y(n_7660)
);

NAND3xp33_ASAP7_75t_L g7661 ( 
.A(n_7457),
.B(n_7029),
.C(n_7020),
.Y(n_7661)
);

NOR3xp33_ASAP7_75t_L g7662 ( 
.A(n_7351),
.B(n_7091),
.C(n_7082),
.Y(n_7662)
);

NAND3xp33_ASAP7_75t_SL g7663 ( 
.A(n_7357),
.B(n_7112),
.C(n_7093),
.Y(n_7663)
);

HB1xp67_ASAP7_75t_L g7664 ( 
.A(n_7132),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7159),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7382),
.Y(n_7666)
);

NAND3xp33_ASAP7_75t_L g7667 ( 
.A(n_7470),
.B(n_7093),
.C(n_7091),
.Y(n_7667)
);

NOR2x1_ASAP7_75t_L g7668 ( 
.A(n_7374),
.B(n_4936),
.Y(n_7668)
);

AND2x2_ASAP7_75t_L g7669 ( 
.A(n_7401),
.B(n_7102),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_7382),
.Y(n_7670)
);

OR2x2_ASAP7_75t_L g7671 ( 
.A(n_7359),
.B(n_6160),
.Y(n_7671)
);

AND2x2_ASAP7_75t_L g7672 ( 
.A(n_7436),
.B(n_5707),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7387),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_7387),
.Y(n_7674)
);

OAI211xp5_ASAP7_75t_L g7675 ( 
.A1(n_7291),
.A2(n_5301),
.B(n_5415),
.C(n_5402),
.Y(n_7675)
);

NAND4xp75_ASAP7_75t_L g7676 ( 
.A(n_7420),
.B(n_6500),
.C(n_6686),
.D(n_6683),
.Y(n_7676)
);

NAND3xp33_ASAP7_75t_L g7677 ( 
.A(n_7199),
.B(n_5992),
.C(n_5988),
.Y(n_7677)
);

NAND2xp5_ASAP7_75t_L g7678 ( 
.A(n_7146),
.B(n_5912),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7155),
.B(n_6208),
.Y(n_7679)
);

NAND3xp33_ASAP7_75t_L g7680 ( 
.A(n_7337),
.B(n_7352),
.C(n_7339),
.Y(n_7680)
);

INVx2_ASAP7_75t_L g7681 ( 
.A(n_7225),
.Y(n_7681)
);

NAND2xp5_ASAP7_75t_L g7682 ( 
.A(n_7225),
.B(n_6209),
.Y(n_7682)
);

NAND3xp33_ASAP7_75t_L g7683 ( 
.A(n_7274),
.B(n_7264),
.C(n_7254),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_7156),
.B(n_6213),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7450),
.Y(n_7685)
);

AND2x4_ASAP7_75t_L g7686 ( 
.A(n_7456),
.B(n_4780),
.Y(n_7686)
);

AND2x2_ASAP7_75t_L g7687 ( 
.A(n_7360),
.B(n_5707),
.Y(n_7687)
);

AND2x2_ASAP7_75t_L g7688 ( 
.A(n_7363),
.B(n_5707),
.Y(n_7688)
);

HB1xp67_ASAP7_75t_L g7689 ( 
.A(n_7191),
.Y(n_7689)
);

AO21x2_ASAP7_75t_L g7690 ( 
.A1(n_7194),
.A2(n_6392),
.B(n_6391),
.Y(n_7690)
);

NAND2xp5_ASAP7_75t_L g7691 ( 
.A(n_7340),
.B(n_6216),
.Y(n_7691)
);

NAND3xp33_ASAP7_75t_L g7692 ( 
.A(n_7362),
.B(n_5992),
.C(n_6391),
.Y(n_7692)
);

NOR4xp25_ASAP7_75t_L g7693 ( 
.A(n_7298),
.B(n_6398),
.C(n_6399),
.D(n_6392),
.Y(n_7693)
);

AND2x2_ASAP7_75t_L g7694 ( 
.A(n_7234),
.B(n_5638),
.Y(n_7694)
);

AND2x2_ASAP7_75t_L g7695 ( 
.A(n_7454),
.B(n_5062),
.Y(n_7695)
);

INVx1_ASAP7_75t_SL g7696 ( 
.A(n_7456),
.Y(n_7696)
);

OR2x2_ASAP7_75t_L g7697 ( 
.A(n_7443),
.B(n_5952),
.Y(n_7697)
);

OR2x2_ASAP7_75t_L g7698 ( 
.A(n_7447),
.B(n_5952),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7450),
.Y(n_7699)
);

NAND3xp33_ASAP7_75t_L g7700 ( 
.A(n_7262),
.B(n_6410),
.C(n_6399),
.Y(n_7700)
);

AOI22xp33_ASAP7_75t_L g7701 ( 
.A1(n_7302),
.A2(n_6695),
.B1(n_6696),
.B2(n_6686),
.Y(n_7701)
);

NOR2x1_ASAP7_75t_SL g7702 ( 
.A(n_7221),
.B(n_5401),
.Y(n_7702)
);

NOR2x1_ASAP7_75t_R g7703 ( 
.A(n_7161),
.B(n_4936),
.Y(n_7703)
);

NAND4xp75_ASAP7_75t_L g7704 ( 
.A(n_7223),
.B(n_6696),
.C(n_6695),
.D(n_6405),
.Y(n_7704)
);

NAND3xp33_ASAP7_75t_L g7705 ( 
.A(n_7256),
.B(n_6405),
.C(n_6398),
.Y(n_7705)
);

OAI21xp5_ASAP7_75t_L g7706 ( 
.A1(n_7138),
.A2(n_5841),
.B(n_5820),
.Y(n_7706)
);

NOR3xp33_ASAP7_75t_SL g7707 ( 
.A(n_7334),
.B(n_5081),
.C(n_5078),
.Y(n_7707)
);

INVx2_ASAP7_75t_SL g7708 ( 
.A(n_7425),
.Y(n_7708)
);

OR2x2_ASAP7_75t_L g7709 ( 
.A(n_7453),
.B(n_6227),
.Y(n_7709)
);

AND2x2_ASAP7_75t_L g7710 ( 
.A(n_7458),
.B(n_5458),
.Y(n_7710)
);

INVxp67_ASAP7_75t_L g7711 ( 
.A(n_7399),
.Y(n_7711)
);

NAND2xp5_ASAP7_75t_SL g7712 ( 
.A(n_7325),
.B(n_7239),
.Y(n_7712)
);

AND2x2_ASAP7_75t_L g7713 ( 
.A(n_7480),
.B(n_5458),
.Y(n_7713)
);

AOI22xp33_ASAP7_75t_SL g7714 ( 
.A1(n_7307),
.A2(n_5402),
.B1(n_5468),
.B2(n_5436),
.Y(n_7714)
);

AND2x2_ASAP7_75t_L g7715 ( 
.A(n_7368),
.B(n_5473),
.Y(n_7715)
);

XNOR2xp5_ASAP7_75t_L g7716 ( 
.A(n_7176),
.B(n_4445),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7465),
.Y(n_7717)
);

NAND2xp5_ASAP7_75t_L g7718 ( 
.A(n_7259),
.B(n_7271),
.Y(n_7718)
);

NAND4xp75_ASAP7_75t_L g7719 ( 
.A(n_7247),
.B(n_6410),
.C(n_6412),
.D(n_6406),
.Y(n_7719)
);

OR2x2_ASAP7_75t_L g7720 ( 
.A(n_7481),
.B(n_6227),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_7465),
.Y(n_7721)
);

NAND2xp5_ASAP7_75t_L g7722 ( 
.A(n_7394),
.B(n_6251),
.Y(n_7722)
);

AND2x2_ASAP7_75t_L g7723 ( 
.A(n_7373),
.B(n_5473),
.Y(n_7723)
);

AND2x2_ASAP7_75t_L g7724 ( 
.A(n_7379),
.B(n_5479),
.Y(n_7724)
);

NOR2xp33_ASAP7_75t_L g7725 ( 
.A(n_7374),
.B(n_5093),
.Y(n_7725)
);

OR2x2_ASAP7_75t_L g7726 ( 
.A(n_7358),
.B(n_6217),
.Y(n_7726)
);

INVxp67_ASAP7_75t_L g7727 ( 
.A(n_7239),
.Y(n_7727)
);

AND2x2_ASAP7_75t_L g7728 ( 
.A(n_7405),
.B(n_5479),
.Y(n_7728)
);

OR2x2_ASAP7_75t_L g7729 ( 
.A(n_7212),
.B(n_6237),
.Y(n_7729)
);

AND2x2_ASAP7_75t_L g7730 ( 
.A(n_7414),
.B(n_5551),
.Y(n_7730)
);

NAND4xp75_ASAP7_75t_L g7731 ( 
.A(n_7258),
.B(n_6412),
.C(n_6418),
.D(n_6406),
.Y(n_7731)
);

NAND2xp5_ASAP7_75t_L g7732 ( 
.A(n_7197),
.B(n_6220),
.Y(n_7732)
);

AND2x2_ASAP7_75t_L g7733 ( 
.A(n_7432),
.B(n_5551),
.Y(n_7733)
);

NAND2xp5_ASAP7_75t_SL g7734 ( 
.A(n_7325),
.B(n_5618),
.Y(n_7734)
);

NAND2xp5_ASAP7_75t_L g7735 ( 
.A(n_7211),
.B(n_6228),
.Y(n_7735)
);

AND2x2_ASAP7_75t_L g7736 ( 
.A(n_7260),
.B(n_5523),
.Y(n_7736)
);

AOI22xp33_ASAP7_75t_L g7737 ( 
.A1(n_7308),
.A2(n_6418),
.B1(n_6609),
.B2(n_6597),
.Y(n_7737)
);

OAI22xp33_ASAP7_75t_L g7738 ( 
.A1(n_7451),
.A2(n_5476),
.B1(n_7333),
.B2(n_7336),
.Y(n_7738)
);

OAI211xp5_ASAP7_75t_L g7739 ( 
.A1(n_7221),
.A2(n_5436),
.B(n_5478),
.C(n_5468),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_7408),
.Y(n_7740)
);

OR2x2_ASAP7_75t_L g7741 ( 
.A(n_7378),
.B(n_6230),
.Y(n_7741)
);

NAND2x1p5_ASAP7_75t_L g7742 ( 
.A(n_7221),
.B(n_5105),
.Y(n_7742)
);

NAND3xp33_ASAP7_75t_SL g7743 ( 
.A(n_7372),
.B(n_5704),
.C(n_5556),
.Y(n_7743)
);

NAND3xp33_ASAP7_75t_L g7744 ( 
.A(n_7210),
.B(n_6609),
.C(n_6597),
.Y(n_7744)
);

HB1xp67_ASAP7_75t_L g7745 ( 
.A(n_7331),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_L g7746 ( 
.A(n_7214),
.B(n_6241),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7408),
.Y(n_7747)
);

NOR3xp33_ASAP7_75t_SL g7748 ( 
.A(n_7311),
.B(n_4496),
.C(n_4685),
.Y(n_7748)
);

OR2x2_ASAP7_75t_L g7749 ( 
.A(n_7428),
.B(n_6245),
.Y(n_7749)
);

NOR3xp33_ASAP7_75t_L g7750 ( 
.A(n_7431),
.B(n_6610),
.C(n_5819),
.Y(n_7750)
);

NAND4xp75_ASAP7_75t_L g7751 ( 
.A(n_7442),
.B(n_6610),
.C(n_5777),
.D(n_5778),
.Y(n_7751)
);

NAND4xp75_ASAP7_75t_L g7752 ( 
.A(n_7232),
.B(n_5777),
.C(n_5778),
.D(n_5773),
.Y(n_7752)
);

NAND2xp5_ASAP7_75t_SL g7753 ( 
.A(n_7200),
.B(n_5618),
.Y(n_7753)
);

AND2x2_ASAP7_75t_L g7754 ( 
.A(n_7260),
.B(n_5523),
.Y(n_7754)
);

NAND3xp33_ASAP7_75t_L g7755 ( 
.A(n_7236),
.B(n_5819),
.C(n_5812),
.Y(n_7755)
);

OAI22xp5_ASAP7_75t_L g7756 ( 
.A1(n_7415),
.A2(n_5633),
.B1(n_5704),
.B2(n_5556),
.Y(n_7756)
);

AND2x2_ASAP7_75t_L g7757 ( 
.A(n_7415),
.B(n_5239),
.Y(n_7757)
);

AND2x2_ASAP7_75t_L g7758 ( 
.A(n_7384),
.B(n_5268),
.Y(n_7758)
);

AND2x2_ASAP7_75t_L g7759 ( 
.A(n_7375),
.B(n_5268),
.Y(n_7759)
);

AND2x2_ASAP7_75t_L g7760 ( 
.A(n_7356),
.B(n_5676),
.Y(n_7760)
);

NAND3xp33_ASAP7_75t_L g7761 ( 
.A(n_7249),
.B(n_5826),
.C(n_5812),
.Y(n_7761)
);

OR2x2_ASAP7_75t_L g7762 ( 
.A(n_7163),
.B(n_6246),
.Y(n_7762)
);

NAND2xp5_ASAP7_75t_L g7763 ( 
.A(n_7404),
.B(n_7406),
.Y(n_7763)
);

NAND4xp75_ASAP7_75t_L g7764 ( 
.A(n_7201),
.B(n_5780),
.C(n_5789),
.D(n_5773),
.Y(n_7764)
);

OR2x2_ASAP7_75t_L g7765 ( 
.A(n_7170),
.B(n_7315),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7410),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_L g7767 ( 
.A(n_7407),
.B(n_6258),
.Y(n_7767)
);

NOR2xp33_ASAP7_75t_L g7768 ( 
.A(n_7161),
.B(n_5093),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_7410),
.Y(n_7769)
);

AND2x2_ASAP7_75t_L g7770 ( 
.A(n_7367),
.B(n_7130),
.Y(n_7770)
);

NOR3xp33_ASAP7_75t_L g7771 ( 
.A(n_7204),
.B(n_5827),
.C(n_5826),
.Y(n_7771)
);

INVx2_ASAP7_75t_L g7772 ( 
.A(n_7189),
.Y(n_7772)
);

NAND3xp33_ASAP7_75t_L g7773 ( 
.A(n_7205),
.B(n_5468),
.C(n_5436),
.Y(n_7773)
);

OR2x2_ASAP7_75t_SL g7774 ( 
.A(n_7269),
.B(n_4465),
.Y(n_7774)
);

NOR3xp33_ASAP7_75t_L g7775 ( 
.A(n_7338),
.B(n_5833),
.C(n_5827),
.Y(n_7775)
);

AOI211xp5_ASAP7_75t_L g7776 ( 
.A1(n_7298),
.A2(n_7300),
.B(n_7299),
.C(n_7413),
.Y(n_7776)
);

AND2x2_ASAP7_75t_L g7777 ( 
.A(n_7130),
.B(n_5676),
.Y(n_7777)
);

AND2x2_ASAP7_75t_L g7778 ( 
.A(n_7209),
.B(n_5687),
.Y(n_7778)
);

NAND4xp75_ASAP7_75t_L g7779 ( 
.A(n_7208),
.B(n_5789),
.C(n_5792),
.D(n_5780),
.Y(n_7779)
);

AND2x2_ASAP7_75t_L g7780 ( 
.A(n_7209),
.B(n_5687),
.Y(n_7780)
);

NOR2xp33_ASAP7_75t_L g7781 ( 
.A(n_7164),
.B(n_7305),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7421),
.Y(n_7782)
);

OR2x2_ASAP7_75t_L g7783 ( 
.A(n_7316),
.B(n_5994),
.Y(n_7783)
);

OR2x2_ASAP7_75t_L g7784 ( 
.A(n_7157),
.B(n_5994),
.Y(n_7784)
);

AND2x2_ASAP7_75t_L g7785 ( 
.A(n_7241),
.B(n_5269),
.Y(n_7785)
);

NOR2x1_ASAP7_75t_L g7786 ( 
.A(n_7164),
.B(n_5478),
.Y(n_7786)
);

INVx2_ASAP7_75t_SL g7787 ( 
.A(n_7441),
.Y(n_7787)
);

AOI22xp33_ASAP7_75t_L g7788 ( 
.A1(n_7308),
.A2(n_6623),
.B1(n_5802),
.B2(n_5808),
.Y(n_7788)
);

OA211x2_ASAP7_75t_L g7789 ( 
.A1(n_7282),
.A2(n_3898),
.B(n_5618),
.C(n_4354),
.Y(n_7789)
);

NOR2xp33_ASAP7_75t_L g7790 ( 
.A(n_7329),
.B(n_5093),
.Y(n_7790)
);

AOI22xp33_ASAP7_75t_L g7791 ( 
.A1(n_7319),
.A2(n_6623),
.B1(n_5802),
.B2(n_5808),
.Y(n_7791)
);

INVx2_ASAP7_75t_L g7792 ( 
.A(n_7219),
.Y(n_7792)
);

NAND3xp33_ASAP7_75t_L g7793 ( 
.A(n_7213),
.B(n_5494),
.C(n_5478),
.Y(n_7793)
);

AO21x2_ASAP7_75t_L g7794 ( 
.A1(n_7217),
.A2(n_5792),
.B(n_5833),
.Y(n_7794)
);

AND2x2_ASAP7_75t_L g7795 ( 
.A(n_7241),
.B(n_5269),
.Y(n_7795)
);

AO21x2_ASAP7_75t_L g7796 ( 
.A1(n_7218),
.A2(n_5849),
.B(n_5846),
.Y(n_7796)
);

OR2x2_ASAP7_75t_L g7797 ( 
.A(n_7416),
.B(n_5999),
.Y(n_7797)
);

AOI22xp33_ASAP7_75t_L g7798 ( 
.A1(n_7319),
.A2(n_5849),
.B1(n_5855),
.B2(n_5846),
.Y(n_7798)
);

BUFx2_ASAP7_75t_L g7799 ( 
.A(n_7537),
.Y(n_7799)
);

AO31x2_ASAP7_75t_L g7800 ( 
.A1(n_7740),
.A2(n_7229),
.A3(n_7231),
.B(n_7227),
.Y(n_7800)
);

AND2x2_ASAP7_75t_L g7801 ( 
.A(n_7485),
.B(n_7475),
.Y(n_7801)
);

AND2x2_ASAP7_75t_L g7802 ( 
.A(n_7529),
.B(n_7530),
.Y(n_7802)
);

OR2x2_ASAP7_75t_L g7803 ( 
.A(n_7523),
.B(n_7417),
.Y(n_7803)
);

INVx4_ASAP7_75t_L g7804 ( 
.A(n_7547),
.Y(n_7804)
);

AND2x2_ASAP7_75t_L g7805 ( 
.A(n_7534),
.B(n_7459),
.Y(n_7805)
);

OR2x2_ASAP7_75t_L g7806 ( 
.A(n_7508),
.B(n_7418),
.Y(n_7806)
);

NOR3xp33_ASAP7_75t_SL g7807 ( 
.A(n_7620),
.B(n_7278),
.C(n_7355),
.Y(n_7807)
);

OAI21xp5_ASAP7_75t_L g7808 ( 
.A1(n_7680),
.A2(n_7257),
.B(n_7446),
.Y(n_7808)
);

AND2x2_ASAP7_75t_L g7809 ( 
.A(n_7632),
.B(n_7460),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7493),
.Y(n_7810)
);

OR2x2_ASAP7_75t_L g7811 ( 
.A(n_7543),
.B(n_7423),
.Y(n_7811)
);

INVx4_ASAP7_75t_L g7812 ( 
.A(n_7489),
.Y(n_7812)
);

AND2x2_ASAP7_75t_L g7813 ( 
.A(n_7505),
.B(n_7462),
.Y(n_7813)
);

NAND3xp33_ASAP7_75t_SL g7814 ( 
.A(n_7502),
.B(n_7300),
.C(n_7299),
.Y(n_7814)
);

NAND2x1p5_ASAP7_75t_L g7815 ( 
.A(n_7696),
.B(n_7600),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_7520),
.Y(n_7816)
);

NOR3xp33_ASAP7_75t_L g7817 ( 
.A(n_7506),
.B(n_7252),
.C(n_7246),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7520),
.Y(n_7818)
);

NAND2xp5_ASAP7_75t_L g7819 ( 
.A(n_7636),
.B(n_7426),
.Y(n_7819)
);

AOI22xp33_ASAP7_75t_L g7820 ( 
.A1(n_7750),
.A2(n_7610),
.B1(n_7612),
.B2(n_7608),
.Y(n_7820)
);

NOR2x1p5_ASAP7_75t_L g7821 ( 
.A(n_7578),
.B(n_7592),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_7527),
.Y(n_7822)
);

AOI33xp33_ASAP7_75t_L g7823 ( 
.A1(n_7502),
.A2(n_7455),
.A3(n_7438),
.B1(n_7469),
.B2(n_7439),
.B3(n_7427),
.Y(n_7823)
);

AND2x2_ASAP7_75t_L g7824 ( 
.A(n_7532),
.B(n_7398),
.Y(n_7824)
);

BUFx2_ASAP7_75t_L g7825 ( 
.A(n_7509),
.Y(n_7825)
);

AND2x2_ASAP7_75t_L g7826 ( 
.A(n_7490),
.B(n_7419),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7527),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_7541),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_7539),
.B(n_7342),
.Y(n_7829)
);

BUFx2_ASAP7_75t_L g7830 ( 
.A(n_7509),
.Y(n_7830)
);

INVx2_ASAP7_75t_L g7831 ( 
.A(n_7540),
.Y(n_7831)
);

NOR2xp33_ASAP7_75t_L g7832 ( 
.A(n_7588),
.B(n_7540),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7747),
.Y(n_7833)
);

INVx1_ASAP7_75t_SL g7834 ( 
.A(n_7487),
.Y(n_7834)
);

HB1xp67_ASAP7_75t_L g7835 ( 
.A(n_7553),
.Y(n_7835)
);

AND2x2_ASAP7_75t_L g7836 ( 
.A(n_7566),
.B(n_7580),
.Y(n_7836)
);

NAND2xp5_ASAP7_75t_L g7837 ( 
.A(n_7647),
.B(n_7342),
.Y(n_7837)
);

INVx4_ASAP7_75t_L g7838 ( 
.A(n_7686),
.Y(n_7838)
);

AND2x2_ASAP7_75t_L g7839 ( 
.A(n_7669),
.B(n_7429),
.Y(n_7839)
);

NAND2xp5_ASAP7_75t_L g7840 ( 
.A(n_7745),
.B(n_7343),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_7766),
.Y(n_7841)
);

AOI222xp33_ASAP7_75t_L g7842 ( 
.A1(n_7769),
.A2(n_7321),
.B1(n_7332),
.B2(n_7324),
.C1(n_7370),
.C2(n_7364),
.Y(n_7842)
);

AND2x2_ASAP7_75t_L g7843 ( 
.A(n_7556),
.B(n_7449),
.Y(n_7843)
);

OAI31xp33_ASAP7_75t_L g7844 ( 
.A1(n_7501),
.A2(n_7346),
.A3(n_7471),
.B(n_7376),
.Y(n_7844)
);

OR2x2_ASAP7_75t_L g7845 ( 
.A(n_7497),
.B(n_7343),
.Y(n_7845)
);

HB1xp67_ASAP7_75t_L g7846 ( 
.A(n_7553),
.Y(n_7846)
);

OAI21xp5_ASAP7_75t_L g7847 ( 
.A1(n_7498),
.A2(n_7281),
.B(n_7412),
.Y(n_7847)
);

AND2x2_ASAP7_75t_L g7848 ( 
.A(n_7503),
.B(n_7504),
.Y(n_7848)
);

AO21x2_ASAP7_75t_L g7849 ( 
.A1(n_7782),
.A2(n_7369),
.B(n_7327),
.Y(n_7849)
);

NAND4xp25_ASAP7_75t_L g7850 ( 
.A(n_7484),
.B(n_7354),
.C(n_7474),
.D(n_7472),
.Y(n_7850)
);

AND2x2_ASAP7_75t_L g7851 ( 
.A(n_7528),
.B(n_7354),
.Y(n_7851)
);

AND2x2_ASAP7_75t_SL g7852 ( 
.A(n_7686),
.B(n_7328),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7565),
.Y(n_7853)
);

AND2x2_ASAP7_75t_L g7854 ( 
.A(n_7604),
.B(n_7472),
.Y(n_7854)
);

NAND2xp5_ASAP7_75t_SL g7855 ( 
.A(n_7611),
.B(n_7474),
.Y(n_7855)
);

AND2x4_ASAP7_75t_L g7856 ( 
.A(n_7626),
.B(n_7476),
.Y(n_7856)
);

NAND2xp5_ASAP7_75t_L g7857 ( 
.A(n_7689),
.B(n_7713),
.Y(n_7857)
);

AND2x2_ASAP7_75t_L g7858 ( 
.A(n_7587),
.B(n_7476),
.Y(n_7858)
);

NAND2xp5_ASAP7_75t_L g7859 ( 
.A(n_7715),
.B(n_7723),
.Y(n_7859)
);

BUFx3_ASAP7_75t_L g7860 ( 
.A(n_7681),
.Y(n_7860)
);

AND2x2_ASAP7_75t_L g7861 ( 
.A(n_7631),
.B(n_7478),
.Y(n_7861)
);

OAI33xp33_ASAP7_75t_L g7862 ( 
.A1(n_7495),
.A2(n_7483),
.A3(n_7479),
.B1(n_7482),
.B2(n_7478),
.B3(n_7390),
.Y(n_7862)
);

NAND2xp5_ASAP7_75t_L g7863 ( 
.A(n_7724),
.B(n_7482),
.Y(n_7863)
);

INVx1_ASAP7_75t_SL g7864 ( 
.A(n_7526),
.Y(n_7864)
);

AND2x4_ASAP7_75t_L g7865 ( 
.A(n_7611),
.B(n_7479),
.Y(n_7865)
);

NAND3xp33_ASAP7_75t_L g7866 ( 
.A(n_7510),
.B(n_7483),
.C(n_7383),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7565),
.Y(n_7867)
);

NAND2xp5_ASAP7_75t_L g7868 ( 
.A(n_7728),
.B(n_7369),
.Y(n_7868)
);

AND2x2_ASAP7_75t_L g7869 ( 
.A(n_7630),
.B(n_7238),
.Y(n_7869)
);

INVx2_ASAP7_75t_L g7870 ( 
.A(n_7589),
.Y(n_7870)
);

BUFx2_ASAP7_75t_L g7871 ( 
.A(n_7646),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_7582),
.Y(n_7872)
);

OAI31xp33_ASAP7_75t_SL g7873 ( 
.A1(n_7498),
.A2(n_7409),
.A3(n_7350),
.B(n_7326),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7582),
.Y(n_7874)
);

OR2x2_ASAP7_75t_L g7875 ( 
.A(n_7571),
.B(n_7307),
.Y(n_7875)
);

INVx1_ASAP7_75t_L g7876 ( 
.A(n_7542),
.Y(n_7876)
);

BUFx3_ASAP7_75t_L g7877 ( 
.A(n_7658),
.Y(n_7877)
);

OR2x2_ASAP7_75t_L g7878 ( 
.A(n_7627),
.B(n_7421),
.Y(n_7878)
);

AOI33xp33_ASAP7_75t_L g7879 ( 
.A1(n_7577),
.A2(n_7510),
.A3(n_7558),
.B1(n_7659),
.B2(n_7512),
.B3(n_7776),
.Y(n_7879)
);

OR2x2_ASAP7_75t_L g7880 ( 
.A(n_7628),
.B(n_7473),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7634),
.Y(n_7881)
);

AOI22xp33_ASAP7_75t_L g7882 ( 
.A1(n_7637),
.A2(n_7324),
.B1(n_7332),
.B2(n_7321),
.Y(n_7882)
);

OAI33xp33_ASAP7_75t_L g7883 ( 
.A1(n_7496),
.A2(n_7400),
.A3(n_7385),
.B1(n_7402),
.B2(n_7391),
.B3(n_7371),
.Y(n_7883)
);

OAI221xp5_ASAP7_75t_L g7884 ( 
.A1(n_7651),
.A2(n_7411),
.B1(n_7403),
.B2(n_7171),
.C(n_7151),
.Y(n_7884)
);

INVx1_ASAP7_75t_L g7885 ( 
.A(n_7641),
.Y(n_7885)
);

INVx1_ASAP7_75t_L g7886 ( 
.A(n_7649),
.Y(n_7886)
);

INVx2_ASAP7_75t_L g7887 ( 
.A(n_7589),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_7660),
.Y(n_7888)
);

OR2x2_ASAP7_75t_L g7889 ( 
.A(n_7671),
.B(n_6000),
.Y(n_7889)
);

OR2x2_ASAP7_75t_L g7890 ( 
.A(n_7555),
.B(n_6000),
.Y(n_7890)
);

AND2x2_ASAP7_75t_L g7891 ( 
.A(n_7590),
.B(n_5269),
.Y(n_7891)
);

OR2x2_ASAP7_75t_L g7892 ( 
.A(n_7596),
.B(n_6036),
.Y(n_7892)
);

HB1xp67_ASAP7_75t_L g7893 ( 
.A(n_7642),
.Y(n_7893)
);

INVx2_ASAP7_75t_L g7894 ( 
.A(n_7794),
.Y(n_7894)
);

INVx1_ASAP7_75t_L g7895 ( 
.A(n_7666),
.Y(n_7895)
);

AND2x4_ASAP7_75t_L g7896 ( 
.A(n_7519),
.B(n_7646),
.Y(n_7896)
);

AND2x2_ASAP7_75t_L g7897 ( 
.A(n_7777),
.B(n_7778),
.Y(n_7897)
);

NOR3xp33_ASAP7_75t_L g7898 ( 
.A(n_7711),
.B(n_7496),
.C(n_7518),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_7670),
.Y(n_7899)
);

OR2x2_ASAP7_75t_L g7900 ( 
.A(n_7709),
.B(n_6036),
.Y(n_7900)
);

NAND2xp5_ASAP7_75t_L g7901 ( 
.A(n_7730),
.B(n_7185),
.Y(n_7901)
);

NAND2xp5_ASAP7_75t_L g7902 ( 
.A(n_7733),
.B(n_7694),
.Y(n_7902)
);

NAND4xp25_ASAP7_75t_L g7903 ( 
.A(n_7484),
.B(n_5105),
.C(n_5047),
.D(n_4387),
.Y(n_7903)
);

AND2x2_ASAP7_75t_L g7904 ( 
.A(n_7780),
.B(n_5269),
.Y(n_7904)
);

AND4x1_ASAP7_75t_L g7905 ( 
.A(n_7488),
.B(n_5096),
.C(n_4691),
.D(n_4858),
.Y(n_7905)
);

AOI22xp33_ASAP7_75t_SL g7906 ( 
.A1(n_7638),
.A2(n_7151),
.B1(n_7171),
.B2(n_7144),
.Y(n_7906)
);

HB1xp67_ASAP7_75t_L g7907 ( 
.A(n_7727),
.Y(n_7907)
);

OR2x2_ASAP7_75t_L g7908 ( 
.A(n_7698),
.B(n_6012),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_7673),
.Y(n_7909)
);

AND2x2_ASAP7_75t_L g7910 ( 
.A(n_7708),
.B(n_5269),
.Y(n_7910)
);

OR2x2_ASAP7_75t_L g7911 ( 
.A(n_7499),
.B(n_6012),
.Y(n_7911)
);

INVx1_ASAP7_75t_L g7912 ( 
.A(n_7674),
.Y(n_7912)
);

INVx2_ASAP7_75t_L g7913 ( 
.A(n_7794),
.Y(n_7913)
);

INVx1_ASAP7_75t_SL g7914 ( 
.A(n_7770),
.Y(n_7914)
);

INVx2_ASAP7_75t_L g7915 ( 
.A(n_7796),
.Y(n_7915)
);

INVx1_ASAP7_75t_L g7916 ( 
.A(n_7685),
.Y(n_7916)
);

AO21x2_ASAP7_75t_L g7917 ( 
.A1(n_7699),
.A2(n_7185),
.B(n_7144),
.Y(n_7917)
);

AND2x2_ASAP7_75t_L g7918 ( 
.A(n_7607),
.B(n_5269),
.Y(n_7918)
);

AOI211xp5_ASAP7_75t_SL g7919 ( 
.A1(n_7552),
.A2(n_5494),
.B(n_5530),
.C(n_5478),
.Y(n_7919)
);

OAI33xp33_ASAP7_75t_L g7920 ( 
.A1(n_7501),
.A2(n_5869),
.A3(n_5861),
.B1(n_5884),
.B2(n_5866),
.B3(n_5855),
.Y(n_7920)
);

AND2x2_ASAP7_75t_L g7921 ( 
.A(n_7622),
.B(n_5269),
.Y(n_7921)
);

INVx3_ASAP7_75t_L g7922 ( 
.A(n_7796),
.Y(n_7922)
);

BUFx3_ASAP7_75t_L g7923 ( 
.A(n_7538),
.Y(n_7923)
);

AND2x4_ASAP7_75t_L g7924 ( 
.A(n_7640),
.B(n_5679),
.Y(n_7924)
);

INVx2_ASAP7_75t_L g7925 ( 
.A(n_7774),
.Y(n_7925)
);

AOI211xp5_ASAP7_75t_L g7926 ( 
.A1(n_7492),
.A2(n_5494),
.B(n_5573),
.C(n_5530),
.Y(n_7926)
);

NAND4xp25_ASAP7_75t_L g7927 ( 
.A(n_7619),
.B(n_5105),
.C(n_5047),
.D(n_4387),
.Y(n_7927)
);

NOR2x1_ASAP7_75t_L g7928 ( 
.A(n_7574),
.B(n_7605),
.Y(n_7928)
);

NAND2xp5_ASAP7_75t_L g7929 ( 
.A(n_7710),
.B(n_5999),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_L g7930 ( 
.A(n_7664),
.B(n_6020),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7717),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7721),
.Y(n_7932)
);

INVx4_ASAP7_75t_L g7933 ( 
.A(n_7516),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_7651),
.Y(n_7934)
);

AOI22xp5_ASAP7_75t_L g7935 ( 
.A1(n_7751),
.A2(n_5866),
.B1(n_5869),
.B2(n_5861),
.Y(n_7935)
);

OAI21xp5_ASAP7_75t_L g7936 ( 
.A1(n_7517),
.A2(n_5841),
.B(n_5820),
.Y(n_7936)
);

INVx2_ASAP7_75t_L g7937 ( 
.A(n_7617),
.Y(n_7937)
);

HB1xp67_ASAP7_75t_L g7938 ( 
.A(n_7531),
.Y(n_7938)
);

INVx3_ASAP7_75t_L g7939 ( 
.A(n_7500),
.Y(n_7939)
);

AND2x2_ASAP7_75t_L g7940 ( 
.A(n_7606),
.B(n_5269),
.Y(n_7940)
);

AND2x4_ASAP7_75t_L g7941 ( 
.A(n_7515),
.B(n_5679),
.Y(n_7941)
);

AND2x4_ASAP7_75t_L g7942 ( 
.A(n_7525),
.B(n_5679),
.Y(n_7942)
);

AND2x2_ASAP7_75t_L g7943 ( 
.A(n_7569),
.B(n_5269),
.Y(n_7943)
);

INVx2_ASAP7_75t_SL g7944 ( 
.A(n_7544),
.Y(n_7944)
);

NAND2xp5_ASAP7_75t_L g7945 ( 
.A(n_7662),
.B(n_6020),
.Y(n_7945)
);

NAND2xp5_ASAP7_75t_L g7946 ( 
.A(n_7593),
.B(n_6021),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7683),
.Y(n_7947)
);

OR2x2_ASAP7_75t_L g7948 ( 
.A(n_7765),
.B(n_6058),
.Y(n_7948)
);

NAND2xp5_ASAP7_75t_L g7949 ( 
.A(n_7652),
.B(n_6021),
.Y(n_7949)
);

HB1xp67_ASAP7_75t_L g7950 ( 
.A(n_7486),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7690),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7690),
.Y(n_7952)
);

OAI221xp5_ASAP7_75t_L g7953 ( 
.A1(n_7512),
.A2(n_5573),
.B1(n_5530),
.B2(n_5494),
.C(n_5884),
.Y(n_7953)
);

INVx3_ASAP7_75t_L g7954 ( 
.A(n_7742),
.Y(n_7954)
);

AND2x2_ASAP7_75t_L g7955 ( 
.A(n_7695),
.B(n_5673),
.Y(n_7955)
);

AOI21xp5_ASAP7_75t_L g7956 ( 
.A1(n_7702),
.A2(n_5891),
.B(n_5888),
.Y(n_7956)
);

AND2x2_ASAP7_75t_L g7957 ( 
.A(n_7548),
.B(n_5673),
.Y(n_7957)
);

BUFx2_ASAP7_75t_SL g7958 ( 
.A(n_7511),
.Y(n_7958)
);

INVxp67_ASAP7_75t_L g7959 ( 
.A(n_7572),
.Y(n_7959)
);

INVx3_ASAP7_75t_L g7960 ( 
.A(n_7522),
.Y(n_7960)
);

INVx2_ASAP7_75t_L g7961 ( 
.A(n_7760),
.Y(n_7961)
);

INVx2_ASAP7_75t_L g7962 ( 
.A(n_7752),
.Y(n_7962)
);

AO21x2_ASAP7_75t_L g7963 ( 
.A1(n_7683),
.A2(n_5891),
.B(n_5888),
.Y(n_7963)
);

OR2x2_ASAP7_75t_L g7964 ( 
.A(n_7598),
.B(n_6029),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7507),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_7726),
.Y(n_7966)
);

INVx2_ASAP7_75t_L g7967 ( 
.A(n_7759),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_7729),
.Y(n_7968)
);

OAI33xp33_ASAP7_75t_L g7969 ( 
.A1(n_7655),
.A2(n_5907),
.A3(n_5895),
.B1(n_6044),
.B2(n_6047),
.B3(n_6029),
.Y(n_7969)
);

AND2x2_ASAP7_75t_L g7970 ( 
.A(n_7757),
.B(n_7736),
.Y(n_7970)
);

OAI21xp5_ASAP7_75t_SL g7971 ( 
.A1(n_7624),
.A2(n_4511),
.B(n_4494),
.Y(n_7971)
);

AOI22xp33_ASAP7_75t_L g7972 ( 
.A1(n_7692),
.A2(n_5895),
.B1(n_5907),
.B2(n_5702),
.Y(n_7972)
);

OAI211xp5_ASAP7_75t_SL g7973 ( 
.A1(n_7650),
.A2(n_5530),
.B(n_5573),
.C(n_5162),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_7741),
.Y(n_7974)
);

AOI221xp5_ASAP7_75t_L g7975 ( 
.A1(n_7514),
.A2(n_5573),
.B1(n_5914),
.B2(n_5911),
.C(n_5910),
.Y(n_7975)
);

HB1xp67_ASAP7_75t_L g7976 ( 
.A(n_7633),
.Y(n_7976)
);

INVx1_ASAP7_75t_L g7977 ( 
.A(n_7749),
.Y(n_7977)
);

INVx3_ASAP7_75t_L g7978 ( 
.A(n_7785),
.Y(n_7978)
);

OAI22xp5_ASAP7_75t_L g7979 ( 
.A1(n_7748),
.A2(n_5633),
.B1(n_5730),
.B2(n_5594),
.Y(n_7979)
);

OA211x2_ASAP7_75t_L g7980 ( 
.A1(n_7712),
.A2(n_4347),
.B(n_4275),
.C(n_3604),
.Y(n_7980)
);

AOI33xp33_ASAP7_75t_L g7981 ( 
.A1(n_7776),
.A2(n_6049),
.A3(n_6047),
.B1(n_6050),
.B2(n_6048),
.B3(n_6044),
.Y(n_7981)
);

AND2x2_ASAP7_75t_L g7982 ( 
.A(n_7754),
.B(n_5600),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_L g7983 ( 
.A(n_7654),
.B(n_6048),
.Y(n_7983)
);

OAI221xp5_ASAP7_75t_L g7984 ( 
.A1(n_7771),
.A2(n_6049),
.B1(n_6081),
.B2(n_6058),
.C(n_6050),
.Y(n_7984)
);

INVx1_ASAP7_75t_SL g7985 ( 
.A(n_7625),
.Y(n_7985)
);

INVx1_ASAP7_75t_L g7986 ( 
.A(n_7667),
.Y(n_7986)
);

AND2x2_ASAP7_75t_L g7987 ( 
.A(n_7672),
.B(n_7687),
.Y(n_7987)
);

INVx1_ASAP7_75t_SL g7988 ( 
.A(n_7784),
.Y(n_7988)
);

INVx1_ASAP7_75t_SL g7989 ( 
.A(n_7613),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7720),
.Y(n_7990)
);

BUFx2_ASAP7_75t_L g7991 ( 
.A(n_7668),
.Y(n_7991)
);

BUFx2_ASAP7_75t_L g7992 ( 
.A(n_7554),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_7559),
.Y(n_7993)
);

OAI21xp33_ASAP7_75t_L g7994 ( 
.A1(n_7535),
.A2(n_6084),
.B(n_6081),
.Y(n_7994)
);

INVx1_ASAP7_75t_SL g7995 ( 
.A(n_7718),
.Y(n_7995)
);

AND2x2_ASAP7_75t_L g7996 ( 
.A(n_7688),
.B(n_5600),
.Y(n_7996)
);

NAND2xp5_ASAP7_75t_L g7997 ( 
.A(n_7557),
.B(n_6084),
.Y(n_7997)
);

INVx1_ASAP7_75t_L g7998 ( 
.A(n_7560),
.Y(n_7998)
);

AND2x2_ASAP7_75t_L g7999 ( 
.A(n_7513),
.B(n_5559),
.Y(n_7999)
);

INVx2_ASAP7_75t_L g8000 ( 
.A(n_7758),
.Y(n_8000)
);

INVx1_ASAP7_75t_L g8001 ( 
.A(n_7564),
.Y(n_8001)
);

OR2x2_ASAP7_75t_L g8002 ( 
.A(n_7697),
.B(n_6105),
.Y(n_8002)
);

AOI22xp33_ASAP7_75t_L g8003 ( 
.A1(n_7788),
.A2(n_5702),
.B1(n_5911),
.B2(n_5910),
.Y(n_8003)
);

AND2x2_ASAP7_75t_L g8004 ( 
.A(n_7533),
.B(n_5559),
.Y(n_8004)
);

OAI22xp5_ASAP7_75t_SL g8005 ( 
.A1(n_7585),
.A2(n_4511),
.B1(n_4644),
.B2(n_4494),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7648),
.Y(n_8006)
);

NAND3xp33_ASAP7_75t_L g8007 ( 
.A(n_7615),
.B(n_7521),
.C(n_7621),
.Y(n_8007)
);

AND2x2_ASAP7_75t_L g8008 ( 
.A(n_7614),
.B(n_5576),
.Y(n_8008)
);

NAND2xp5_ASAP7_75t_L g8009 ( 
.A(n_7568),
.B(n_6099),
.Y(n_8009)
);

NAND2xp5_ASAP7_75t_SL g8010 ( 
.A(n_7551),
.B(n_4494),
.Y(n_8010)
);

AND2x2_ASAP7_75t_L g8011 ( 
.A(n_7707),
.B(n_5576),
.Y(n_8011)
);

NAND4xp25_ASAP7_75t_L g8012 ( 
.A(n_7619),
.B(n_5047),
.C(n_4387),
.D(n_4391),
.Y(n_8012)
);

NOR2x1_ASAP7_75t_L g8013 ( 
.A(n_7524),
.B(n_5047),
.Y(n_8013)
);

OAI22xp5_ASAP7_75t_L g8014 ( 
.A1(n_7586),
.A2(n_5633),
.B1(n_5730),
.B2(n_5464),
.Y(n_8014)
);

OAI21x1_ASAP7_75t_SL g8015 ( 
.A1(n_7716),
.A2(n_6105),
.B(n_6099),
.Y(n_8015)
);

OAI221xp5_ASAP7_75t_L g8016 ( 
.A1(n_7601),
.A2(n_6109),
.B1(n_6120),
.B2(n_6117),
.C(n_6114),
.Y(n_8016)
);

INVx2_ASAP7_75t_L g8017 ( 
.A(n_7764),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7586),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7704),
.Y(n_8019)
);

OR2x2_ASAP7_75t_L g8020 ( 
.A(n_7663),
.B(n_6187),
.Y(n_8020)
);

INVx1_ASAP7_75t_L g8021 ( 
.A(n_7783),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7691),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7581),
.B(n_6109),
.Y(n_8023)
);

AOI22xp33_ASAP7_75t_L g8024 ( 
.A1(n_7791),
.A2(n_5702),
.B1(n_5923),
.B2(n_5914),
.Y(n_8024)
);

OR2x6_ASAP7_75t_L g8025 ( 
.A(n_7597),
.B(n_5725),
.Y(n_8025)
);

INVx1_ASAP7_75t_L g8026 ( 
.A(n_7797),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7491),
.B(n_5589),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7725),
.B(n_5589),
.Y(n_8028)
);

AOI22xp5_ASAP7_75t_L g8029 ( 
.A1(n_7656),
.A2(n_5470),
.B1(n_5469),
.B2(n_5499),
.Y(n_8029)
);

AND2x2_ASAP7_75t_L g8030 ( 
.A(n_7665),
.B(n_5656),
.Y(n_8030)
);

NOR2x1_ASAP7_75t_L g8031 ( 
.A(n_7644),
.B(n_6114),
.Y(n_8031)
);

INVx1_ASAP7_75t_L g8032 ( 
.A(n_7616),
.Y(n_8032)
);

INVx2_ASAP7_75t_SL g8033 ( 
.A(n_7795),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7645),
.Y(n_8034)
);

INVx3_ASAP7_75t_L g8035 ( 
.A(n_7772),
.Y(n_8035)
);

OAI21xp5_ASAP7_75t_SL g8036 ( 
.A1(n_7594),
.A2(n_4511),
.B(n_4494),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_7679),
.Y(n_8037)
);

AND2x2_ASAP7_75t_L g8038 ( 
.A(n_7787),
.B(n_7790),
.Y(n_8038)
);

INVx1_ASAP7_75t_L g8039 ( 
.A(n_7719),
.Y(n_8039)
);

AND2x2_ASAP7_75t_L g8040 ( 
.A(n_7781),
.B(n_5656),
.Y(n_8040)
);

AOI221x1_ASAP7_75t_L g8041 ( 
.A1(n_7563),
.A2(n_7573),
.B1(n_7591),
.B2(n_7576),
.C(n_7575),
.Y(n_8041)
);

AND2x2_ASAP7_75t_L g8042 ( 
.A(n_7768),
.B(n_5667),
.Y(n_8042)
);

INVx1_ASAP7_75t_L g8043 ( 
.A(n_7762),
.Y(n_8043)
);

NAND2xp5_ASAP7_75t_L g8044 ( 
.A(n_7599),
.B(n_6117),
.Y(n_8044)
);

AND2x2_ASAP7_75t_L g8045 ( 
.A(n_7550),
.B(n_7678),
.Y(n_8045)
);

AND2x4_ASAP7_75t_L g8046 ( 
.A(n_7609),
.B(n_5730),
.Y(n_8046)
);

INVx1_ASAP7_75t_L g8047 ( 
.A(n_7684),
.Y(n_8047)
);

AND2x2_ASAP7_75t_L g8048 ( 
.A(n_7570),
.B(n_5667),
.Y(n_8048)
);

NAND3xp33_ASAP7_75t_L g8049 ( 
.A(n_7653),
.B(n_7661),
.C(n_7657),
.Y(n_8049)
);

AND2x2_ASAP7_75t_L g8050 ( 
.A(n_7583),
.B(n_5730),
.Y(n_8050)
);

INVx1_ASAP7_75t_L g8051 ( 
.A(n_7732),
.Y(n_8051)
);

OAI33xp33_ASAP7_75t_L g8052 ( 
.A1(n_7738),
.A2(n_6120),
.A3(n_6137),
.B1(n_6147),
.B2(n_6142),
.B3(n_6129),
.Y(n_8052)
);

BUFx2_ASAP7_75t_L g8053 ( 
.A(n_7703),
.Y(n_8053)
);

AND2x2_ASAP7_75t_L g8054 ( 
.A(n_7792),
.B(n_4494),
.Y(n_8054)
);

INVx2_ASAP7_75t_L g8055 ( 
.A(n_7779),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_7786),
.Y(n_8056)
);

AND2x4_ASAP7_75t_L g8057 ( 
.A(n_7643),
.B(n_6142),
.Y(n_8057)
);

NOR2xp33_ASAP7_75t_R g8058 ( 
.A(n_7635),
.B(n_4494),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_7676),
.Y(n_8059)
);

OR2x2_ASAP7_75t_L g8060 ( 
.A(n_7494),
.B(n_6221),
.Y(n_8060)
);

HB1xp67_ASAP7_75t_L g8061 ( 
.A(n_7629),
.Y(n_8061)
);

INVx2_ASAP7_75t_L g8062 ( 
.A(n_7731),
.Y(n_8062)
);

OR2x2_ASAP7_75t_L g8063 ( 
.A(n_7763),
.B(n_6221),
.Y(n_8063)
);

INVx1_ASAP7_75t_L g8064 ( 
.A(n_7735),
.Y(n_8064)
);

INVx2_ASAP7_75t_L g8065 ( 
.A(n_7682),
.Y(n_8065)
);

NAND2xp5_ASAP7_75t_L g8066 ( 
.A(n_7561),
.B(n_6129),
.Y(n_8066)
);

NAND2xp5_ASAP7_75t_L g8067 ( 
.A(n_7775),
.B(n_6137),
.Y(n_8067)
);

BUFx2_ASAP7_75t_L g8068 ( 
.A(n_7703),
.Y(n_8068)
);

NOR3xp33_ASAP7_75t_SL g8069 ( 
.A(n_7536),
.B(n_4681),
.C(n_4859),
.Y(n_8069)
);

INVx2_ASAP7_75t_L g8070 ( 
.A(n_7545),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7746),
.Y(n_8071)
);

INVx3_ASAP7_75t_L g8072 ( 
.A(n_7595),
.Y(n_8072)
);

AND2x2_ASAP7_75t_L g8073 ( 
.A(n_7722),
.B(n_4511),
.Y(n_8073)
);

OAI221xp5_ASAP7_75t_L g8074 ( 
.A1(n_7623),
.A2(n_6152),
.B1(n_6177),
.B2(n_6161),
.C(n_6147),
.Y(n_8074)
);

OR2x2_ASAP7_75t_L g8075 ( 
.A(n_7584),
.B(n_6212),
.Y(n_8075)
);

INVx1_ASAP7_75t_L g8076 ( 
.A(n_7602),
.Y(n_8076)
);

AOI221xp5_ASAP7_75t_L g8077 ( 
.A1(n_7693),
.A2(n_5930),
.B1(n_5932),
.B2(n_5923),
.C(n_5501),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7602),
.Y(n_8078)
);

INVx2_ASAP7_75t_L g8079 ( 
.A(n_7629),
.Y(n_8079)
);

NAND2xp5_ASAP7_75t_SL g8080 ( 
.A(n_7546),
.B(n_4511),
.Y(n_8080)
);

AND2x2_ASAP7_75t_L g8081 ( 
.A(n_7603),
.B(n_4511),
.Y(n_8081)
);

INVx1_ASAP7_75t_L g8082 ( 
.A(n_7700),
.Y(n_8082)
);

INVx1_ASAP7_75t_L g8083 ( 
.A(n_7603),
.Y(n_8083)
);

NOR2xp33_ASAP7_75t_L g8084 ( 
.A(n_7562),
.B(n_5093),
.Y(n_8084)
);

AND2x2_ASAP7_75t_L g8085 ( 
.A(n_7753),
.B(n_4644),
.Y(n_8085)
);

INVx4_ASAP7_75t_L g8086 ( 
.A(n_7639),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7639),
.Y(n_8087)
);

INVx5_ASAP7_75t_SL g8088 ( 
.A(n_7789),
.Y(n_8088)
);

OAI211xp5_ASAP7_75t_SL g8089 ( 
.A1(n_7675),
.A2(n_5162),
.B(n_5280),
.C(n_5253),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_7922),
.Y(n_8090)
);

NAND2x1_ASAP7_75t_L g8091 ( 
.A(n_7825),
.B(n_7773),
.Y(n_8091)
);

NAND2xp5_ASAP7_75t_L g8092 ( 
.A(n_7848),
.B(n_7767),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_7922),
.Y(n_8093)
);

INVx2_ASAP7_75t_L g8094 ( 
.A(n_7877),
.Y(n_8094)
);

INVx2_ASAP7_75t_L g8095 ( 
.A(n_7896),
.Y(n_8095)
);

INVx1_ASAP7_75t_L g8096 ( 
.A(n_7917),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_7849),
.Y(n_8097)
);

OR2x2_ASAP7_75t_L g8098 ( 
.A(n_7947),
.B(n_7677),
.Y(n_8098)
);

AND2x2_ASAP7_75t_L g8099 ( 
.A(n_7802),
.B(n_7734),
.Y(n_8099)
);

OR2x2_ASAP7_75t_L g8100 ( 
.A(n_7947),
.B(n_7755),
.Y(n_8100)
);

AOI22xp5_ASAP7_75t_L g8101 ( 
.A1(n_7934),
.A2(n_7761),
.B1(n_7705),
.B2(n_7744),
.Y(n_8101)
);

OR2x2_ASAP7_75t_L g8102 ( 
.A(n_7985),
.B(n_7743),
.Y(n_8102)
);

NAND2xp5_ASAP7_75t_L g8103 ( 
.A(n_7836),
.B(n_7798),
.Y(n_8103)
);

AND2x2_ASAP7_75t_L g8104 ( 
.A(n_7896),
.B(n_7756),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_L g8105 ( 
.A(n_7871),
.B(n_7579),
.Y(n_8105)
);

INVxp67_ASAP7_75t_L g8106 ( 
.A(n_7830),
.Y(n_8106)
);

INVx1_ASAP7_75t_L g8107 ( 
.A(n_7893),
.Y(n_8107)
);

BUFx2_ASAP7_75t_L g8108 ( 
.A(n_7804),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7815),
.Y(n_8109)
);

NAND2x1_ASAP7_75t_L g8110 ( 
.A(n_7838),
.B(n_7773),
.Y(n_8110)
);

AND2x2_ASAP7_75t_L g8111 ( 
.A(n_7804),
.B(n_7706),
.Y(n_8111)
);

AND2x2_ASAP7_75t_L g8112 ( 
.A(n_7801),
.B(n_7714),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7858),
.Y(n_8113)
);

NOR2xp33_ASAP7_75t_L g8114 ( 
.A(n_7838),
.B(n_7618),
.Y(n_8114)
);

INVx1_ASAP7_75t_L g8115 ( 
.A(n_7835),
.Y(n_8115)
);

HB1xp67_ASAP7_75t_L g8116 ( 
.A(n_8076),
.Y(n_8116)
);

AND2x2_ASAP7_75t_L g8117 ( 
.A(n_7809),
.B(n_7793),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7846),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_7799),
.Y(n_8119)
);

HB1xp67_ASAP7_75t_L g8120 ( 
.A(n_8076),
.Y(n_8120)
);

NAND2xp5_ASAP7_75t_L g8121 ( 
.A(n_7834),
.B(n_7549),
.Y(n_8121)
);

INVx2_ASAP7_75t_L g8122 ( 
.A(n_7860),
.Y(n_8122)
);

AND2x2_ASAP7_75t_L g8123 ( 
.A(n_7851),
.B(n_7793),
.Y(n_8123)
);

INVx2_ASAP7_75t_L g8124 ( 
.A(n_7856),
.Y(n_8124)
);

OR2x2_ASAP7_75t_L g8125 ( 
.A(n_7806),
.B(n_7739),
.Y(n_8125)
);

NAND2xp5_ASAP7_75t_L g8126 ( 
.A(n_7861),
.B(n_7567),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_7854),
.B(n_7701),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_7907),
.Y(n_8128)
);

AND2x4_ASAP7_75t_L g8129 ( 
.A(n_7805),
.B(n_6259),
.Y(n_8129)
);

NAND2xp5_ASAP7_75t_L g8130 ( 
.A(n_7939),
.B(n_7737),
.Y(n_8130)
);

AND2x2_ASAP7_75t_L g8131 ( 
.A(n_7843),
.B(n_4644),
.Y(n_8131)
);

AND2x2_ASAP7_75t_L g8132 ( 
.A(n_7813),
.B(n_4644),
.Y(n_8132)
);

INVx2_ASAP7_75t_SL g8133 ( 
.A(n_7824),
.Y(n_8133)
);

NAND2xp5_ASAP7_75t_L g8134 ( 
.A(n_7939),
.B(n_6152),
.Y(n_8134)
);

O2A1O1Ixp5_ASAP7_75t_R g8135 ( 
.A1(n_7857),
.A2(n_7789),
.B(n_5253),
.C(n_5280),
.Y(n_8135)
);

INVxp67_ASAP7_75t_L g8136 ( 
.A(n_7938),
.Y(n_8136)
);

AND2x2_ASAP7_75t_L g8137 ( 
.A(n_7839),
.B(n_4644),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7856),
.Y(n_8138)
);

AND2x2_ASAP7_75t_L g8139 ( 
.A(n_7897),
.B(n_4644),
.Y(n_8139)
);

OR2x2_ASAP7_75t_L g8140 ( 
.A(n_7811),
.B(n_6161),
.Y(n_8140)
);

OR2x2_ASAP7_75t_L g8141 ( 
.A(n_7803),
.B(n_6177),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7951),
.Y(n_8142)
);

INVx2_ASAP7_75t_L g8143 ( 
.A(n_7812),
.Y(n_8143)
);

INVx2_ASAP7_75t_L g8144 ( 
.A(n_7812),
.Y(n_8144)
);

AND2x2_ASAP7_75t_L g8145 ( 
.A(n_7914),
.B(n_4658),
.Y(n_8145)
);

NOR2xp33_ASAP7_75t_L g8146 ( 
.A(n_7933),
.B(n_4683),
.Y(n_8146)
);

NOR2xp67_ASAP7_75t_SL g8147 ( 
.A(n_7958),
.B(n_4658),
.Y(n_8147)
);

INVx1_ASAP7_75t_L g8148 ( 
.A(n_7952),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7894),
.Y(n_8149)
);

INVx2_ASAP7_75t_L g8150 ( 
.A(n_7924),
.Y(n_8150)
);

INVx1_ASAP7_75t_SL g8151 ( 
.A(n_7992),
.Y(n_8151)
);

INVx2_ASAP7_75t_L g8152 ( 
.A(n_7924),
.Y(n_8152)
);

INVxp67_ASAP7_75t_L g8153 ( 
.A(n_7928),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_SL g8154 ( 
.A(n_7933),
.B(n_4658),
.Y(n_8154)
);

INVx2_ASAP7_75t_L g8155 ( 
.A(n_7865),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7913),
.Y(n_8156)
);

NAND2xp5_ASAP7_75t_L g8157 ( 
.A(n_7865),
.B(n_6180),
.Y(n_8157)
);

OR2x2_ASAP7_75t_L g8158 ( 
.A(n_8086),
.B(n_6180),
.Y(n_8158)
);

OAI21xp5_ASAP7_75t_SL g8159 ( 
.A1(n_7971),
.A2(n_8087),
.B(n_8078),
.Y(n_8159)
);

INVx2_ASAP7_75t_SL g8160 ( 
.A(n_7941),
.Y(n_8160)
);

INVx2_ASAP7_75t_SL g8161 ( 
.A(n_7941),
.Y(n_8161)
);

INVx1_ASAP7_75t_L g8162 ( 
.A(n_7915),
.Y(n_8162)
);

NAND2x1p5_ASAP7_75t_L g8163 ( 
.A(n_7923),
.B(n_4658),
.Y(n_8163)
);

AND2x2_ASAP7_75t_L g8164 ( 
.A(n_7955),
.B(n_4658),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_7870),
.Y(n_8165)
);

INVx1_ASAP7_75t_L g8166 ( 
.A(n_7800),
.Y(n_8166)
);

NAND2xp5_ASAP7_75t_SL g8167 ( 
.A(n_8086),
.B(n_4658),
.Y(n_8167)
);

AND2x2_ASAP7_75t_L g8168 ( 
.A(n_7937),
.B(n_4683),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7800),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_7800),
.Y(n_8170)
);

INVx1_ASAP7_75t_L g8171 ( 
.A(n_7816),
.Y(n_8171)
);

INVx1_ASAP7_75t_L g8172 ( 
.A(n_7818),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7822),
.Y(n_8173)
);

INVx1_ASAP7_75t_SL g8174 ( 
.A(n_7869),
.Y(n_8174)
);

OR2x2_ASAP7_75t_L g8175 ( 
.A(n_7995),
.B(n_6187),
.Y(n_8175)
);

AND2x2_ASAP7_75t_L g8176 ( 
.A(n_7807),
.B(n_4683),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_7827),
.Y(n_8177)
);

NAND2xp5_ASAP7_75t_SL g8178 ( 
.A(n_7960),
.B(n_4683),
.Y(n_8178)
);

BUFx2_ASAP7_75t_L g8179 ( 
.A(n_8058),
.Y(n_8179)
);

NAND2xp5_ASAP7_75t_L g8180 ( 
.A(n_7988),
.B(n_6205),
.Y(n_8180)
);

NOR2x1_ASAP7_75t_L g8181 ( 
.A(n_8078),
.B(n_6205),
.Y(n_8181)
);

AND2x2_ASAP7_75t_L g8182 ( 
.A(n_7826),
.B(n_4683),
.Y(n_8182)
);

HB1xp67_ASAP7_75t_L g8183 ( 
.A(n_8087),
.Y(n_8183)
);

NOR2x1p5_ASAP7_75t_L g8184 ( 
.A(n_7837),
.B(n_4683),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7840),
.Y(n_8185)
);

NAND2x1p5_ASAP7_75t_L g8186 ( 
.A(n_7954),
.B(n_4739),
.Y(n_8186)
);

NAND2xp5_ASAP7_75t_L g8187 ( 
.A(n_7887),
.B(n_6206),
.Y(n_8187)
);

OR2x2_ASAP7_75t_L g8188 ( 
.A(n_7845),
.B(n_6206),
.Y(n_8188)
);

NAND2xp5_ASAP7_75t_L g8189 ( 
.A(n_7831),
.B(n_6210),
.Y(n_8189)
);

INVx2_ASAP7_75t_SL g8190 ( 
.A(n_7942),
.Y(n_8190)
);

NOR2xp67_ASAP7_75t_L g8191 ( 
.A(n_7927),
.B(n_6229),
.Y(n_8191)
);

INVx1_ASAP7_75t_L g8192 ( 
.A(n_7878),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7863),
.Y(n_8193)
);

AND2x2_ASAP7_75t_L g8194 ( 
.A(n_7821),
.B(n_4739),
.Y(n_8194)
);

HB1xp67_ASAP7_75t_L g8195 ( 
.A(n_7963),
.Y(n_8195)
);

AND2x2_ASAP7_75t_L g8196 ( 
.A(n_7999),
.B(n_4739),
.Y(n_8196)
);

OR2x2_ASAP7_75t_L g8197 ( 
.A(n_7990),
.B(n_6210),
.Y(n_8197)
);

NAND2xp5_ASAP7_75t_SL g8198 ( 
.A(n_7960),
.B(n_7852),
.Y(n_8198)
);

NAND2xp5_ASAP7_75t_L g8199 ( 
.A(n_8048),
.B(n_6212),
.Y(n_8199)
);

AND2x4_ASAP7_75t_L g8200 ( 
.A(n_7967),
.B(n_6248),
.Y(n_8200)
);

INVx2_ASAP7_75t_L g8201 ( 
.A(n_7942),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7948),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_7964),
.Y(n_8203)
);

AND2x4_ASAP7_75t_L g8204 ( 
.A(n_8000),
.B(n_6248),
.Y(n_8204)
);

NAND2xp5_ASAP7_75t_L g8205 ( 
.A(n_7864),
.B(n_6215),
.Y(n_8205)
);

NAND2xp5_ASAP7_75t_L g8206 ( 
.A(n_8030),
.B(n_6215),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_7829),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_7892),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_7908),
.Y(n_8209)
);

BUFx2_ASAP7_75t_L g8210 ( 
.A(n_8025),
.Y(n_8210)
);

OAI33xp33_ASAP7_75t_L g8211 ( 
.A1(n_8082),
.A2(n_5932),
.A3(n_5930),
.B1(n_6224),
.B2(n_6229),
.B3(n_6223),
.Y(n_8211)
);

INVx1_ASAP7_75t_SL g8212 ( 
.A(n_7989),
.Y(n_8212)
);

AOI21x1_ASAP7_75t_L g8213 ( 
.A1(n_7853),
.A2(n_6224),
.B(n_6223),
.Y(n_8213)
);

INVx1_ASAP7_75t_L g8214 ( 
.A(n_7950),
.Y(n_8214)
);

NAND2xp5_ASAP7_75t_L g8215 ( 
.A(n_7961),
.B(n_6232),
.Y(n_8215)
);

AND2x2_ASAP7_75t_L g8216 ( 
.A(n_8004),
.B(n_7957),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_L g8217 ( 
.A(n_8043),
.B(n_6232),
.Y(n_8217)
);

AND2x2_ASAP7_75t_L g8218 ( 
.A(n_8027),
.B(n_4739),
.Y(n_8218)
);

BUFx2_ASAP7_75t_L g8219 ( 
.A(n_8025),
.Y(n_8219)
);

INVx2_ASAP7_75t_L g8220 ( 
.A(n_7954),
.Y(n_8220)
);

INVx1_ASAP7_75t_L g8221 ( 
.A(n_8002),
.Y(n_8221)
);

INVx1_ASAP7_75t_SL g8222 ( 
.A(n_7987),
.Y(n_8222)
);

OAI22xp5_ASAP7_75t_L g8223 ( 
.A1(n_8083),
.A2(n_7976),
.B1(n_7986),
.B2(n_8007),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_7890),
.Y(n_8224)
);

AND2x4_ASAP7_75t_SL g8225 ( 
.A(n_7970),
.B(n_4739),
.Y(n_8225)
);

INVxp67_ASAP7_75t_SL g8226 ( 
.A(n_8083),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7859),
.Y(n_8227)
);

INVx3_ASAP7_75t_SL g8228 ( 
.A(n_7944),
.Y(n_8228)
);

AND2x2_ASAP7_75t_L g8229 ( 
.A(n_8040),
.B(n_4739),
.Y(n_8229)
);

AND2x2_ASAP7_75t_L g8230 ( 
.A(n_8008),
.B(n_4770),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_8026),
.B(n_6249),
.Y(n_8231)
);

AND2x2_ASAP7_75t_L g8232 ( 
.A(n_8045),
.B(n_4770),
.Y(n_8232)
);

INVx1_ASAP7_75t_L g8233 ( 
.A(n_7900),
.Y(n_8233)
);

AND2x4_ASAP7_75t_SL g8234 ( 
.A(n_7832),
.B(n_4775),
.Y(n_8234)
);

AND2x2_ASAP7_75t_L g8235 ( 
.A(n_8046),
.B(n_4770),
.Y(n_8235)
);

INVx2_ASAP7_75t_L g8236 ( 
.A(n_7996),
.Y(n_8236)
);

INVxp33_ASAP7_75t_L g8237 ( 
.A(n_8084),
.Y(n_8237)
);

OAI22xp33_ASAP7_75t_L g8238 ( 
.A1(n_8082),
.A2(n_5335),
.B1(n_5329),
.B2(n_6249),
.Y(n_8238)
);

INVx1_ASAP7_75t_L g8239 ( 
.A(n_7901),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_8035),
.Y(n_8240)
);

AND2x2_ASAP7_75t_L g8241 ( 
.A(n_8046),
.B(n_8050),
.Y(n_8241)
);

INVx2_ASAP7_75t_L g8242 ( 
.A(n_7889),
.Y(n_8242)
);

AND2x2_ASAP7_75t_L g8243 ( 
.A(n_7982),
.B(n_4770),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_8035),
.Y(n_8244)
);

OAI22xp5_ASAP7_75t_L g8245 ( 
.A1(n_7986),
.A2(n_6259),
.B1(n_6256),
.B2(n_5253),
.Y(n_8245)
);

OAI21xp5_ASAP7_75t_L g8246 ( 
.A1(n_7808),
.A2(n_6235),
.B(n_5856),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_7959),
.B(n_4770),
.Y(n_8247)
);

OR2x2_ASAP7_75t_L g8248 ( 
.A(n_7819),
.B(n_6256),
.Y(n_8248)
);

INVxp67_ASAP7_75t_L g8249 ( 
.A(n_8061),
.Y(n_8249)
);

NAND2xp5_ASAP7_75t_L g8250 ( 
.A(n_8021),
.B(n_5360),
.Y(n_8250)
);

NAND3xp33_ASAP7_75t_L g8251 ( 
.A(n_7879),
.B(n_5501),
.C(n_5446),
.Y(n_8251)
);

INVx2_ASAP7_75t_L g8252 ( 
.A(n_8015),
.Y(n_8252)
);

AND2x2_ASAP7_75t_L g8253 ( 
.A(n_7910),
.B(n_4770),
.Y(n_8253)
);

NOR2xp33_ASAP7_75t_L g8254 ( 
.A(n_8012),
.B(n_4775),
.Y(n_8254)
);

INVx1_ASAP7_75t_L g8255 ( 
.A(n_7867),
.Y(n_8255)
);

INVx1_ASAP7_75t_L g8256 ( 
.A(n_7872),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7874),
.Y(n_8257)
);

HB1xp67_ASAP7_75t_L g8258 ( 
.A(n_7868),
.Y(n_8258)
);

NAND2xp5_ASAP7_75t_L g8259 ( 
.A(n_7968),
.B(n_5360),
.Y(n_8259)
);

NOR2xp33_ASAP7_75t_L g8260 ( 
.A(n_7969),
.B(n_8036),
.Y(n_8260)
);

INVx1_ASAP7_75t_L g8261 ( 
.A(n_7902),
.Y(n_8261)
);

OR2x2_ASAP7_75t_L g8262 ( 
.A(n_7814),
.B(n_5361),
.Y(n_8262)
);

INVx2_ASAP7_75t_SL g8263 ( 
.A(n_8081),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_7881),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_7881),
.Y(n_8265)
);

NAND2xp5_ASAP7_75t_SL g8266 ( 
.A(n_7844),
.B(n_4775),
.Y(n_8266)
);

AND2x2_ASAP7_75t_L g8267 ( 
.A(n_8011),
.B(n_4775),
.Y(n_8267)
);

INVx1_ASAP7_75t_L g8268 ( 
.A(n_7875),
.Y(n_8268)
);

NAND2x1_ASAP7_75t_SL g8269 ( 
.A(n_8013),
.B(n_8072),
.Y(n_8269)
);

AND2x2_ASAP7_75t_L g8270 ( 
.A(n_7876),
.B(n_4775),
.Y(n_8270)
);

AND2x2_ASAP7_75t_L g8271 ( 
.A(n_8028),
.B(n_4775),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_7966),
.B(n_7974),
.Y(n_8272)
);

AND2x2_ASAP7_75t_L g8273 ( 
.A(n_8042),
.B(n_8073),
.Y(n_8273)
);

OAI21xp5_ASAP7_75t_L g8274 ( 
.A1(n_8049),
.A2(n_6235),
.B(n_5856),
.Y(n_8274)
);

HB1xp67_ASAP7_75t_L g8275 ( 
.A(n_7855),
.Y(n_8275)
);

NAND3xp33_ASAP7_75t_L g8276 ( 
.A(n_7898),
.B(n_5446),
.C(n_5442),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_7866),
.Y(n_8277)
);

INVxp67_ASAP7_75t_L g8278 ( 
.A(n_7991),
.Y(n_8278)
);

OR2x2_ASAP7_75t_L g8279 ( 
.A(n_7828),
.B(n_5361),
.Y(n_8279)
);

NOR2xp33_ASAP7_75t_L g8280 ( 
.A(n_7903),
.B(n_4862),
.Y(n_8280)
);

NOR2xp33_ASAP7_75t_L g8281 ( 
.A(n_7920),
.B(n_4862),
.Y(n_8281)
);

INVx1_ASAP7_75t_L g8282 ( 
.A(n_7810),
.Y(n_8282)
);

HB1xp67_ASAP7_75t_L g8283 ( 
.A(n_8072),
.Y(n_8283)
);

INVx1_ASAP7_75t_L g8284 ( 
.A(n_7810),
.Y(n_8284)
);

NAND2xp5_ASAP7_75t_L g8285 ( 
.A(n_7977),
.B(n_5363),
.Y(n_8285)
);

NAND2xp5_ASAP7_75t_L g8286 ( 
.A(n_8018),
.B(n_5363),
.Y(n_8286)
);

AOI21xp33_ASAP7_75t_L g8287 ( 
.A1(n_7873),
.A2(n_6158),
.B(n_6055),
.Y(n_8287)
);

AOI21xp5_ASAP7_75t_L g8288 ( 
.A1(n_7847),
.A2(n_5237),
.B(n_5236),
.Y(n_8288)
);

INVx2_ASAP7_75t_L g8289 ( 
.A(n_8063),
.Y(n_8289)
);

AND2x2_ASAP7_75t_L g8290 ( 
.A(n_8038),
.B(n_4778),
.Y(n_8290)
);

AND2x2_ASAP7_75t_L g8291 ( 
.A(n_8070),
.B(n_4778),
.Y(n_8291)
);

OR2x6_ASAP7_75t_L g8292 ( 
.A(n_7993),
.B(n_5329),
.Y(n_8292)
);

INVx1_ASAP7_75t_SL g8293 ( 
.A(n_7880),
.Y(n_8293)
);

OR3x2_ASAP7_75t_L g8294 ( 
.A(n_7850),
.B(n_3506),
.C(n_3882),
.Y(n_8294)
);

NAND2xp5_ASAP7_75t_L g8295 ( 
.A(n_8018),
.B(n_5364),
.Y(n_8295)
);

AND2x2_ASAP7_75t_L g8296 ( 
.A(n_7925),
.B(n_4778),
.Y(n_8296)
);

AND2x2_ASAP7_75t_L g8297 ( 
.A(n_8032),
.B(n_4778),
.Y(n_8297)
);

INVx3_ASAP7_75t_L g8298 ( 
.A(n_8088),
.Y(n_8298)
);

AND2x2_ASAP7_75t_L g8299 ( 
.A(n_8034),
.B(n_4778),
.Y(n_8299)
);

NAND2xp5_ASAP7_75t_L g8300 ( 
.A(n_8065),
.B(n_5364),
.Y(n_8300)
);

OR2x2_ASAP7_75t_L g8301 ( 
.A(n_7911),
.B(n_5366),
.Y(n_8301)
);

INVx1_ASAP7_75t_L g8302 ( 
.A(n_7906),
.Y(n_8302)
);

AND2x2_ASAP7_75t_L g8303 ( 
.A(n_8006),
.B(n_4778),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_L g8304 ( 
.A(n_8057),
.B(n_5366),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_7842),
.Y(n_8305)
);

NAND2xp5_ASAP7_75t_L g8306 ( 
.A(n_8057),
.B(n_5369),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_7899),
.Y(n_8307)
);

AND2x2_ASAP7_75t_L g8308 ( 
.A(n_7943),
.B(n_8088),
.Y(n_8308)
);

NAND2xp5_ASAP7_75t_L g8309 ( 
.A(n_7823),
.B(n_5369),
.Y(n_8309)
);

AOI22xp5_ASAP7_75t_L g8310 ( 
.A1(n_8019),
.A2(n_5469),
.B1(n_5470),
.B2(n_5451),
.Y(n_8310)
);

OR2x2_ASAP7_75t_L g8311 ( 
.A(n_7930),
.B(n_5380),
.Y(n_8311)
);

AND2x2_ASAP7_75t_L g8312 ( 
.A(n_7998),
.B(n_4783),
.Y(n_8312)
);

INVx3_ASAP7_75t_L g8313 ( 
.A(n_8056),
.Y(n_8313)
);

INVx1_ASAP7_75t_L g8314 ( 
.A(n_7899),
.Y(n_8314)
);

INVx2_ASAP7_75t_L g8315 ( 
.A(n_7891),
.Y(n_8315)
);

INVx2_ASAP7_75t_SL g8316 ( 
.A(n_8060),
.Y(n_8316)
);

AND2x4_ASAP7_75t_L g8317 ( 
.A(n_8041),
.B(n_5287),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_7916),
.Y(n_8318)
);

AND2x2_ASAP7_75t_L g8319 ( 
.A(n_8001),
.B(n_4783),
.Y(n_8319)
);

OAI21xp33_ASAP7_75t_L g8320 ( 
.A1(n_8069),
.A2(n_5242),
.B(n_5236),
.Y(n_8320)
);

OR2x2_ASAP7_75t_L g8321 ( 
.A(n_8075),
.B(n_5380),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7916),
.Y(n_8322)
);

AND2x2_ASAP7_75t_L g8323 ( 
.A(n_7817),
.B(n_4783),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_7931),
.Y(n_8324)
);

AND2x4_ASAP7_75t_L g8325 ( 
.A(n_8053),
.B(n_8068),
.Y(n_8325)
);

BUFx2_ASAP7_75t_L g8326 ( 
.A(n_8031),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_7931),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_L g8328 ( 
.A(n_8037),
.B(n_5381),
.Y(n_8328)
);

NAND2xp5_ASAP7_75t_L g8329 ( 
.A(n_8047),
.B(n_8051),
.Y(n_8329)
);

AND2x2_ASAP7_75t_L g8330 ( 
.A(n_8022),
.B(n_4783),
.Y(n_8330)
);

NOR2xp33_ASAP7_75t_L g8331 ( 
.A(n_8010),
.B(n_4783),
.Y(n_8331)
);

NAND2xp5_ASAP7_75t_SL g8332 ( 
.A(n_8017),
.B(n_4783),
.Y(n_8332)
);

INVx2_ASAP7_75t_SL g8333 ( 
.A(n_8054),
.Y(n_8333)
);

NAND2xp5_ASAP7_75t_L g8334 ( 
.A(n_8064),
.B(n_5381),
.Y(n_8334)
);

NAND2x1_ASAP7_75t_SL g8335 ( 
.A(n_8079),
.B(n_5162),
.Y(n_8335)
);

INVx1_ASAP7_75t_L g8336 ( 
.A(n_7885),
.Y(n_8336)
);

INVxp67_ASAP7_75t_L g8337 ( 
.A(n_8154),
.Y(n_8337)
);

AOI21xp33_ASAP7_75t_L g8338 ( 
.A1(n_8277),
.A2(n_8039),
.B(n_8019),
.Y(n_8338)
);

AND2x2_ASAP7_75t_L g8339 ( 
.A(n_8216),
.B(n_8071),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_8096),
.Y(n_8340)
);

AND2x2_ASAP7_75t_L g8341 ( 
.A(n_8095),
.B(n_8228),
.Y(n_8341)
);

INVx2_ASAP7_75t_L g8342 ( 
.A(n_8108),
.Y(n_8342)
);

AOI22xp33_ASAP7_75t_L g8343 ( 
.A1(n_8305),
.A2(n_8062),
.B1(n_8039),
.B2(n_8059),
.Y(n_8343)
);

INVx1_ASAP7_75t_L g8344 ( 
.A(n_8283),
.Y(n_8344)
);

INVx1_ASAP7_75t_L g8345 ( 
.A(n_8096),
.Y(n_8345)
);

OR2x2_ASAP7_75t_L g8346 ( 
.A(n_8293),
.B(n_8020),
.Y(n_8346)
);

INVx1_ASAP7_75t_L g8347 ( 
.A(n_8195),
.Y(n_8347)
);

NAND2xp5_ASAP7_75t_L g8348 ( 
.A(n_8133),
.B(n_8055),
.Y(n_8348)
);

OR2x2_ASAP7_75t_L g8349 ( 
.A(n_8151),
.B(n_7929),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_8275),
.Y(n_8350)
);

HB1xp67_ASAP7_75t_L g8351 ( 
.A(n_8183),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_8122),
.Y(n_8352)
);

NAND2xp5_ASAP7_75t_L g8353 ( 
.A(n_8222),
.B(n_8033),
.Y(n_8353)
);

NAND2xp5_ASAP7_75t_L g8354 ( 
.A(n_8106),
.B(n_7962),
.Y(n_8354)
);

INVx2_ASAP7_75t_L g8355 ( 
.A(n_8335),
.Y(n_8355)
);

NAND2xp5_ASAP7_75t_SL g8356 ( 
.A(n_8298),
.B(n_8005),
.Y(n_8356)
);

INVx2_ASAP7_75t_L g8357 ( 
.A(n_8163),
.Y(n_8357)
);

OAI322xp33_ASAP7_75t_L g8358 ( 
.A1(n_8277),
.A2(n_7884),
.A3(n_8066),
.B1(n_7945),
.B2(n_8023),
.C1(n_7997),
.C2(n_8044),
.Y(n_8358)
);

INVx3_ASAP7_75t_L g8359 ( 
.A(n_8298),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_8107),
.Y(n_8360)
);

AOI21xp5_ASAP7_75t_L g8361 ( 
.A1(n_8198),
.A2(n_7862),
.B(n_7883),
.Y(n_8361)
);

OAI22xp5_ASAP7_75t_L g8362 ( 
.A1(n_8302),
.A2(n_7820),
.B1(n_7882),
.B2(n_7926),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_8166),
.Y(n_8363)
);

NAND2xp5_ASAP7_75t_L g8364 ( 
.A(n_8155),
.B(n_7978),
.Y(n_8364)
);

OR2x2_ASAP7_75t_L g8365 ( 
.A(n_8113),
.B(n_7946),
.Y(n_8365)
);

O2A1O1Ixp33_ASAP7_75t_L g8366 ( 
.A1(n_8116),
.A2(n_7888),
.B(n_7895),
.C(n_7886),
.Y(n_8366)
);

NOR2xp33_ASAP7_75t_L g8367 ( 
.A(n_8153),
.B(n_8052),
.Y(n_8367)
);

INVx1_ASAP7_75t_L g8368 ( 
.A(n_8169),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_8170),
.Y(n_8369)
);

INVx2_ASAP7_75t_L g8370 ( 
.A(n_8186),
.Y(n_8370)
);

INVx1_ASAP7_75t_L g8371 ( 
.A(n_8226),
.Y(n_8371)
);

AOI21xp33_ASAP7_75t_SL g8372 ( 
.A1(n_8302),
.A2(n_7965),
.B(n_8080),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_8092),
.Y(n_8373)
);

INVx2_ASAP7_75t_L g8374 ( 
.A(n_8269),
.Y(n_8374)
);

NOR2x1_ASAP7_75t_L g8375 ( 
.A(n_8159),
.B(n_7909),
.Y(n_8375)
);

INVx1_ASAP7_75t_SL g8376 ( 
.A(n_8174),
.Y(n_8376)
);

NAND2xp5_ASAP7_75t_L g8377 ( 
.A(n_8129),
.B(n_8160),
.Y(n_8377)
);

AOI22xp33_ASAP7_75t_L g8378 ( 
.A1(n_8305),
.A2(n_8024),
.B1(n_8003),
.B2(n_7972),
.Y(n_8378)
);

OAI21xp5_ASAP7_75t_SL g8379 ( 
.A1(n_8136),
.A2(n_7973),
.B(n_7994),
.Y(n_8379)
);

AND2x2_ASAP7_75t_L g8380 ( 
.A(n_8109),
.B(n_7918),
.Y(n_8380)
);

INVx1_ASAP7_75t_L g8381 ( 
.A(n_8143),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_8144),
.Y(n_8382)
);

OAI22xp33_ASAP7_75t_SL g8383 ( 
.A1(n_8326),
.A2(n_7983),
.B1(n_7949),
.B2(n_8009),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_8184),
.Y(n_8384)
);

AOI211xp5_ASAP7_75t_SL g8385 ( 
.A1(n_8223),
.A2(n_7932),
.B(n_7912),
.C(n_7841),
.Y(n_8385)
);

OR2x2_ASAP7_75t_L g8386 ( 
.A(n_8094),
.B(n_8067),
.Y(n_8386)
);

INVx2_ASAP7_75t_L g8387 ( 
.A(n_8294),
.Y(n_8387)
);

OR2x2_ASAP7_75t_L g8388 ( 
.A(n_8119),
.B(n_7978),
.Y(n_8388)
);

AOI22xp5_ASAP7_75t_L g8389 ( 
.A1(n_8212),
.A2(n_8101),
.B1(n_8120),
.B2(n_8097),
.Y(n_8389)
);

INVx2_ASAP7_75t_L g8390 ( 
.A(n_8129),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_8097),
.Y(n_8391)
);

INVxp67_ASAP7_75t_L g8392 ( 
.A(n_8146),
.Y(n_8392)
);

OR2x2_ASAP7_75t_L g8393 ( 
.A(n_8236),
.B(n_7956),
.Y(n_8393)
);

AND2x2_ASAP7_75t_L g8394 ( 
.A(n_8232),
.B(n_7921),
.Y(n_8394)
);

INVx2_ASAP7_75t_L g8395 ( 
.A(n_8292),
.Y(n_8395)
);

AND2x2_ASAP7_75t_L g8396 ( 
.A(n_8112),
.B(n_7940),
.Y(n_8396)
);

OR2x2_ASAP7_75t_L g8397 ( 
.A(n_8316),
.B(n_8014),
.Y(n_8397)
);

INVx1_ASAP7_75t_L g8398 ( 
.A(n_8213),
.Y(n_8398)
);

INVx1_ASAP7_75t_L g8399 ( 
.A(n_8140),
.Y(n_8399)
);

INVx3_ASAP7_75t_L g8400 ( 
.A(n_8317),
.Y(n_8400)
);

INVxp67_ASAP7_75t_SL g8401 ( 
.A(n_8091),
.Y(n_8401)
);

OR2x2_ASAP7_75t_L g8402 ( 
.A(n_8165),
.B(n_7979),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_8141),
.Y(n_8403)
);

NOR4xp25_ASAP7_75t_L g8404 ( 
.A(n_8098),
.B(n_7833),
.C(n_7936),
.D(n_7953),
.Y(n_8404)
);

AOI21xp33_ASAP7_75t_SL g8405 ( 
.A1(n_8100),
.A2(n_8085),
.B(n_7984),
.Y(n_8405)
);

NOR3xp33_ASAP7_75t_L g8406 ( 
.A(n_8249),
.B(n_7981),
.C(n_8077),
.Y(n_8406)
);

INVx1_ASAP7_75t_SL g8407 ( 
.A(n_8123),
.Y(n_8407)
);

INVx1_ASAP7_75t_L g8408 ( 
.A(n_8181),
.Y(n_8408)
);

INVx1_ASAP7_75t_L g8409 ( 
.A(n_8130),
.Y(n_8409)
);

INVx1_ASAP7_75t_L g8410 ( 
.A(n_8188),
.Y(n_8410)
);

INVx2_ASAP7_75t_L g8411 ( 
.A(n_8292),
.Y(n_8411)
);

OR2x2_ASAP7_75t_L g8412 ( 
.A(n_8161),
.B(n_7904),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_8158),
.Y(n_8413)
);

AOI33xp33_ASAP7_75t_L g8414 ( 
.A1(n_8241),
.A2(n_7935),
.A3(n_7975),
.B1(n_8029),
.B2(n_7919),
.B3(n_8089),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_8128),
.Y(n_8415)
);

AND2x2_ASAP7_75t_L g8416 ( 
.A(n_8290),
.B(n_7905),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_8242),
.Y(n_8417)
);

OAI22xp5_ASAP7_75t_L g8418 ( 
.A1(n_8103),
.A2(n_7980),
.B1(n_8016),
.B2(n_8074),
.Y(n_8418)
);

AND2x2_ASAP7_75t_L g8419 ( 
.A(n_8182),
.B(n_4789),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_8175),
.Y(n_8420)
);

OAI221xp5_ASAP7_75t_L g8421 ( 
.A1(n_8287),
.A2(n_5451),
.B1(n_5455),
.B2(n_5450),
.C(n_5447),
.Y(n_8421)
);

OAI32xp33_ASAP7_75t_L g8422 ( 
.A1(n_8105),
.A2(n_5280),
.A3(n_5287),
.B1(n_5253),
.B2(n_5162),
.Y(n_8422)
);

OR2x2_ASAP7_75t_L g8423 ( 
.A(n_8190),
.B(n_5242),
.Y(n_8423)
);

OAI221xp5_ASAP7_75t_L g8424 ( 
.A1(n_8274),
.A2(n_5450),
.B1(n_5455),
.B2(n_5456),
.C(n_5447),
.Y(n_8424)
);

OR2x2_ASAP7_75t_L g8425 ( 
.A(n_8272),
.B(n_5245),
.Y(n_8425)
);

NOR2xp33_ASAP7_75t_L g8426 ( 
.A(n_8278),
.B(n_4789),
.Y(n_8426)
);

INVx2_ASAP7_75t_L g8427 ( 
.A(n_8137),
.Y(n_8427)
);

NAND2xp5_ASAP7_75t_L g8428 ( 
.A(n_8124),
.B(n_5385),
.Y(n_8428)
);

AND2x4_ASAP7_75t_L g8429 ( 
.A(n_8201),
.B(n_5280),
.Y(n_8429)
);

NAND2x1p5_ASAP7_75t_L g8430 ( 
.A(n_8220),
.B(n_4789),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_8307),
.Y(n_8431)
);

AOI21xp5_ASAP7_75t_L g8432 ( 
.A1(n_8266),
.A2(n_5252),
.B(n_5245),
.Y(n_8432)
);

OR2x2_ASAP7_75t_L g8433 ( 
.A(n_8214),
.B(n_5252),
.Y(n_8433)
);

INVx2_ASAP7_75t_L g8434 ( 
.A(n_8131),
.Y(n_8434)
);

INVx1_ASAP7_75t_L g8435 ( 
.A(n_8307),
.Y(n_8435)
);

AOI21xp5_ASAP7_75t_L g8436 ( 
.A1(n_8317),
.A2(n_5262),
.B(n_5258),
.Y(n_8436)
);

INVx2_ASAP7_75t_L g8437 ( 
.A(n_8132),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_8176),
.B(n_4789),
.Y(n_8438)
);

AO21x1_ASAP7_75t_L g8439 ( 
.A1(n_8110),
.A2(n_5262),
.B(n_5258),
.Y(n_8439)
);

OR2x2_ASAP7_75t_L g8440 ( 
.A(n_8126),
.B(n_5277),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_8138),
.B(n_8273),
.Y(n_8441)
);

AND2x2_ASAP7_75t_SL g8442 ( 
.A(n_8210),
.B(n_5362),
.Y(n_8442)
);

OAI21xp33_ASAP7_75t_SL g8443 ( 
.A1(n_8268),
.A2(n_5298),
.B(n_5287),
.Y(n_8443)
);

INVx2_ASAP7_75t_L g8444 ( 
.A(n_8164),
.Y(n_8444)
);

OAI332xp33_ASAP7_75t_L g8445 ( 
.A1(n_8127),
.A2(n_5456),
.A3(n_5457),
.B1(n_5294),
.B2(n_5289),
.B3(n_5277),
.C1(n_5295),
.C2(n_5285),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_8314),
.Y(n_8446)
);

AND2x2_ASAP7_75t_L g8447 ( 
.A(n_8099),
.B(n_8145),
.Y(n_8447)
);

INVx2_ASAP7_75t_SL g8448 ( 
.A(n_8225),
.Y(n_8448)
);

INVx2_ASAP7_75t_L g8449 ( 
.A(n_8313),
.Y(n_8449)
);

INVx1_ASAP7_75t_L g8450 ( 
.A(n_8314),
.Y(n_8450)
);

INVxp67_ASAP7_75t_SL g8451 ( 
.A(n_8121),
.Y(n_8451)
);

NAND2xp5_ASAP7_75t_L g8452 ( 
.A(n_8313),
.B(n_8289),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_8318),
.Y(n_8453)
);

AOI32xp33_ASAP7_75t_L g8454 ( 
.A1(n_8260),
.A2(n_5287),
.A3(n_5298),
.B1(n_5294),
.B2(n_5289),
.Y(n_8454)
);

INVxp67_ASAP7_75t_L g8455 ( 
.A(n_8147),
.Y(n_8455)
);

INVx1_ASAP7_75t_L g8456 ( 
.A(n_8318),
.Y(n_8456)
);

AND2x2_ASAP7_75t_L g8457 ( 
.A(n_8117),
.B(n_4789),
.Y(n_8457)
);

NAND4xp25_ASAP7_75t_L g8458 ( 
.A(n_8114),
.B(n_4391),
.C(n_4400),
.D(n_4372),
.Y(n_8458)
);

OAI32xp33_ASAP7_75t_L g8459 ( 
.A1(n_8125),
.A2(n_5298),
.A3(n_5295),
.B1(n_5285),
.B2(n_5457),
.Y(n_8459)
);

OAI21xp33_ASAP7_75t_L g8460 ( 
.A1(n_8237),
.A2(n_5298),
.B(n_4818),
.Y(n_8460)
);

INVx2_ASAP7_75t_SL g8461 ( 
.A(n_8139),
.Y(n_8461)
);

NOR2x1_ASAP7_75t_R g8462 ( 
.A(n_8325),
.B(n_4789),
.Y(n_8462)
);

INVx1_ASAP7_75t_L g8463 ( 
.A(n_8322),
.Y(n_8463)
);

AOI32xp33_ASAP7_75t_L g8464 ( 
.A1(n_8281),
.A2(n_5896),
.A3(n_5443),
.B1(n_6001),
.B2(n_5947),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_8322),
.Y(n_8465)
);

NOR2xp33_ASAP7_75t_L g8466 ( 
.A(n_8167),
.B(n_4818),
.Y(n_8466)
);

O2A1O1Ixp5_ASAP7_75t_L g8467 ( 
.A1(n_8178),
.A2(n_5385),
.B(n_5392),
.C(n_5387),
.Y(n_8467)
);

INVx1_ASAP7_75t_L g8468 ( 
.A(n_8090),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_8090),
.Y(n_8469)
);

INVx2_ASAP7_75t_L g8470 ( 
.A(n_8196),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_8324),
.Y(n_8471)
);

AND2x2_ASAP7_75t_L g8472 ( 
.A(n_8104),
.B(n_4818),
.Y(n_8472)
);

OAI21xp5_ASAP7_75t_L g8473 ( 
.A1(n_8251),
.A2(n_5896),
.B(n_5927),
.Y(n_8473)
);

OAI22xp33_ASAP7_75t_L g8474 ( 
.A1(n_8268),
.A2(n_5335),
.B1(n_5329),
.B2(n_5633),
.Y(n_8474)
);

NAND2xp5_ASAP7_75t_L g8475 ( 
.A(n_8200),
.B(n_8204),
.Y(n_8475)
);

INVx1_ASAP7_75t_L g8476 ( 
.A(n_8324),
.Y(n_8476)
);

INVx2_ASAP7_75t_L g8477 ( 
.A(n_8229),
.Y(n_8477)
);

INVx1_ASAP7_75t_L g8478 ( 
.A(n_8327),
.Y(n_8478)
);

AOI21xp5_ASAP7_75t_L g8479 ( 
.A1(n_8332),
.A2(n_5392),
.B(n_5387),
.Y(n_8479)
);

INVx1_ASAP7_75t_L g8480 ( 
.A(n_8327),
.Y(n_8480)
);

INVxp67_ASAP7_75t_L g8481 ( 
.A(n_8219),
.Y(n_8481)
);

OAI21xp33_ASAP7_75t_SL g8482 ( 
.A1(n_8135),
.A2(n_5734),
.B(n_5727),
.Y(n_8482)
);

NAND2xp5_ASAP7_75t_L g8483 ( 
.A(n_8200),
.B(n_5403),
.Y(n_8483)
);

INVx1_ASAP7_75t_L g8484 ( 
.A(n_8209),
.Y(n_8484)
);

INVx1_ASAP7_75t_L g8485 ( 
.A(n_8221),
.Y(n_8485)
);

AOI32xp33_ASAP7_75t_L g8486 ( 
.A1(n_8111),
.A2(n_5443),
.A3(n_6001),
.B1(n_5947),
.B2(n_5927),
.Y(n_8486)
);

HB1xp67_ASAP7_75t_L g8487 ( 
.A(n_8150),
.Y(n_8487)
);

OAI21xp33_ASAP7_75t_SL g8488 ( 
.A1(n_8115),
.A2(n_5734),
.B(n_5406),
.Y(n_8488)
);

NAND2xp33_ASAP7_75t_L g8489 ( 
.A(n_8152),
.B(n_4818),
.Y(n_8489)
);

OR2x2_ASAP7_75t_L g8490 ( 
.A(n_8224),
.B(n_8206),
.Y(n_8490)
);

OR2x2_ASAP7_75t_L g8491 ( 
.A(n_8227),
.B(n_5403),
.Y(n_8491)
);

NAND2x2_ASAP7_75t_L g8492 ( 
.A(n_8102),
.B(n_4403),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_8233),
.Y(n_8493)
);

INVx1_ASAP7_75t_SL g8494 ( 
.A(n_8194),
.Y(n_8494)
);

OR2x2_ASAP7_75t_L g8495 ( 
.A(n_8261),
.B(n_5406),
.Y(n_8495)
);

INVx1_ASAP7_75t_L g8496 ( 
.A(n_8134),
.Y(n_8496)
);

NAND2xp5_ASAP7_75t_L g8497 ( 
.A(n_8204),
.B(n_5409),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_8197),
.Y(n_8498)
);

INVx2_ASAP7_75t_L g8499 ( 
.A(n_8230),
.Y(n_8499)
);

INVx1_ASAP7_75t_SL g8500 ( 
.A(n_8168),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_8205),
.Y(n_8501)
);

INVx1_ASAP7_75t_L g8502 ( 
.A(n_8202),
.Y(n_8502)
);

AOI22xp5_ASAP7_75t_L g8503 ( 
.A1(n_8192),
.A2(n_5299),
.B1(n_5309),
.B2(n_5306),
.Y(n_8503)
);

AOI22xp5_ASAP7_75t_L g8504 ( 
.A1(n_8239),
.A2(n_5299),
.B1(n_5309),
.B2(n_5306),
.Y(n_8504)
);

NAND2x1p5_ASAP7_75t_L g8505 ( 
.A(n_8308),
.B(n_4818),
.Y(n_8505)
);

INVx1_ASAP7_75t_L g8506 ( 
.A(n_8203),
.Y(n_8506)
);

INVxp67_ASAP7_75t_SL g8507 ( 
.A(n_8208),
.Y(n_8507)
);

INVx1_ASAP7_75t_L g8508 ( 
.A(n_8199),
.Y(n_8508)
);

INVx2_ASAP7_75t_SL g8509 ( 
.A(n_8234),
.Y(n_8509)
);

NAND2x1p5_ASAP7_75t_L g8510 ( 
.A(n_8325),
.B(n_4818),
.Y(n_8510)
);

INVxp67_ASAP7_75t_SL g8511 ( 
.A(n_8258),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8248),
.Y(n_8512)
);

INVx1_ASAP7_75t_L g8513 ( 
.A(n_8180),
.Y(n_8513)
);

AOI22xp5_ASAP7_75t_L g8514 ( 
.A1(n_8240),
.A2(n_5312),
.B1(n_5316),
.B2(n_5314),
.Y(n_8514)
);

AOI21xp33_ASAP7_75t_SL g8515 ( 
.A1(n_8263),
.A2(n_5725),
.B(n_5461),
.Y(n_8515)
);

OAI32xp33_ASAP7_75t_L g8516 ( 
.A1(n_8262),
.A2(n_5461),
.A3(n_5316),
.B1(n_5334),
.B2(n_5314),
.Y(n_8516)
);

INVx1_ASAP7_75t_L g8517 ( 
.A(n_8244),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_8157),
.Y(n_8518)
);

INVx1_ASAP7_75t_L g8519 ( 
.A(n_8329),
.Y(n_8519)
);

BUFx2_ASAP7_75t_L g8520 ( 
.A(n_8179),
.Y(n_8520)
);

INVx2_ASAP7_75t_L g8521 ( 
.A(n_8243),
.Y(n_8521)
);

INVx2_ASAP7_75t_SL g8522 ( 
.A(n_8271),
.Y(n_8522)
);

AOI22xp5_ASAP7_75t_L g8523 ( 
.A1(n_8246),
.A2(n_5312),
.B1(n_5336),
.B2(n_5334),
.Y(n_8523)
);

INVx1_ASAP7_75t_L g8524 ( 
.A(n_8301),
.Y(n_8524)
);

AOI22xp5_ASAP7_75t_L g8525 ( 
.A1(n_8149),
.A2(n_5340),
.B1(n_5343),
.B2(n_5336),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_8282),
.Y(n_8526)
);

OAI21xp33_ASAP7_75t_L g8527 ( 
.A1(n_8267),
.A2(n_4862),
.B(n_4854),
.Y(n_8527)
);

BUFx2_ASAP7_75t_L g8528 ( 
.A(n_8247),
.Y(n_8528)
);

AOI32xp33_ASAP7_75t_L g8529 ( 
.A1(n_8323),
.A2(n_6031),
.A3(n_6134),
.B1(n_6108),
.B2(n_5240),
.Y(n_8529)
);

NAND2xp5_ASAP7_75t_L g8530 ( 
.A(n_8291),
.B(n_5409),
.Y(n_8530)
);

INVx1_ASAP7_75t_L g8531 ( 
.A(n_8282),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_8270),
.Y(n_8532)
);

NAND2xp5_ASAP7_75t_L g8533 ( 
.A(n_8333),
.B(n_5424),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_L g8534 ( 
.A(n_8297),
.B(n_5424),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_8299),
.B(n_5426),
.Y(n_8535)
);

INVx2_ASAP7_75t_L g8536 ( 
.A(n_8330),
.Y(n_8536)
);

OAI21xp33_ASAP7_75t_L g8537 ( 
.A1(n_8254),
.A2(n_4862),
.B(n_4854),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_8284),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_8284),
.Y(n_8539)
);

AND2x2_ASAP7_75t_L g8540 ( 
.A(n_8218),
.B(n_4854),
.Y(n_8540)
);

OR2x2_ASAP7_75t_L g8541 ( 
.A(n_8215),
.B(n_5426),
.Y(n_8541)
);

INVx2_ASAP7_75t_L g8542 ( 
.A(n_8303),
.Y(n_8542)
);

INVx2_ASAP7_75t_L g8543 ( 
.A(n_8312),
.Y(n_8543)
);

AND2x2_ASAP7_75t_L g8544 ( 
.A(n_8296),
.B(n_4854),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_8093),
.Y(n_8545)
);

INVx1_ASAP7_75t_L g8546 ( 
.A(n_8093),
.Y(n_8546)
);

OR2x2_ASAP7_75t_L g8547 ( 
.A(n_8193),
.B(n_5432),
.Y(n_8547)
);

OAI21xp33_ASAP7_75t_L g8548 ( 
.A1(n_8280),
.A2(n_4862),
.B(n_4854),
.Y(n_8548)
);

AND2x2_ASAP7_75t_L g8549 ( 
.A(n_8319),
.B(n_4854),
.Y(n_8549)
);

INVx1_ASAP7_75t_L g8550 ( 
.A(n_8264),
.Y(n_8550)
);

A2O1A1Ixp33_ASAP7_75t_L g8551 ( 
.A1(n_8118),
.A2(n_6108),
.B(n_6134),
.C(n_6031),
.Y(n_8551)
);

INVx1_ASAP7_75t_L g8552 ( 
.A(n_8265),
.Y(n_8552)
);

NAND3xp33_ASAP7_75t_L g8553 ( 
.A(n_8185),
.B(n_4897),
.C(n_4862),
.Y(n_8553)
);

NAND2xp5_ASAP7_75t_L g8554 ( 
.A(n_8207),
.B(n_5432),
.Y(n_8554)
);

OA21x2_ASAP7_75t_L g8555 ( 
.A1(n_8142),
.A2(n_5240),
.B(n_5135),
.Y(n_8555)
);

INVx1_ASAP7_75t_L g8556 ( 
.A(n_8217),
.Y(n_8556)
);

NAND3xp33_ASAP7_75t_L g8557 ( 
.A(n_8336),
.B(n_4981),
.C(n_4897),
.Y(n_8557)
);

INVx1_ASAP7_75t_L g8558 ( 
.A(n_8187),
.Y(n_8558)
);

AOI21xp5_ASAP7_75t_L g8559 ( 
.A1(n_8309),
.A2(n_5435),
.B(n_5434),
.Y(n_8559)
);

OAI22xp5_ASAP7_75t_L g8560 ( 
.A1(n_8191),
.A2(n_5435),
.B1(n_5439),
.B2(n_5434),
.Y(n_8560)
);

HB1xp67_ASAP7_75t_L g8561 ( 
.A(n_8252),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_8148),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_8189),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_8231),
.Y(n_8564)
);

BUFx3_ASAP7_75t_L g8565 ( 
.A(n_8341),
.Y(n_8565)
);

AND2x4_ASAP7_75t_L g8566 ( 
.A(n_8359),
.B(n_8315),
.Y(n_8566)
);

BUFx6f_ASAP7_75t_L g8567 ( 
.A(n_8359),
.Y(n_8567)
);

NAND2xp5_ASAP7_75t_L g8568 ( 
.A(n_8401),
.B(n_8300),
.Y(n_8568)
);

NAND2xp5_ASAP7_75t_L g8569 ( 
.A(n_8487),
.B(n_8250),
.Y(n_8569)
);

NAND2xp5_ASAP7_75t_L g8570 ( 
.A(n_8351),
.B(n_8376),
.Y(n_8570)
);

INVxp67_ASAP7_75t_L g8571 ( 
.A(n_8462),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_8375),
.Y(n_8572)
);

NOR2x1_ASAP7_75t_L g8573 ( 
.A(n_8400),
.B(n_8171),
.Y(n_8573)
);

NAND2xp5_ASAP7_75t_L g8574 ( 
.A(n_8511),
.B(n_8259),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_8398),
.Y(n_8575)
);

AND2x2_ASAP7_75t_L g8576 ( 
.A(n_8447),
.B(n_8339),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_8400),
.Y(n_8577)
);

NAND2xp5_ASAP7_75t_L g8578 ( 
.A(n_8407),
.B(n_8285),
.Y(n_8578)
);

NAND3xp33_ASAP7_75t_SL g8579 ( 
.A(n_8361),
.B(n_8162),
.C(n_8156),
.Y(n_8579)
);

INVxp67_ASAP7_75t_L g8580 ( 
.A(n_8520),
.Y(n_8580)
);

INVx2_ASAP7_75t_L g8581 ( 
.A(n_8510),
.Y(n_8581)
);

NAND2xp5_ASAP7_75t_L g8582 ( 
.A(n_8371),
.B(n_8328),
.Y(n_8582)
);

CKINVDCx14_ASAP7_75t_R g8583 ( 
.A(n_8346),
.Y(n_8583)
);

INVx2_ASAP7_75t_SL g8584 ( 
.A(n_8472),
.Y(n_8584)
);

NAND2x1_ASAP7_75t_L g8585 ( 
.A(n_8374),
.B(n_8235),
.Y(n_8585)
);

AND2x2_ASAP7_75t_L g8586 ( 
.A(n_8457),
.B(n_8253),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_8452),
.Y(n_8587)
);

INVx1_ASAP7_75t_L g8588 ( 
.A(n_8441),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_8505),
.Y(n_8589)
);

INVx2_ASAP7_75t_L g8590 ( 
.A(n_8430),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_8507),
.Y(n_8591)
);

INVx2_ASAP7_75t_SL g8592 ( 
.A(n_8449),
.Y(n_8592)
);

AND2x2_ASAP7_75t_L g8593 ( 
.A(n_8350),
.B(n_8331),
.Y(n_8593)
);

INVx2_ASAP7_75t_L g8594 ( 
.A(n_8416),
.Y(n_8594)
);

INVx2_ASAP7_75t_L g8595 ( 
.A(n_8442),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_8475),
.Y(n_8596)
);

INVx1_ASAP7_75t_SL g8597 ( 
.A(n_8349),
.Y(n_8597)
);

INVx2_ASAP7_75t_L g8598 ( 
.A(n_8355),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_8408),
.Y(n_8599)
);

NAND2xp5_ASAP7_75t_SL g8600 ( 
.A(n_8404),
.B(n_8276),
.Y(n_8600)
);

NAND3xp33_ASAP7_75t_L g8601 ( 
.A(n_8385),
.B(n_8256),
.C(n_8255),
.Y(n_8601)
);

NAND2xp5_ASAP7_75t_L g8602 ( 
.A(n_8451),
.B(n_8334),
.Y(n_8602)
);

INVx2_ASAP7_75t_L g8603 ( 
.A(n_8490),
.Y(n_8603)
);

OR2x2_ASAP7_75t_L g8604 ( 
.A(n_8377),
.B(n_8321),
.Y(n_8604)
);

INVx3_ASAP7_75t_L g8605 ( 
.A(n_8429),
.Y(n_8605)
);

INVx1_ASAP7_75t_L g8606 ( 
.A(n_8347),
.Y(n_8606)
);

AND2x2_ASAP7_75t_L g8607 ( 
.A(n_8396),
.B(n_8494),
.Y(n_8607)
);

NOR2xp33_ASAP7_75t_L g8608 ( 
.A(n_8481),
.B(n_8211),
.Y(n_8608)
);

BUFx3_ASAP7_75t_L g8609 ( 
.A(n_8528),
.Y(n_8609)
);

NAND3xp33_ASAP7_75t_L g8610 ( 
.A(n_8389),
.B(n_8257),
.C(n_8173),
.Y(n_8610)
);

OR2x2_ASAP7_75t_L g8611 ( 
.A(n_8393),
.B(n_8279),
.Y(n_8611)
);

AND2x4_ASAP7_75t_L g8612 ( 
.A(n_8390),
.B(n_8286),
.Y(n_8612)
);

BUFx3_ASAP7_75t_L g8613 ( 
.A(n_8417),
.Y(n_8613)
);

INVxp67_ASAP7_75t_L g8614 ( 
.A(n_8561),
.Y(n_8614)
);

AOI22xp33_ASAP7_75t_L g8615 ( 
.A1(n_8367),
.A2(n_8177),
.B1(n_8172),
.B2(n_8310),
.Y(n_8615)
);

INVx1_ASAP7_75t_SL g8616 ( 
.A(n_8397),
.Y(n_8616)
);

OAI22xp5_ASAP7_75t_L g8617 ( 
.A1(n_8492),
.A2(n_8295),
.B1(n_8320),
.B2(n_8306),
.Y(n_8617)
);

AND2x2_ASAP7_75t_L g8618 ( 
.A(n_8500),
.B(n_8311),
.Y(n_8618)
);

NAND2xp5_ASAP7_75t_L g8619 ( 
.A(n_8461),
.B(n_8409),
.Y(n_8619)
);

AND2x2_ASAP7_75t_L g8620 ( 
.A(n_8522),
.B(n_8304),
.Y(n_8620)
);

INVxp33_ASAP7_75t_SL g8621 ( 
.A(n_8353),
.Y(n_8621)
);

AOI22xp5_ASAP7_75t_L g8622 ( 
.A1(n_8343),
.A2(n_8238),
.B1(n_8245),
.B2(n_8288),
.Y(n_8622)
);

AOI22xp5_ASAP7_75t_L g8623 ( 
.A1(n_8406),
.A2(n_5343),
.B1(n_5340),
.B2(n_6006),
.Y(n_8623)
);

INVx1_ASAP7_75t_L g8624 ( 
.A(n_8364),
.Y(n_8624)
);

OR2x2_ASAP7_75t_L g8625 ( 
.A(n_8388),
.B(n_5439),
.Y(n_8625)
);

NAND2xp5_ASAP7_75t_L g8626 ( 
.A(n_8498),
.B(n_5441),
.Y(n_8626)
);

INVxp67_ASAP7_75t_L g8627 ( 
.A(n_8426),
.Y(n_8627)
);

INVx2_ASAP7_75t_L g8628 ( 
.A(n_8365),
.Y(n_8628)
);

AND2x2_ASAP7_75t_L g8629 ( 
.A(n_8352),
.B(n_4897),
.Y(n_8629)
);

INVx3_ASAP7_75t_SL g8630 ( 
.A(n_8342),
.Y(n_8630)
);

INVx1_ASAP7_75t_SL g8631 ( 
.A(n_8386),
.Y(n_8631)
);

INVxp67_ASAP7_75t_L g8632 ( 
.A(n_8413),
.Y(n_8632)
);

INVx3_ASAP7_75t_L g8633 ( 
.A(n_8429),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_8420),
.Y(n_8634)
);

BUFx3_ASAP7_75t_L g8635 ( 
.A(n_8512),
.Y(n_8635)
);

AND2x4_ASAP7_75t_SL g8636 ( 
.A(n_8470),
.B(n_4897),
.Y(n_8636)
);

INVx2_ASAP7_75t_SL g8637 ( 
.A(n_8412),
.Y(n_8637)
);

HB1xp67_ASAP7_75t_L g8638 ( 
.A(n_8526),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_8531),
.Y(n_8639)
);

NAND2xp5_ASAP7_75t_L g8640 ( 
.A(n_8373),
.B(n_5441),
.Y(n_8640)
);

AND2x2_ASAP7_75t_L g8641 ( 
.A(n_8427),
.B(n_4897),
.Y(n_8641)
);

AND2x2_ASAP7_75t_L g8642 ( 
.A(n_8434),
.B(n_4897),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_8366),
.Y(n_8643)
);

NAND2xp5_ASAP7_75t_L g8644 ( 
.A(n_8410),
.B(n_5448),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_L g8645 ( 
.A(n_8519),
.B(n_5448),
.Y(n_8645)
);

BUFx3_ASAP7_75t_L g8646 ( 
.A(n_8484),
.Y(n_8646)
);

AND2x2_ASAP7_75t_L g8647 ( 
.A(n_8437),
.B(n_4981),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_8340),
.Y(n_8648)
);

BUFx2_ASAP7_75t_L g8649 ( 
.A(n_8399),
.Y(n_8649)
);

INVx4_ASAP7_75t_L g8650 ( 
.A(n_8381),
.Y(n_8650)
);

NAND2xp5_ASAP7_75t_L g8651 ( 
.A(n_8403),
.B(n_5460),
.Y(n_8651)
);

INVx1_ASAP7_75t_L g8652 ( 
.A(n_8538),
.Y(n_8652)
);

NAND2xp5_ASAP7_75t_L g8653 ( 
.A(n_8524),
.B(n_5460),
.Y(n_8653)
);

INVx2_ASAP7_75t_SL g8654 ( 
.A(n_8544),
.Y(n_8654)
);

OR2x2_ASAP7_75t_L g8655 ( 
.A(n_8344),
.B(n_5462),
.Y(n_8655)
);

AOI22xp33_ASAP7_75t_L g8656 ( 
.A1(n_8378),
.A2(n_6171),
.B1(n_6190),
.B2(n_6176),
.Y(n_8656)
);

AND2x2_ASAP7_75t_L g8657 ( 
.A(n_8477),
.B(n_4981),
.Y(n_8657)
);

INVx1_ASAP7_75t_SL g8658 ( 
.A(n_8402),
.Y(n_8658)
);

NOR2xp33_ASAP7_75t_L g8659 ( 
.A(n_8455),
.B(n_4981),
.Y(n_8659)
);

INVx1_ASAP7_75t_L g8660 ( 
.A(n_8539),
.Y(n_8660)
);

NAND2xp5_ASAP7_75t_L g8661 ( 
.A(n_8532),
.B(n_5462),
.Y(n_8661)
);

INVx1_ASAP7_75t_SL g8662 ( 
.A(n_8380),
.Y(n_8662)
);

OR2x2_ASAP7_75t_L g8663 ( 
.A(n_8485),
.B(n_5466),
.Y(n_8663)
);

AO21x1_ASAP7_75t_L g8664 ( 
.A1(n_8362),
.A2(n_5471),
.B(n_5466),
.Y(n_8664)
);

OR2x2_ASAP7_75t_L g8665 ( 
.A(n_8493),
.B(n_5471),
.Y(n_8665)
);

HB1xp67_ASAP7_75t_L g8666 ( 
.A(n_8499),
.Y(n_8666)
);

OR2x2_ASAP7_75t_L g8667 ( 
.A(n_8502),
.B(n_5477),
.Y(n_8667)
);

NAND2xp5_ASAP7_75t_L g8668 ( 
.A(n_8536),
.B(n_5477),
.Y(n_8668)
);

OR2x2_ASAP7_75t_L g8669 ( 
.A(n_8506),
.B(n_5481),
.Y(n_8669)
);

AOI22xp33_ASAP7_75t_L g8670 ( 
.A1(n_8338),
.A2(n_6171),
.B1(n_6190),
.B2(n_6176),
.Y(n_8670)
);

INVx1_ASAP7_75t_L g8671 ( 
.A(n_8431),
.Y(n_8671)
);

INVx1_ASAP7_75t_SL g8672 ( 
.A(n_8348),
.Y(n_8672)
);

AND2x2_ASAP7_75t_L g8673 ( 
.A(n_8444),
.B(n_8521),
.Y(n_8673)
);

AND2x2_ASAP7_75t_L g8674 ( 
.A(n_8394),
.B(n_4981),
.Y(n_8674)
);

AND2x2_ASAP7_75t_L g8675 ( 
.A(n_8542),
.B(n_4981),
.Y(n_8675)
);

AND2x2_ASAP7_75t_L g8676 ( 
.A(n_8543),
.B(n_5056),
.Y(n_8676)
);

AND3x1_ASAP7_75t_L g8677 ( 
.A(n_8379),
.B(n_4672),
.C(n_4638),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_8435),
.Y(n_8678)
);

INVx1_ASAP7_75t_SL g8679 ( 
.A(n_8440),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8549),
.Y(n_8680)
);

INVx2_ASAP7_75t_L g8681 ( 
.A(n_8419),
.Y(n_8681)
);

INVx1_ASAP7_75t_L g8682 ( 
.A(n_8446),
.Y(n_8682)
);

CKINVDCx16_ASAP7_75t_R g8683 ( 
.A(n_8387),
.Y(n_8683)
);

AND2x2_ASAP7_75t_L g8684 ( 
.A(n_8438),
.B(n_5056),
.Y(n_8684)
);

NOR2x1_ASAP7_75t_L g8685 ( 
.A(n_8450),
.B(n_5056),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_8453),
.Y(n_8686)
);

AOI21xp5_ASAP7_75t_L g8687 ( 
.A1(n_8356),
.A2(n_5483),
.B(n_5481),
.Y(n_8687)
);

INVx2_ASAP7_75t_L g8688 ( 
.A(n_8540),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_8340),
.Y(n_8689)
);

NAND2xp5_ASAP7_75t_L g8690 ( 
.A(n_8508),
.B(n_5483),
.Y(n_8690)
);

BUFx3_ASAP7_75t_L g8691 ( 
.A(n_8382),
.Y(n_8691)
);

OR2x2_ASAP7_75t_L g8692 ( 
.A(n_8423),
.B(n_5487),
.Y(n_8692)
);

NOR2x1_ASAP7_75t_L g8693 ( 
.A(n_8456),
.B(n_5056),
.Y(n_8693)
);

AND2x4_ASAP7_75t_L g8694 ( 
.A(n_8509),
.B(n_5056),
.Y(n_8694)
);

AND2x4_ASAP7_75t_L g8695 ( 
.A(n_8360),
.B(n_5056),
.Y(n_8695)
);

INVx2_ASAP7_75t_L g8696 ( 
.A(n_8463),
.Y(n_8696)
);

INVx1_ASAP7_75t_SL g8697 ( 
.A(n_8354),
.Y(n_8697)
);

NAND2xp5_ASAP7_75t_L g8698 ( 
.A(n_8558),
.B(n_5487),
.Y(n_8698)
);

HB1xp67_ASAP7_75t_L g8699 ( 
.A(n_8465),
.Y(n_8699)
);

INVx2_ASAP7_75t_L g8700 ( 
.A(n_8471),
.Y(n_8700)
);

AND2x2_ASAP7_75t_L g8701 ( 
.A(n_8448),
.B(n_5064),
.Y(n_8701)
);

AND2x2_ASAP7_75t_L g8702 ( 
.A(n_8337),
.B(n_5064),
.Y(n_8702)
);

NAND2xp5_ASAP7_75t_SL g8703 ( 
.A(n_8383),
.B(n_5064),
.Y(n_8703)
);

INVx1_ASAP7_75t_SL g8704 ( 
.A(n_8425),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_8476),
.Y(n_8705)
);

AND2x2_ASAP7_75t_L g8706 ( 
.A(n_8415),
.B(n_5064),
.Y(n_8706)
);

AO21x2_ASAP7_75t_L g8707 ( 
.A1(n_8391),
.A2(n_5953),
.B(n_5935),
.Y(n_8707)
);

INVx2_ASAP7_75t_L g8708 ( 
.A(n_8478),
.Y(n_8708)
);

INVx2_ASAP7_75t_L g8709 ( 
.A(n_8480),
.Y(n_8709)
);

INVx2_ASAP7_75t_L g8710 ( 
.A(n_8491),
.Y(n_8710)
);

NAND2xp5_ASAP7_75t_SL g8711 ( 
.A(n_8372),
.B(n_5064),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8468),
.Y(n_8712)
);

INVx1_ASAP7_75t_SL g8713 ( 
.A(n_8513),
.Y(n_8713)
);

AND2x2_ASAP7_75t_L g8714 ( 
.A(n_8384),
.B(n_5064),
.Y(n_8714)
);

INVx2_ASAP7_75t_SL g8715 ( 
.A(n_8357),
.Y(n_8715)
);

INVx1_ASAP7_75t_L g8716 ( 
.A(n_8468),
.Y(n_8716)
);

OR2x6_ASAP7_75t_L g8717 ( 
.A(n_8395),
.B(n_8411),
.Y(n_8717)
);

INVx1_ASAP7_75t_L g8718 ( 
.A(n_8469),
.Y(n_8718)
);

INVx1_ASAP7_75t_SL g8719 ( 
.A(n_8489),
.Y(n_8719)
);

INVx2_ASAP7_75t_L g8720 ( 
.A(n_8495),
.Y(n_8720)
);

AND2x2_ASAP7_75t_L g8721 ( 
.A(n_8370),
.B(n_5069),
.Y(n_8721)
);

INVx1_ASAP7_75t_L g8722 ( 
.A(n_8469),
.Y(n_8722)
);

AND2x2_ASAP7_75t_L g8723 ( 
.A(n_8517),
.B(n_5069),
.Y(n_8723)
);

HB1xp67_ASAP7_75t_L g8724 ( 
.A(n_8439),
.Y(n_8724)
);

INVx2_ASAP7_75t_L g8725 ( 
.A(n_8547),
.Y(n_8725)
);

INVxp67_ASAP7_75t_L g8726 ( 
.A(n_8550),
.Y(n_8726)
);

AND2x2_ASAP7_75t_L g8727 ( 
.A(n_8405),
.B(n_5069),
.Y(n_8727)
);

OR2x2_ASAP7_75t_L g8728 ( 
.A(n_8433),
.B(n_5488),
.Y(n_8728)
);

INVx1_ASAP7_75t_L g8729 ( 
.A(n_8345),
.Y(n_8729)
);

HB1xp67_ASAP7_75t_L g8730 ( 
.A(n_8545),
.Y(n_8730)
);

INVx2_ASAP7_75t_L g8731 ( 
.A(n_8467),
.Y(n_8731)
);

INVx1_ASAP7_75t_L g8732 ( 
.A(n_8546),
.Y(n_8732)
);

AND2x2_ASAP7_75t_L g8733 ( 
.A(n_8414),
.B(n_5069),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8358),
.Y(n_8734)
);

CKINVDCx16_ASAP7_75t_R g8735 ( 
.A(n_8501),
.Y(n_8735)
);

AND3x1_ASAP7_75t_L g8736 ( 
.A(n_8552),
.B(n_8460),
.C(n_8556),
.Y(n_8736)
);

INVx3_ASAP7_75t_SL g8737 ( 
.A(n_8563),
.Y(n_8737)
);

NOR2xp33_ASAP7_75t_L g8738 ( 
.A(n_8564),
.B(n_5069),
.Y(n_8738)
);

INVx1_ASAP7_75t_L g8739 ( 
.A(n_8483),
.Y(n_8739)
);

AOI22xp33_ASAP7_75t_L g8740 ( 
.A1(n_8473),
.A2(n_8421),
.B1(n_8424),
.B2(n_8496),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_L g8741 ( 
.A(n_8518),
.B(n_8392),
.Y(n_8741)
);

HB1xp67_ASAP7_75t_L g8742 ( 
.A(n_8562),
.Y(n_8742)
);

INVx1_ASAP7_75t_SL g8743 ( 
.A(n_8554),
.Y(n_8743)
);

CKINVDCx16_ASAP7_75t_R g8744 ( 
.A(n_8418),
.Y(n_8744)
);

INVxp67_ASAP7_75t_SL g8745 ( 
.A(n_8562),
.Y(n_8745)
);

INVx2_ASAP7_75t_L g8746 ( 
.A(n_8541),
.Y(n_8746)
);

AND2x4_ASAP7_75t_L g8747 ( 
.A(n_8428),
.B(n_5069),
.Y(n_8747)
);

AND2x2_ASAP7_75t_L g8748 ( 
.A(n_8515),
.B(n_5488),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_8555),
.Y(n_8749)
);

NAND2xp5_ASAP7_75t_L g8750 ( 
.A(n_8534),
.B(n_5490),
.Y(n_8750)
);

AOI22xp5_ASAP7_75t_L g8751 ( 
.A1(n_8488),
.A2(n_6055),
.B1(n_6091),
.B2(n_6006),
.Y(n_8751)
);

NAND2xp5_ASAP7_75t_L g8752 ( 
.A(n_8576),
.B(n_8533),
.Y(n_8752)
);

OAI31xp33_ASAP7_75t_L g8753 ( 
.A1(n_8600),
.A2(n_8551),
.A3(n_8560),
.B(n_8368),
.Y(n_8753)
);

INVxp33_ASAP7_75t_L g8754 ( 
.A(n_8666),
.Y(n_8754)
);

NAND2x1_ASAP7_75t_L g8755 ( 
.A(n_8650),
.B(n_8557),
.Y(n_8755)
);

AND2x2_ASAP7_75t_L g8756 ( 
.A(n_8607),
.B(n_8466),
.Y(n_8756)
);

OAI321xp33_ASAP7_75t_L g8757 ( 
.A1(n_8572),
.A2(n_8454),
.A3(n_8464),
.B1(n_8486),
.B2(n_8529),
.C(n_8553),
.Y(n_8757)
);

AOI21xp5_ASAP7_75t_L g8758 ( 
.A1(n_8572),
.A2(n_8459),
.B(n_8497),
.Y(n_8758)
);

INVxp67_ASAP7_75t_SL g8759 ( 
.A(n_8567),
.Y(n_8759)
);

INVx1_ASAP7_75t_SL g8760 ( 
.A(n_8658),
.Y(n_8760)
);

NAND3xp33_ASAP7_75t_L g8761 ( 
.A(n_8583),
.B(n_8369),
.C(n_8363),
.Y(n_8761)
);

NAND2xp5_ASAP7_75t_SL g8762 ( 
.A(n_8567),
.B(n_8443),
.Y(n_8762)
);

AOI32xp33_ASAP7_75t_L g8763 ( 
.A1(n_8643),
.A2(n_8482),
.A3(n_8530),
.B1(n_8535),
.B2(n_8537),
.Y(n_8763)
);

NAND2xp5_ASAP7_75t_L g8764 ( 
.A(n_8567),
.B(n_8559),
.Y(n_8764)
);

AND2x2_ASAP7_75t_L g8765 ( 
.A(n_8609),
.B(n_8527),
.Y(n_8765)
);

OR2x2_ASAP7_75t_L g8766 ( 
.A(n_8616),
.B(n_8458),
.Y(n_8766)
);

NAND2xp5_ASAP7_75t_L g8767 ( 
.A(n_8597),
.B(n_8445),
.Y(n_8767)
);

INVx1_ASAP7_75t_L g8768 ( 
.A(n_8724),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_8649),
.Y(n_8769)
);

AOI22xp5_ASAP7_75t_SL g8770 ( 
.A1(n_8621),
.A2(n_8555),
.B1(n_8436),
.B2(n_8479),
.Y(n_8770)
);

INVx1_ASAP7_75t_L g8771 ( 
.A(n_8742),
.Y(n_8771)
);

NAND2xp5_ASAP7_75t_L g8772 ( 
.A(n_8631),
.B(n_8504),
.Y(n_8772)
);

NAND2xp5_ASAP7_75t_L g8773 ( 
.A(n_8662),
.B(n_8566),
.Y(n_8773)
);

INVx3_ASAP7_75t_L g8774 ( 
.A(n_8565),
.Y(n_8774)
);

AOI31xp33_ASAP7_75t_L g8775 ( 
.A1(n_8580),
.A2(n_8548),
.A3(n_8432),
.B(n_8474),
.Y(n_8775)
);

AOI22xp33_ASAP7_75t_L g8776 ( 
.A1(n_8579),
.A2(n_8523),
.B1(n_8525),
.B2(n_8503),
.Y(n_8776)
);

OAI22xp5_ASAP7_75t_L g8777 ( 
.A1(n_8614),
.A2(n_8672),
.B1(n_8735),
.B2(n_8603),
.Y(n_8777)
);

AND2x2_ASAP7_75t_L g8778 ( 
.A(n_8673),
.B(n_8459),
.Y(n_8778)
);

OAI21xp33_ASAP7_75t_SL g8779 ( 
.A1(n_8643),
.A2(n_8514),
.B(n_8422),
.Y(n_8779)
);

O2A1O1Ixp33_ASAP7_75t_SL g8780 ( 
.A1(n_8711),
.A2(n_8422),
.B(n_8516),
.C(n_5493),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_8566),
.Y(n_8781)
);

OAI33xp33_ASAP7_75t_L g8782 ( 
.A1(n_8617),
.A2(n_8516),
.A3(n_5497),
.B1(n_5493),
.B2(n_5498),
.B3(n_5496),
.Y(n_8782)
);

INVx2_ASAP7_75t_L g8783 ( 
.A(n_8611),
.Y(n_8783)
);

NAND2xp5_ASAP7_75t_L g8784 ( 
.A(n_8697),
.B(n_5490),
.Y(n_8784)
);

INVx1_ASAP7_75t_L g8785 ( 
.A(n_8730),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_8745),
.Y(n_8786)
);

INVx2_ASAP7_75t_SL g8787 ( 
.A(n_8613),
.Y(n_8787)
);

INVx2_ASAP7_75t_L g8788 ( 
.A(n_8628),
.Y(n_8788)
);

INVx2_ASAP7_75t_SL g8789 ( 
.A(n_8691),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_8630),
.B(n_5496),
.Y(n_8790)
);

NOR2xp33_ASAP7_75t_L g8791 ( 
.A(n_8650),
.B(n_5991),
.Y(n_8791)
);

NAND2x1p5_ASAP7_75t_L g8792 ( 
.A(n_8635),
.B(n_4391),
.Y(n_8792)
);

AND2x4_ASAP7_75t_L g8793 ( 
.A(n_8637),
.B(n_4400),
.Y(n_8793)
);

AOI21xp5_ASAP7_75t_SL g8794 ( 
.A1(n_8570),
.A2(n_4403),
.B(n_4400),
.Y(n_8794)
);

INVx1_ASAP7_75t_L g8795 ( 
.A(n_8573),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_8638),
.Y(n_8796)
);

INVx1_ASAP7_75t_L g8797 ( 
.A(n_8699),
.Y(n_8797)
);

INVx1_ASAP7_75t_L g8798 ( 
.A(n_8594),
.Y(n_8798)
);

INVx2_ASAP7_75t_L g8799 ( 
.A(n_8618),
.Y(n_8799)
);

OR2x2_ASAP7_75t_L g8800 ( 
.A(n_8619),
.B(n_5497),
.Y(n_8800)
);

NAND2xp5_ASAP7_75t_L g8801 ( 
.A(n_8683),
.B(n_5498),
.Y(n_8801)
);

OAI211xp5_ASAP7_75t_L g8802 ( 
.A1(n_8585),
.A2(n_4876),
.B(n_5725),
.C(n_4403),
.Y(n_8802)
);

INVx1_ASAP7_75t_L g8803 ( 
.A(n_8569),
.Y(n_8803)
);

NOR2xp33_ASAP7_75t_L g8804 ( 
.A(n_8737),
.B(n_5991),
.Y(n_8804)
);

A2O1A1Ixp33_ASAP7_75t_L g8805 ( 
.A1(n_8608),
.A2(n_5609),
.B(n_5614),
.C(n_5610),
.Y(n_8805)
);

AOI221xp5_ASAP7_75t_L g8806 ( 
.A1(n_8734),
.A2(n_8615),
.B1(n_8749),
.B2(n_8656),
.C(n_8670),
.Y(n_8806)
);

INVx1_ASAP7_75t_L g8807 ( 
.A(n_8577),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_8591),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_8679),
.B(n_5500),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8605),
.Y(n_8810)
);

INVx1_ASAP7_75t_L g8811 ( 
.A(n_8605),
.Y(n_8811)
);

AOI21xp5_ASAP7_75t_L g8812 ( 
.A1(n_8703),
.A2(n_5506),
.B(n_5500),
.Y(n_8812)
);

INVx1_ASAP7_75t_L g8813 ( 
.A(n_8633),
.Y(n_8813)
);

NOR2xp67_ASAP7_75t_L g8814 ( 
.A(n_8633),
.B(n_5506),
.Y(n_8814)
);

INVx2_ASAP7_75t_L g8815 ( 
.A(n_8604),
.Y(n_8815)
);

AOI21xp5_ASAP7_75t_L g8816 ( 
.A1(n_8578),
.A2(n_5513),
.B(n_5509),
.Y(n_8816)
);

INVx1_ASAP7_75t_L g8817 ( 
.A(n_8612),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8612),
.Y(n_8818)
);

NOR2xp33_ASAP7_75t_L g8819 ( 
.A(n_8744),
.B(n_5991),
.Y(n_8819)
);

AOI21xp5_ASAP7_75t_L g8820 ( 
.A1(n_8568),
.A2(n_5513),
.B(n_5509),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_8646),
.Y(n_8821)
);

AOI322xp5_ASAP7_75t_L g8822 ( 
.A1(n_8734),
.A2(n_5630),
.A3(n_5610),
.B1(n_5632),
.B2(n_5639),
.C1(n_5614),
.C2(n_5609),
.Y(n_8822)
);

INVxp33_ASAP7_75t_L g8823 ( 
.A(n_8574),
.Y(n_8823)
);

NAND2xp5_ASAP7_75t_L g8824 ( 
.A(n_8704),
.B(n_5516),
.Y(n_8824)
);

OR2x2_ASAP7_75t_L g8825 ( 
.A(n_8592),
.B(n_5516),
.Y(n_8825)
);

INVx1_ASAP7_75t_L g8826 ( 
.A(n_8602),
.Y(n_8826)
);

INVx1_ASAP7_75t_L g8827 ( 
.A(n_8588),
.Y(n_8827)
);

NAND3xp33_ASAP7_75t_L g8828 ( 
.A(n_8601),
.B(n_6158),
.C(n_6171),
.Y(n_8828)
);

AOI22xp5_ASAP7_75t_L g8829 ( 
.A1(n_8623),
.A2(n_6091),
.B1(n_6136),
.B2(n_6055),
.Y(n_8829)
);

A2O1A1Ixp33_ASAP7_75t_L g8830 ( 
.A1(n_8731),
.A2(n_5630),
.B(n_5639),
.C(n_5632),
.Y(n_8830)
);

OAI211xp5_ASAP7_75t_SL g8831 ( 
.A1(n_8571),
.A2(n_5096),
.B(n_5520),
.C(n_5519),
.Y(n_8831)
);

OAI22xp5_ASAP7_75t_L g8832 ( 
.A1(n_8632),
.A2(n_8713),
.B1(n_8719),
.B2(n_8598),
.Y(n_8832)
);

NAND2xp5_ASAP7_75t_L g8833 ( 
.A(n_8584),
.B(n_5519),
.Y(n_8833)
);

OR2x2_ASAP7_75t_L g8834 ( 
.A(n_8715),
.B(n_5520),
.Y(n_8834)
);

AOI22xp5_ASAP7_75t_L g8835 ( 
.A1(n_8595),
.A2(n_6136),
.B1(n_6151),
.B2(n_6091),
.Y(n_8835)
);

NAND2xp33_ASAP7_75t_L g8836 ( 
.A(n_8654),
.B(n_5725),
.Y(n_8836)
);

INVx1_ASAP7_75t_L g8837 ( 
.A(n_8712),
.Y(n_8837)
);

CKINVDCx16_ASAP7_75t_R g8838 ( 
.A(n_8593),
.Y(n_8838)
);

NAND2xp5_ASAP7_75t_L g8839 ( 
.A(n_8743),
.B(n_5521),
.Y(n_8839)
);

OR2x2_ASAP7_75t_L g8840 ( 
.A(n_8710),
.B(n_5521),
.Y(n_8840)
);

INVx1_ASAP7_75t_SL g8841 ( 
.A(n_8629),
.Y(n_8841)
);

INVx1_ASAP7_75t_L g8842 ( 
.A(n_8716),
.Y(n_8842)
);

INVx2_ASAP7_75t_L g8843 ( 
.A(n_8674),
.Y(n_8843)
);

OAI211xp5_ASAP7_75t_SL g8844 ( 
.A1(n_8726),
.A2(n_5526),
.B(n_5532),
.C(n_5525),
.Y(n_8844)
);

NAND2x1_ASAP7_75t_L g8845 ( 
.A(n_8685),
.B(n_5089),
.Y(n_8845)
);

NOR2xp33_ASAP7_75t_L g8846 ( 
.A(n_8681),
.B(n_6030),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_8718),
.Y(n_8847)
);

AOI22xp5_ASAP7_75t_L g8848 ( 
.A1(n_8575),
.A2(n_6151),
.B1(n_6136),
.B2(n_6158),
.Y(n_8848)
);

O2A1O1Ixp33_ASAP7_75t_L g8849 ( 
.A1(n_8606),
.A2(n_6045),
.B(n_6030),
.C(n_6176),
.Y(n_8849)
);

INVx2_ASAP7_75t_L g8850 ( 
.A(n_8586),
.Y(n_8850)
);

OR2x2_ASAP7_75t_L g8851 ( 
.A(n_8720),
.B(n_5525),
.Y(n_8851)
);

INVx2_ASAP7_75t_L g8852 ( 
.A(n_8725),
.Y(n_8852)
);

AND2x2_ASAP7_75t_L g8853 ( 
.A(n_8641),
.B(n_5480),
.Y(n_8853)
);

INVx1_ASAP7_75t_L g8854 ( 
.A(n_8722),
.Y(n_8854)
);

INVx2_ASAP7_75t_SL g8855 ( 
.A(n_8636),
.Y(n_8855)
);

NAND4xp25_ASAP7_75t_L g8856 ( 
.A(n_8622),
.B(n_5362),
.C(n_4741),
.D(n_4804),
.Y(n_8856)
);

AOI21xp5_ASAP7_75t_L g8857 ( 
.A1(n_8741),
.A2(n_5532),
.B(n_5526),
.Y(n_8857)
);

AOI21xp5_ASAP7_75t_L g8858 ( 
.A1(n_8693),
.A2(n_5547),
.B(n_5540),
.Y(n_8858)
);

AND2x2_ASAP7_75t_L g8859 ( 
.A(n_8642),
.B(n_5480),
.Y(n_8859)
);

AOI21xp33_ASAP7_75t_SL g8860 ( 
.A1(n_8610),
.A2(n_6045),
.B(n_6030),
.Y(n_8860)
);

NAND2xp5_ASAP7_75t_L g8861 ( 
.A(n_8747),
.B(n_5540),
.Y(n_8861)
);

INVx2_ASAP7_75t_L g8862 ( 
.A(n_8747),
.Y(n_8862)
);

OAI221xp5_ASAP7_75t_L g8863 ( 
.A1(n_8740),
.A2(n_6190),
.B1(n_6201),
.B2(n_6195),
.C(n_6045),
.Y(n_8863)
);

NAND2xp5_ASAP7_75t_L g8864 ( 
.A(n_8746),
.B(n_5547),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_8694),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_8620),
.Y(n_8866)
);

NAND2xp5_ASAP7_75t_L g8867 ( 
.A(n_8695),
.B(n_5555),
.Y(n_8867)
);

NAND2xp5_ASAP7_75t_L g8868 ( 
.A(n_8695),
.B(n_5555),
.Y(n_8868)
);

OAI22xp33_ASAP7_75t_L g8869 ( 
.A1(n_8751),
.A2(n_5335),
.B1(n_5329),
.B2(n_6195),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_8664),
.Y(n_8870)
);

NAND2xp5_ASAP7_75t_L g8871 ( 
.A(n_8727),
.B(n_5557),
.Y(n_8871)
);

AOI322xp5_ASAP7_75t_L g8872 ( 
.A1(n_8575),
.A2(n_5654),
.A3(n_5643),
.B1(n_5657),
.B2(n_5658),
.C1(n_5644),
.C2(n_5641),
.Y(n_8872)
);

INVx1_ASAP7_75t_SL g8873 ( 
.A(n_8706),
.Y(n_8873)
);

INVx1_ASAP7_75t_SL g8874 ( 
.A(n_8723),
.Y(n_8874)
);

NAND2xp5_ASAP7_75t_SL g8875 ( 
.A(n_8694),
.B(n_5362),
.Y(n_8875)
);

INVx1_ASAP7_75t_L g8876 ( 
.A(n_8732),
.Y(n_8876)
);

INVx2_ASAP7_75t_L g8877 ( 
.A(n_8647),
.Y(n_8877)
);

AND2x2_ASAP7_75t_L g8878 ( 
.A(n_8657),
.B(n_5480),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_8732),
.Y(n_8879)
);

NAND2xp5_ASAP7_75t_L g8880 ( 
.A(n_8675),
.B(n_5557),
.Y(n_8880)
);

NAND3xp33_ASAP7_75t_L g8881 ( 
.A(n_8599),
.B(n_6201),
.C(n_6195),
.Y(n_8881)
);

OAI221xp5_ASAP7_75t_L g8882 ( 
.A1(n_8599),
.A2(n_6201),
.B1(n_6068),
.B2(n_5335),
.C(n_5329),
.Y(n_8882)
);

INVxp67_ASAP7_75t_SL g8883 ( 
.A(n_8696),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_8648),
.Y(n_8884)
);

OAI22xp33_ASAP7_75t_L g8885 ( 
.A1(n_8634),
.A2(n_8606),
.B1(n_8705),
.B2(n_8700),
.Y(n_8885)
);

NAND2xp5_ASAP7_75t_L g8886 ( 
.A(n_8676),
.B(n_5562),
.Y(n_8886)
);

INVx1_ASAP7_75t_L g8887 ( 
.A(n_8648),
.Y(n_8887)
);

AND2x2_ASAP7_75t_L g8888 ( 
.A(n_8701),
.B(n_5480),
.Y(n_8888)
);

NAND2xp5_ASAP7_75t_L g8889 ( 
.A(n_8708),
.B(n_5562),
.Y(n_8889)
);

OAI22xp5_ASAP7_75t_L g8890 ( 
.A1(n_8587),
.A2(n_5590),
.B1(n_5635),
.B2(n_5569),
.Y(n_8890)
);

OAI22xp33_ASAP7_75t_L g8891 ( 
.A1(n_8709),
.A2(n_5335),
.B1(n_6068),
.B2(n_6207),
.Y(n_8891)
);

AOI22xp5_ASAP7_75t_L g8892 ( 
.A1(n_8596),
.A2(n_6151),
.B1(n_6153),
.B2(n_5953),
.Y(n_8892)
);

NOR2x1_ASAP7_75t_L g8893 ( 
.A(n_8689),
.B(n_5567),
.Y(n_8893)
);

AND2x2_ASAP7_75t_L g8894 ( 
.A(n_8688),
.B(n_5594),
.Y(n_8894)
);

AOI21xp5_ASAP7_75t_L g8895 ( 
.A1(n_8582),
.A2(n_5569),
.B(n_5567),
.Y(n_8895)
);

OR2x2_ASAP7_75t_L g8896 ( 
.A(n_8680),
.B(n_5570),
.Y(n_8896)
);

INVx1_ASAP7_75t_SL g8897 ( 
.A(n_8702),
.Y(n_8897)
);

NAND2xp5_ASAP7_75t_L g8898 ( 
.A(n_8624),
.B(n_8590),
.Y(n_8898)
);

OAI22xp33_ASAP7_75t_L g8899 ( 
.A1(n_8589),
.A2(n_6068),
.B1(n_6219),
.B2(n_6207),
.Y(n_8899)
);

AOI22xp33_ASAP7_75t_L g8900 ( 
.A1(n_8707),
.A2(n_5953),
.B1(n_5935),
.B2(n_6207),
.Y(n_8900)
);

INVx2_ASAP7_75t_L g8901 ( 
.A(n_8625),
.Y(n_8901)
);

INVx1_ASAP7_75t_SL g8902 ( 
.A(n_8733),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_L g8903 ( 
.A(n_8738),
.B(n_5570),
.Y(n_8903)
);

OAI22xp5_ASAP7_75t_L g8904 ( 
.A1(n_8736),
.A2(n_5627),
.B1(n_5664),
.B2(n_5581),
.Y(n_8904)
);

INVx1_ASAP7_75t_L g8905 ( 
.A(n_8689),
.Y(n_8905)
);

NOR3xp33_ASAP7_75t_L g8906 ( 
.A(n_8639),
.B(n_4670),
.C(n_4667),
.Y(n_8906)
);

NAND3xp33_ASAP7_75t_L g8907 ( 
.A(n_8652),
.B(n_6219),
.C(n_6098),
.Y(n_8907)
);

OR2x2_ASAP7_75t_L g8908 ( 
.A(n_8660),
.B(n_5581),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8728),
.Y(n_8909)
);

INVxp67_ASAP7_75t_SL g8910 ( 
.A(n_8671),
.Y(n_8910)
);

AOI21xp33_ASAP7_75t_L g8911 ( 
.A1(n_8717),
.A2(n_6219),
.B(n_6098),
.Y(n_8911)
);

OAI21xp5_ASAP7_75t_L g8912 ( 
.A1(n_8659),
.A2(n_5135),
.B(n_5149),
.Y(n_8912)
);

OAI21xp5_ASAP7_75t_SL g8913 ( 
.A1(n_8721),
.A2(n_5362),
.B(n_5461),
.Y(n_8913)
);

INVx2_ASAP7_75t_L g8914 ( 
.A(n_8692),
.Y(n_8914)
);

OAI22xp5_ASAP7_75t_L g8915 ( 
.A1(n_8581),
.A2(n_5672),
.B1(n_5710),
.B2(n_5622),
.Y(n_8915)
);

AO22x2_ASAP7_75t_L g8916 ( 
.A1(n_8729),
.A2(n_5643),
.B1(n_5654),
.B2(n_5644),
.Y(n_8916)
);

AOI222xp33_ASAP7_75t_L g8917 ( 
.A1(n_8729),
.A2(n_5657),
.B1(n_5658),
.B2(n_5669),
.C1(n_5666),
.C2(n_5641),
.Y(n_8917)
);

INVx2_ASAP7_75t_L g8918 ( 
.A(n_8684),
.Y(n_8918)
);

AND2x2_ASAP7_75t_L g8919 ( 
.A(n_8714),
.B(n_5594),
.Y(n_8919)
);

AOI22xp33_ASAP7_75t_SL g8920 ( 
.A1(n_8678),
.A2(n_5286),
.B1(n_6098),
.B2(n_5619),
.Y(n_8920)
);

INVx1_ASAP7_75t_SL g8921 ( 
.A(n_8682),
.Y(n_8921)
);

INVxp67_ASAP7_75t_SL g8922 ( 
.A(n_8686),
.Y(n_8922)
);

AOI22xp5_ASAP7_75t_L g8923 ( 
.A1(n_8768),
.A2(n_8739),
.B1(n_8627),
.B2(n_8677),
.Y(n_8923)
);

AOI222xp33_ASAP7_75t_L g8924 ( 
.A1(n_8828),
.A2(n_8739),
.B1(n_8748),
.B2(n_8651),
.C1(n_8644),
.C2(n_8626),
.Y(n_8924)
);

AOI22xp33_ASAP7_75t_L g8925 ( 
.A1(n_8806),
.A2(n_8717),
.B1(n_8750),
.B2(n_8653),
.Y(n_8925)
);

INVx2_ASAP7_75t_L g8926 ( 
.A(n_8838),
.Y(n_8926)
);

OAI21xp5_ASAP7_75t_L g8927 ( 
.A1(n_8754),
.A2(n_8640),
.B(n_8645),
.Y(n_8927)
);

NAND3xp33_ASAP7_75t_L g8928 ( 
.A(n_8795),
.B(n_8698),
.C(n_8690),
.Y(n_8928)
);

NAND2xp33_ASAP7_75t_L g8929 ( 
.A(n_8760),
.B(n_8655),
.Y(n_8929)
);

NOR2xp33_ASAP7_75t_L g8930 ( 
.A(n_8823),
.B(n_8661),
.Y(n_8930)
);

NAND2x1_ASAP7_75t_L g8931 ( 
.A(n_8774),
.B(n_8663),
.Y(n_8931)
);

AOI22xp5_ASAP7_75t_L g8932 ( 
.A1(n_8804),
.A2(n_8668),
.B1(n_8667),
.B2(n_8665),
.Y(n_8932)
);

AND2x2_ASAP7_75t_L g8933 ( 
.A(n_8774),
.B(n_8815),
.Y(n_8933)
);

AOI221x1_ASAP7_75t_L g8934 ( 
.A1(n_8832),
.A2(n_8687),
.B1(n_8669),
.B2(n_5590),
.C(n_5591),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8759),
.B(n_5583),
.Y(n_8935)
);

OAI22xp5_ASAP7_75t_L g8936 ( 
.A1(n_8883),
.A2(n_5587),
.B1(n_5591),
.B2(n_5583),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_8773),
.Y(n_8937)
);

INVx1_ASAP7_75t_L g8938 ( 
.A(n_8781),
.Y(n_8938)
);

AND2x2_ASAP7_75t_L g8939 ( 
.A(n_8850),
.B(n_5594),
.Y(n_8939)
);

INVx1_ASAP7_75t_L g8940 ( 
.A(n_8817),
.Y(n_8940)
);

OAI21xp33_ASAP7_75t_L g8941 ( 
.A1(n_8798),
.A2(n_5596),
.B(n_5587),
.Y(n_8941)
);

INVxp67_ASAP7_75t_SL g8942 ( 
.A(n_8788),
.Y(n_8942)
);

AOI21xp5_ASAP7_75t_L g8943 ( 
.A1(n_8762),
.A2(n_5605),
.B(n_5596),
.Y(n_8943)
);

A2O1A1Ixp33_ASAP7_75t_L g8944 ( 
.A1(n_8860),
.A2(n_8770),
.B(n_8753),
.C(n_8791),
.Y(n_8944)
);

INVx1_ASAP7_75t_L g8945 ( 
.A(n_8818),
.Y(n_8945)
);

NAND2xp5_ASAP7_75t_L g8946 ( 
.A(n_8787),
.B(n_5605),
.Y(n_8946)
);

AND2x2_ASAP7_75t_L g8947 ( 
.A(n_8894),
.B(n_5597),
.Y(n_8947)
);

A2O1A1Ixp33_ASAP7_75t_L g8948 ( 
.A1(n_8846),
.A2(n_5669),
.B(n_5670),
.C(n_5666),
.Y(n_8948)
);

INVx1_ASAP7_75t_L g8949 ( 
.A(n_8783),
.Y(n_8949)
);

NAND2xp5_ASAP7_75t_L g8950 ( 
.A(n_8789),
.B(n_5608),
.Y(n_8950)
);

INVx2_ASAP7_75t_SL g8951 ( 
.A(n_8799),
.Y(n_8951)
);

INVx1_ASAP7_75t_L g8952 ( 
.A(n_8769),
.Y(n_8952)
);

AND2x2_ASAP7_75t_SL g8953 ( 
.A(n_8756),
.B(n_5597),
.Y(n_8953)
);

AOI21xp5_ASAP7_75t_SL g8954 ( 
.A1(n_8777),
.A2(n_5619),
.B(n_5597),
.Y(n_8954)
);

AND2x2_ASAP7_75t_L g8955 ( 
.A(n_8919),
.B(n_5597),
.Y(n_8955)
);

INVx1_ASAP7_75t_L g8956 ( 
.A(n_8910),
.Y(n_8956)
);

OAI22xp5_ASAP7_75t_SL g8957 ( 
.A1(n_8866),
.A2(n_5034),
.B1(n_5046),
.B2(n_5000),
.Y(n_8957)
);

NOR2xp33_ASAP7_75t_L g8958 ( 
.A(n_8779),
.B(n_6153),
.Y(n_8958)
);

AOI21xp33_ASAP7_75t_SL g8959 ( 
.A1(n_8761),
.A2(n_5193),
.B(n_6116),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_8922),
.Y(n_8960)
);

INVxp67_ASAP7_75t_SL g8961 ( 
.A(n_8752),
.Y(n_8961)
);

AND2x2_ASAP7_75t_L g8962 ( 
.A(n_8853),
.B(n_5619),
.Y(n_8962)
);

OR2x2_ASAP7_75t_L g8963 ( 
.A(n_8852),
.B(n_5608),
.Y(n_8963)
);

OAI221xp5_ASAP7_75t_L g8964 ( 
.A1(n_8763),
.A2(n_6116),
.B1(n_6125),
.B2(n_6149),
.C(n_4876),
.Y(n_8964)
);

AOI22xp33_ASAP7_75t_L g8965 ( 
.A1(n_8819),
.A2(n_5935),
.B1(n_6149),
.B2(n_6125),
.Y(n_8965)
);

AND2x2_ASAP7_75t_L g8966 ( 
.A(n_8859),
.B(n_8878),
.Y(n_8966)
);

AOI21xp33_ASAP7_75t_L g8967 ( 
.A1(n_8771),
.A2(n_6149),
.B(n_6116),
.Y(n_8967)
);

AOI221xp5_ASAP7_75t_L g8968 ( 
.A1(n_8757),
.A2(n_6153),
.B1(n_6202),
.B2(n_6203),
.C(n_6157),
.Y(n_8968)
);

NOR2xp33_ASAP7_75t_L g8969 ( 
.A(n_8841),
.B(n_6125),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_8870),
.Y(n_8970)
);

NOR2xp33_ASAP7_75t_L g8971 ( 
.A(n_8786),
.B(n_5266),
.Y(n_8971)
);

INVx1_ASAP7_75t_L g8972 ( 
.A(n_8810),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8811),
.Y(n_8973)
);

INVx1_ASAP7_75t_L g8974 ( 
.A(n_8813),
.Y(n_8974)
);

AND2x2_ASAP7_75t_L g8975 ( 
.A(n_8888),
.B(n_5619),
.Y(n_8975)
);

AOI21xp33_ASAP7_75t_SL g8976 ( 
.A1(n_8885),
.A2(n_5193),
.B(n_5725),
.Y(n_8976)
);

AOI21xp5_ASAP7_75t_L g8977 ( 
.A1(n_8758),
.A2(n_8780),
.B(n_8755),
.Y(n_8977)
);

NAND2xp5_ASAP7_75t_L g8978 ( 
.A(n_8873),
.B(n_5617),
.Y(n_8978)
);

AOI21xp33_ASAP7_75t_L g8979 ( 
.A1(n_8767),
.A2(n_6202),
.B(n_6157),
.Y(n_8979)
);

AOI222xp33_ASAP7_75t_L g8980 ( 
.A1(n_8881),
.A2(n_5682),
.B1(n_5671),
.B2(n_5688),
.C1(n_5680),
.C2(n_5670),
.Y(n_8980)
);

AOI222xp33_ASAP7_75t_L g8981 ( 
.A1(n_8907),
.A2(n_5688),
.B1(n_5680),
.B2(n_5690),
.C1(n_5682),
.C2(n_5671),
.Y(n_8981)
);

NAND2xp5_ASAP7_75t_SL g8982 ( 
.A(n_8763),
.B(n_5650),
.Y(n_8982)
);

NOR2xp33_ASAP7_75t_L g8983 ( 
.A(n_8874),
.B(n_5266),
.Y(n_8983)
);

NAND2xp5_ASAP7_75t_SL g8984 ( 
.A(n_8793),
.B(n_5650),
.Y(n_8984)
);

NAND2xp5_ASAP7_75t_L g8985 ( 
.A(n_8778),
.B(n_5617),
.Y(n_8985)
);

OAI221xp5_ASAP7_75t_L g8986 ( 
.A1(n_8902),
.A2(n_5193),
.B1(n_4409),
.B2(n_5691),
.C(n_5690),
.Y(n_8986)
);

NAND2xp5_ASAP7_75t_L g8987 ( 
.A(n_8921),
.B(n_8793),
.Y(n_8987)
);

AOI21xp5_ASAP7_75t_SL g8988 ( 
.A1(n_8785),
.A2(n_5650),
.B(n_5182),
.Y(n_8988)
);

AOI21xp33_ASAP7_75t_L g8989 ( 
.A1(n_8772),
.A2(n_6202),
.B(n_6157),
.Y(n_8989)
);

OAI221xp5_ASAP7_75t_L g8990 ( 
.A1(n_8796),
.A2(n_8797),
.B1(n_8920),
.B2(n_8805),
.C(n_8776),
.Y(n_8990)
);

OAI21xp5_ASAP7_75t_L g8991 ( 
.A1(n_8898),
.A2(n_5622),
.B(n_5621),
.Y(n_8991)
);

OAI22xp5_ASAP7_75t_L g8992 ( 
.A1(n_8827),
.A2(n_8807),
.B1(n_8897),
.B2(n_8803),
.Y(n_8992)
);

AND2x2_ASAP7_75t_L g8993 ( 
.A(n_8792),
.B(n_5650),
.Y(n_8993)
);

INVxp67_ASAP7_75t_L g8994 ( 
.A(n_8764),
.Y(n_8994)
);

AOI221xp5_ASAP7_75t_L g8995 ( 
.A1(n_8775),
.A2(n_6203),
.B1(n_5711),
.B2(n_5713),
.C(n_5706),
.Y(n_8995)
);

NOR2xp33_ASAP7_75t_L g8996 ( 
.A(n_8865),
.B(n_5266),
.Y(n_8996)
);

AOI322xp5_ASAP7_75t_L g8997 ( 
.A1(n_8884),
.A2(n_5735),
.A3(n_5716),
.B1(n_5713),
.B2(n_5714),
.C1(n_5706),
.C2(n_5711),
.Y(n_8997)
);

OAI21xp33_ASAP7_75t_L g8998 ( 
.A1(n_8794),
.A2(n_5626),
.B(n_5621),
.Y(n_8998)
);

NOR2xp33_ASAP7_75t_L g8999 ( 
.A(n_8782),
.B(n_5313),
.Y(n_8999)
);

INVx2_ASAP7_75t_L g9000 ( 
.A(n_8901),
.Y(n_9000)
);

INVxp67_ASAP7_75t_L g9001 ( 
.A(n_8821),
.Y(n_9001)
);

AOI222xp33_ASAP7_75t_L g9002 ( 
.A1(n_8863),
.A2(n_5722),
.B1(n_5714),
.B2(n_5735),
.C1(n_5716),
.C2(n_5691),
.Y(n_9002)
);

OAI21xp33_ASAP7_75t_L g9003 ( 
.A1(n_8826),
.A2(n_5627),
.B(n_5626),
.Y(n_9003)
);

AND2x2_ASAP7_75t_L g9004 ( 
.A(n_8843),
.B(n_5628),
.Y(n_9004)
);

NAND2xp5_ASAP7_75t_SL g9005 ( 
.A(n_8914),
.B(n_5286),
.Y(n_9005)
);

OAI31xp33_ASAP7_75t_L g9006 ( 
.A1(n_8830),
.A2(n_5286),
.A3(n_5722),
.B(n_4726),
.Y(n_9006)
);

OAI21xp5_ASAP7_75t_L g9007 ( 
.A1(n_8801),
.A2(n_5629),
.B(n_5628),
.Y(n_9007)
);

OR2x2_ASAP7_75t_L g9008 ( 
.A(n_8766),
.B(n_5629),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_8887),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8905),
.Y(n_9010)
);

O2A1O1Ixp33_ASAP7_75t_L g9011 ( 
.A1(n_8876),
.A2(n_6203),
.B(n_5193),
.C(n_5371),
.Y(n_9011)
);

OR2x2_ASAP7_75t_L g9012 ( 
.A(n_8918),
.B(n_8877),
.Y(n_9012)
);

INVx1_ASAP7_75t_L g9013 ( 
.A(n_8879),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8893),
.Y(n_9014)
);

INVx1_ASAP7_75t_L g9015 ( 
.A(n_8893),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_8837),
.Y(n_9016)
);

AOI22xp5_ASAP7_75t_L g9017 ( 
.A1(n_8808),
.A2(n_5286),
.B1(n_5386),
.B2(n_5313),
.Y(n_9017)
);

NAND2xp5_ASAP7_75t_L g9018 ( 
.A(n_8909),
.B(n_5631),
.Y(n_9018)
);

AOI21xp33_ASAP7_75t_SL g9019 ( 
.A1(n_8855),
.A2(n_5371),
.B(n_4680),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8842),
.Y(n_9020)
);

OAI21xp33_ASAP7_75t_SL g9021 ( 
.A1(n_8875),
.A2(n_5635),
.B(n_5631),
.Y(n_9021)
);

AOI21xp33_ASAP7_75t_L g9022 ( 
.A1(n_8847),
.A2(n_5386),
.B(n_5313),
.Y(n_9022)
);

AND2x2_ASAP7_75t_L g9023 ( 
.A(n_8765),
.B(n_5640),
.Y(n_9023)
);

AOI22xp5_ASAP7_75t_L g9024 ( 
.A1(n_8854),
.A2(n_5386),
.B1(n_5515),
.B2(n_5511),
.Y(n_9024)
);

OAI32xp33_ASAP7_75t_L g9025 ( 
.A1(n_8790),
.A2(n_5655),
.A3(n_5661),
.B1(n_5653),
.B2(n_5640),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_L g9026 ( 
.A(n_8862),
.B(n_5653),
.Y(n_9026)
);

OAI21xp5_ASAP7_75t_SL g9027 ( 
.A1(n_8802),
.A2(n_5182),
.B(n_5171),
.Y(n_9027)
);

OAI21xp33_ASAP7_75t_SL g9028 ( 
.A1(n_8833),
.A2(n_5661),
.B(n_5655),
.Y(n_9028)
);

OAI21xp33_ASAP7_75t_L g9029 ( 
.A1(n_8836),
.A2(n_5665),
.B(n_5664),
.Y(n_9029)
);

AOI222xp33_ASAP7_75t_L g9030 ( 
.A1(n_8899),
.A2(n_5515),
.B1(n_5518),
.B2(n_5531),
.C1(n_5522),
.C2(n_5511),
.Y(n_9030)
);

AND2x2_ASAP7_75t_L g9031 ( 
.A(n_8814),
.B(n_5665),
.Y(n_9031)
);

OAI31xp33_ASAP7_75t_L g9032 ( 
.A1(n_8869),
.A2(n_4822),
.A3(n_4812),
.B(n_4763),
.Y(n_9032)
);

AOI21xp33_ASAP7_75t_L g9033 ( 
.A1(n_8784),
.A2(n_5522),
.B(n_5518),
.Y(n_9033)
);

NAND2xp5_ASAP7_75t_L g9034 ( 
.A(n_8904),
.B(n_5672),
.Y(n_9034)
);

BUFx2_ASAP7_75t_L g9035 ( 
.A(n_8834),
.Y(n_9035)
);

NOR2xp33_ASAP7_75t_L g9036 ( 
.A(n_8809),
.B(n_5674),
.Y(n_9036)
);

INVx2_ASAP7_75t_SL g9037 ( 
.A(n_8896),
.Y(n_9037)
);

NOR2xp33_ASAP7_75t_L g9038 ( 
.A(n_8824),
.B(n_5674),
.Y(n_9038)
);

OAI21xp5_ASAP7_75t_SL g9039 ( 
.A1(n_8839),
.A2(n_5182),
.B(n_5171),
.Y(n_9039)
);

NAND2xp5_ASAP7_75t_L g9040 ( 
.A(n_8816),
.B(n_5678),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_8825),
.Y(n_9041)
);

NAND3x2_ASAP7_75t_L g9042 ( 
.A(n_8840),
.B(n_5681),
.C(n_5678),
.Y(n_9042)
);

INVx1_ASAP7_75t_L g9043 ( 
.A(n_8851),
.Y(n_9043)
);

NOR3xp33_ASAP7_75t_L g9044 ( 
.A(n_8911),
.B(n_4631),
.C(n_4671),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_8908),
.Y(n_9045)
);

OAI33xp33_ASAP7_75t_L g9046 ( 
.A1(n_8889),
.A2(n_5684),
.A3(n_5685),
.B1(n_5694),
.B2(n_5692),
.B3(n_5681),
.Y(n_9046)
);

INVx1_ASAP7_75t_SL g9047 ( 
.A(n_8800),
.Y(n_9047)
);

AOI22xp33_ASAP7_75t_SL g9048 ( 
.A1(n_8882),
.A2(n_5171),
.B1(n_5182),
.B2(n_5371),
.Y(n_9048)
);

OR2x2_ASAP7_75t_L g9049 ( 
.A(n_8864),
.B(n_5684),
.Y(n_9049)
);

AOI21xp33_ASAP7_75t_L g9050 ( 
.A1(n_8891),
.A2(n_8849),
.B(n_8829),
.Y(n_9050)
);

AO32x1_ASAP7_75t_L g9051 ( 
.A1(n_8915),
.A2(n_5685),
.A3(n_5695),
.B1(n_5694),
.B2(n_5692),
.Y(n_9051)
);

AOI22xp33_ASAP7_75t_L g9052 ( 
.A1(n_8906),
.A2(n_5531),
.B1(n_5536),
.B2(n_5535),
.Y(n_9052)
);

AOI22xp33_ASAP7_75t_L g9053 ( 
.A1(n_8900),
.A2(n_5535),
.B1(n_5538),
.B2(n_5536),
.Y(n_9053)
);

INVx1_ASAP7_75t_SL g9054 ( 
.A(n_8880),
.Y(n_9054)
);

OAI221xp5_ASAP7_75t_L g9055 ( 
.A1(n_8871),
.A2(n_4409),
.B1(n_5696),
.B2(n_5544),
.C(n_4445),
.Y(n_9055)
);

AOI221xp5_ASAP7_75t_SL g9056 ( 
.A1(n_8820),
.A2(n_5695),
.B1(n_5719),
.B2(n_5712),
.C(n_5710),
.Y(n_9056)
);

NOR2xp67_ASAP7_75t_L g9057 ( 
.A(n_8857),
.B(n_5712),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_8886),
.Y(n_9058)
);

NAND2xp5_ASAP7_75t_L g9059 ( 
.A(n_8895),
.B(n_5719),
.Y(n_9059)
);

NAND2xp5_ASAP7_75t_SL g9060 ( 
.A(n_8848),
.B(n_5171),
.Y(n_9060)
);

O2A1O1Ixp5_ASAP7_75t_L g9061 ( 
.A1(n_8845),
.A2(n_5724),
.B(n_5729),
.C(n_5720),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8861),
.Y(n_9062)
);

AOI22xp5_ASAP7_75t_L g9063 ( 
.A1(n_8831),
.A2(n_5571),
.B1(n_5578),
.B2(n_5564),
.Y(n_9063)
);

AOI221xp5_ASAP7_75t_L g9064 ( 
.A1(n_8912),
.A2(n_5585),
.B1(n_5578),
.B2(n_5571),
.C(n_5550),
.Y(n_9064)
);

OAI21xp33_ASAP7_75t_L g9065 ( 
.A1(n_8856),
.A2(n_5729),
.B(n_5724),
.Y(n_9065)
);

NAND2xp5_ASAP7_75t_L g9066 ( 
.A(n_8903),
.B(n_8867),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8933),
.Y(n_9067)
);

INVx1_ASAP7_75t_L g9068 ( 
.A(n_8942),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_8931),
.Y(n_9069)
);

NAND2xp5_ASAP7_75t_L g9070 ( 
.A(n_8926),
.B(n_8868),
.Y(n_9070)
);

NAND2x1p5_ASAP7_75t_L g9071 ( 
.A(n_8949),
.B(n_8812),
.Y(n_9071)
);

AND2x2_ASAP7_75t_L g9072 ( 
.A(n_8953),
.B(n_8913),
.Y(n_9072)
);

NAND2xp5_ASAP7_75t_L g9073 ( 
.A(n_8961),
.B(n_8822),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_9012),
.Y(n_9074)
);

NOR2xp33_ASAP7_75t_L g9075 ( 
.A(n_8956),
.B(n_8844),
.Y(n_9075)
);

AND2x2_ASAP7_75t_L g9076 ( 
.A(n_8966),
.B(n_8939),
.Y(n_9076)
);

NOR2xp67_ASAP7_75t_SL g9077 ( 
.A(n_8960),
.B(n_8858),
.Y(n_9077)
);

CKINVDCx16_ASAP7_75t_R g9078 ( 
.A(n_8951),
.Y(n_9078)
);

NAND2xp5_ASAP7_75t_L g9079 ( 
.A(n_9047),
.B(n_8890),
.Y(n_9079)
);

NAND2xp5_ASAP7_75t_L g9080 ( 
.A(n_9035),
.B(n_8835),
.Y(n_9080)
);

INVx2_ASAP7_75t_L g9081 ( 
.A(n_8955),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8929),
.Y(n_9082)
);

NAND2x1_ASAP7_75t_SL g9083 ( 
.A(n_8937),
.B(n_8892),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_9000),
.Y(n_9084)
);

INVx2_ASAP7_75t_L g9085 ( 
.A(n_8962),
.Y(n_9085)
);

AND2x2_ASAP7_75t_L g9086 ( 
.A(n_8947),
.B(n_8916),
.Y(n_9086)
);

NAND2xp5_ASAP7_75t_L g9087 ( 
.A(n_9037),
.B(n_8872),
.Y(n_9087)
);

AND2x2_ASAP7_75t_L g9088 ( 
.A(n_8975),
.B(n_8916),
.Y(n_9088)
);

INVx1_ASAP7_75t_L g9089 ( 
.A(n_8987),
.Y(n_9089)
);

INVx2_ASAP7_75t_L g9090 ( 
.A(n_8993),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_9014),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_L g9092 ( 
.A(n_8930),
.B(n_8917),
.Y(n_9092)
);

NAND2xp5_ASAP7_75t_L g9093 ( 
.A(n_8977),
.B(n_5732),
.Y(n_9093)
);

NOR2x1_ASAP7_75t_L g9094 ( 
.A(n_8928),
.B(n_5732),
.Y(n_9094)
);

INVxp67_ASAP7_75t_L g9095 ( 
.A(n_8958),
.Y(n_9095)
);

AND2x2_ASAP7_75t_L g9096 ( 
.A(n_8938),
.B(n_5733),
.Y(n_9096)
);

AND2x2_ASAP7_75t_L g9097 ( 
.A(n_9054),
.B(n_5733),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_9015),
.Y(n_9098)
);

OR2x2_ASAP7_75t_L g9099 ( 
.A(n_8992),
.B(n_5371),
.Y(n_9099)
);

INVx1_ASAP7_75t_SL g9100 ( 
.A(n_8940),
.Y(n_9100)
);

NAND2xp5_ASAP7_75t_L g9101 ( 
.A(n_9045),
.B(n_4578),
.Y(n_9101)
);

NOR2xp67_ASAP7_75t_L g9102 ( 
.A(n_9001),
.B(n_8923),
.Y(n_9102)
);

OAI22xp5_ASAP7_75t_L g9103 ( 
.A1(n_8923),
.A2(n_5034),
.B1(n_5046),
.B2(n_5000),
.Y(n_9103)
);

NAND2xp5_ASAP7_75t_L g9104 ( 
.A(n_9043),
.B(n_4578),
.Y(n_9104)
);

NAND2xp5_ASAP7_75t_L g9105 ( 
.A(n_8925),
.B(n_4578),
.Y(n_9105)
);

OR2x2_ASAP7_75t_L g9106 ( 
.A(n_8945),
.B(n_8972),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_9009),
.Y(n_9107)
);

NAND2xp5_ASAP7_75t_SL g9108 ( 
.A(n_9010),
.B(n_4607),
.Y(n_9108)
);

NAND2xp5_ASAP7_75t_L g9109 ( 
.A(n_9013),
.B(n_4578),
.Y(n_9109)
);

AND2x2_ASAP7_75t_L g9110 ( 
.A(n_8952),
.B(n_5000),
.Y(n_9110)
);

INVx1_ASAP7_75t_L g9111 ( 
.A(n_8973),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8974),
.Y(n_9112)
);

AND2x2_ASAP7_75t_L g9113 ( 
.A(n_8954),
.B(n_5000),
.Y(n_9113)
);

OR2x2_ASAP7_75t_L g9114 ( 
.A(n_9016),
.B(n_3994),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_9020),
.Y(n_9115)
);

OR2x2_ASAP7_75t_L g9116 ( 
.A(n_9041),
.B(n_8985),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_L g9117 ( 
.A(n_8994),
.B(n_9023),
.Y(n_9117)
);

AND2x2_ASAP7_75t_L g9118 ( 
.A(n_8988),
.B(n_5034),
.Y(n_9118)
);

AND2x2_ASAP7_75t_L g9119 ( 
.A(n_8927),
.B(n_5034),
.Y(n_9119)
);

NAND2xp5_ASAP7_75t_L g9120 ( 
.A(n_9004),
.B(n_5538),
.Y(n_9120)
);

NAND2xp5_ASAP7_75t_L g9121 ( 
.A(n_8932),
.B(n_5548),
.Y(n_9121)
);

NAND2xp5_ASAP7_75t_L g9122 ( 
.A(n_9058),
.B(n_5548),
.Y(n_9122)
);

INVx1_ASAP7_75t_L g9123 ( 
.A(n_9031),
.Y(n_9123)
);

NAND2xp5_ASAP7_75t_L g9124 ( 
.A(n_8969),
.B(n_5550),
.Y(n_9124)
);

INVx1_ASAP7_75t_L g9125 ( 
.A(n_8963),
.Y(n_9125)
);

AND2x2_ASAP7_75t_L g9126 ( 
.A(n_8984),
.B(n_5046),
.Y(n_9126)
);

INVx2_ASAP7_75t_SL g9127 ( 
.A(n_8982),
.Y(n_9127)
);

AND2x2_ASAP7_75t_L g9128 ( 
.A(n_9005),
.B(n_5046),
.Y(n_9128)
);

INVx1_ASAP7_75t_SL g9129 ( 
.A(n_9066),
.Y(n_9129)
);

INVx1_ASAP7_75t_L g9130 ( 
.A(n_9051),
.Y(n_9130)
);

NAND2xp5_ASAP7_75t_SL g9131 ( 
.A(n_8944),
.B(n_8924),
.Y(n_9131)
);

OAI221xp5_ASAP7_75t_L g9132 ( 
.A1(n_8990),
.A2(n_5544),
.B1(n_5696),
.B2(n_5564),
.C(n_5560),
.Y(n_9132)
);

NAND2xp5_ASAP7_75t_L g9133 ( 
.A(n_8934),
.B(n_5553),
.Y(n_9133)
);

NAND2xp5_ASAP7_75t_L g9134 ( 
.A(n_9036),
.B(n_5553),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_9049),
.Y(n_9135)
);

NAND2xp5_ASAP7_75t_L g9136 ( 
.A(n_9038),
.B(n_5560),
.Y(n_9136)
);

NOR2xp33_ASAP7_75t_L g9137 ( 
.A(n_8976),
.B(n_5585),
.Y(n_9137)
);

INVx2_ASAP7_75t_L g9138 ( 
.A(n_9061),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_9051),
.Y(n_9139)
);

AND2x2_ASAP7_75t_L g9140 ( 
.A(n_9062),
.B(n_9039),
.Y(n_9140)
);

INVx1_ASAP7_75t_SL g9141 ( 
.A(n_9008),
.Y(n_9141)
);

AND2x2_ASAP7_75t_L g9142 ( 
.A(n_9027),
.B(n_5067),
.Y(n_9142)
);

INVx1_ASAP7_75t_L g9143 ( 
.A(n_8978),
.Y(n_9143)
);

INVxp67_ASAP7_75t_L g9144 ( 
.A(n_8970),
.Y(n_9144)
);

INVx1_ASAP7_75t_L g9145 ( 
.A(n_9051),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_9059),
.Y(n_9146)
);

NOR2xp33_ASAP7_75t_L g9147 ( 
.A(n_9060),
.B(n_5267),
.Y(n_9147)
);

INVx1_ASAP7_75t_L g9148 ( 
.A(n_9040),
.Y(n_9148)
);

INVx2_ASAP7_75t_L g9149 ( 
.A(n_8935),
.Y(n_9149)
);

OAI22xp5_ASAP7_75t_L g9150 ( 
.A1(n_8964),
.A2(n_5067),
.B1(n_4589),
.B2(n_4909),
.Y(n_9150)
);

NAND2xp5_ASAP7_75t_L g9151 ( 
.A(n_9057),
.B(n_5149),
.Y(n_9151)
);

OR2x2_ASAP7_75t_L g9152 ( 
.A(n_9026),
.B(n_3994),
.Y(n_9152)
);

NAND2xp5_ASAP7_75t_L g9153 ( 
.A(n_8983),
.B(n_4861),
.Y(n_9153)
);

INVx1_ASAP7_75t_L g9154 ( 
.A(n_9018),
.Y(n_9154)
);

INVx1_ASAP7_75t_L g9155 ( 
.A(n_8946),
.Y(n_9155)
);

INVx2_ASAP7_75t_SL g9156 ( 
.A(n_8950),
.Y(n_9156)
);

NAND2x1_ASAP7_75t_L g9157 ( 
.A(n_8991),
.B(n_5089),
.Y(n_9157)
);

BUFx4f_ASAP7_75t_SL g9158 ( 
.A(n_9042),
.Y(n_9158)
);

NAND2x1_ASAP7_75t_SL g9159 ( 
.A(n_8971),
.B(n_8999),
.Y(n_9159)
);

AND2x4_ASAP7_75t_L g9160 ( 
.A(n_9007),
.B(n_4607),
.Y(n_9160)
);

NAND2xp5_ASAP7_75t_L g9161 ( 
.A(n_9056),
.B(n_4861),
.Y(n_9161)
);

NAND2xp5_ASAP7_75t_L g9162 ( 
.A(n_8943),
.B(n_4861),
.Y(n_9162)
);

INVx1_ASAP7_75t_L g9163 ( 
.A(n_9034),
.Y(n_9163)
);

NAND2xp5_ASAP7_75t_L g9164 ( 
.A(n_8996),
.B(n_4861),
.Y(n_9164)
);

NAND2xp5_ASAP7_75t_L g9165 ( 
.A(n_8995),
.B(n_4885),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_9028),
.Y(n_9166)
);

AND2x2_ASAP7_75t_L g9167 ( 
.A(n_9048),
.B(n_5067),
.Y(n_9167)
);

INVxp67_ASAP7_75t_L g9168 ( 
.A(n_9050),
.Y(n_9168)
);

NAND2x1_ASAP7_75t_SL g9169 ( 
.A(n_9024),
.B(n_4401),
.Y(n_9169)
);

NOR2xp33_ASAP7_75t_L g9170 ( 
.A(n_9021),
.B(n_5267),
.Y(n_9170)
);

AO22x2_ASAP7_75t_L g9171 ( 
.A1(n_8979),
.A2(n_4160),
.B1(n_4331),
.B2(n_4427),
.Y(n_9171)
);

OR2x2_ASAP7_75t_L g9172 ( 
.A(n_9065),
.B(n_3994),
.Y(n_9172)
);

INVx1_ASAP7_75t_SL g9173 ( 
.A(n_8957),
.Y(n_9173)
);

HB1xp67_ASAP7_75t_L g9174 ( 
.A(n_8967),
.Y(n_9174)
);

AND2x2_ASAP7_75t_L g9175 ( 
.A(n_8959),
.B(n_5067),
.Y(n_9175)
);

AND2x2_ASAP7_75t_L g9176 ( 
.A(n_8941),
.B(n_4607),
.Y(n_9176)
);

NOR3xp33_ASAP7_75t_L g9177 ( 
.A(n_8989),
.B(n_4575),
.C(n_4572),
.Y(n_9177)
);

HB1xp67_ASAP7_75t_L g9178 ( 
.A(n_8968),
.Y(n_9178)
);

HB1xp67_ASAP7_75t_L g9179 ( 
.A(n_9022),
.Y(n_9179)
);

INVx1_ASAP7_75t_L g9180 ( 
.A(n_9003),
.Y(n_9180)
);

CKINVDCx16_ASAP7_75t_R g9181 ( 
.A(n_8936),
.Y(n_9181)
);

INVx1_ASAP7_75t_L g9182 ( 
.A(n_8998),
.Y(n_9182)
);

NAND2xp5_ASAP7_75t_L g9183 ( 
.A(n_9029),
.B(n_4885),
.Y(n_9183)
);

NOR2xp33_ASAP7_75t_L g9184 ( 
.A(n_9046),
.B(n_5272),
.Y(n_9184)
);

NOR2xp33_ASAP7_75t_L g9185 ( 
.A(n_9168),
.B(n_8986),
.Y(n_9185)
);

NOR3x1_ASAP7_75t_L g9186 ( 
.A(n_9127),
.B(n_9055),
.C(n_9032),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_L g9187 ( 
.A(n_9078),
.B(n_9076),
.Y(n_9187)
);

AOI21xp33_ASAP7_75t_L g9188 ( 
.A1(n_9100),
.A2(n_8965),
.B(n_9002),
.Y(n_9188)
);

OAI21xp5_ASAP7_75t_SL g9189 ( 
.A1(n_9067),
.A2(n_9019),
.B(n_9006),
.Y(n_9189)
);

INVx1_ASAP7_75t_L g9190 ( 
.A(n_9067),
.Y(n_9190)
);

INVxp67_ASAP7_75t_L g9191 ( 
.A(n_9069),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_9074),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_SL g9193 ( 
.A(n_9069),
.B(n_9017),
.Y(n_9193)
);

NAND2xp5_ASAP7_75t_L g9194 ( 
.A(n_9129),
.B(n_9030),
.Y(n_9194)
);

NAND3xp33_ASAP7_75t_L g9195 ( 
.A(n_9131),
.B(n_9033),
.C(n_9052),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_9088),
.B(n_9086),
.Y(n_9196)
);

NOR2xp33_ASAP7_75t_SL g9197 ( 
.A(n_9084),
.B(n_9011),
.Y(n_9197)
);

CKINVDCx14_ASAP7_75t_R g9198 ( 
.A(n_9082),
.Y(n_9198)
);

AOI211xp5_ASAP7_75t_SL g9199 ( 
.A1(n_9102),
.A2(n_9044),
.B(n_8948),
.C(n_9025),
.Y(n_9199)
);

INVx2_ASAP7_75t_L g9200 ( 
.A(n_9071),
.Y(n_9200)
);

INVx1_ASAP7_75t_L g9201 ( 
.A(n_9106),
.Y(n_9201)
);

AOI21xp5_ASAP7_75t_L g9202 ( 
.A1(n_9068),
.A2(n_9053),
.B(n_9063),
.Y(n_9202)
);

NAND2xp5_ASAP7_75t_L g9203 ( 
.A(n_9068),
.B(n_8997),
.Y(n_9203)
);

INVx2_ASAP7_75t_L g9204 ( 
.A(n_9116),
.Y(n_9204)
);

NOR3x1_ASAP7_75t_L g9205 ( 
.A(n_9079),
.B(n_4917),
.C(n_4887),
.Y(n_9205)
);

O2A1O1Ixp33_ASAP7_75t_SL g9206 ( 
.A1(n_9093),
.A2(n_9064),
.B(n_3801),
.C(n_5102),
.Y(n_9206)
);

NOR3xp33_ASAP7_75t_L g9207 ( 
.A(n_9144),
.B(n_8981),
.C(n_8980),
.Y(n_9207)
);

NAND3xp33_ASAP7_75t_SL g9208 ( 
.A(n_9141),
.B(n_4414),
.C(n_4645),
.Y(n_9208)
);

INVx1_ASAP7_75t_L g9209 ( 
.A(n_9081),
.Y(n_9209)
);

INVx1_ASAP7_75t_L g9210 ( 
.A(n_9085),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_9117),
.Y(n_9211)
);

INVx2_ASAP7_75t_L g9212 ( 
.A(n_9118),
.Y(n_9212)
);

AOI211xp5_ASAP7_75t_L g9213 ( 
.A1(n_9075),
.A2(n_4759),
.B(n_4902),
.C(n_4955),
.Y(n_9213)
);

NOR2xp67_ASAP7_75t_L g9214 ( 
.A(n_9089),
.B(n_4426),
.Y(n_9214)
);

OAI21xp33_ASAP7_75t_L g9215 ( 
.A1(n_9110),
.A2(n_4085),
.B(n_3977),
.Y(n_9215)
);

AOI211x1_ASAP7_75t_L g9216 ( 
.A1(n_9077),
.A2(n_9108),
.B(n_9132),
.C(n_9113),
.Y(n_9216)
);

NOR4xp25_ASAP7_75t_L g9217 ( 
.A(n_9095),
.B(n_4259),
.C(n_4852),
.D(n_4846),
.Y(n_9217)
);

NOR3x1_ASAP7_75t_L g9218 ( 
.A(n_9156),
.B(n_9112),
.C(n_9111),
.Y(n_9218)
);

OAI22xp5_ASAP7_75t_SL g9219 ( 
.A1(n_9181),
.A2(n_5696),
.B1(n_5544),
.B2(n_4792),
.Y(n_9219)
);

NOR3xp33_ASAP7_75t_L g9220 ( 
.A(n_9070),
.B(n_5168),
.C(n_5157),
.Y(n_9220)
);

NAND2xp5_ASAP7_75t_SL g9221 ( 
.A(n_9090),
.B(n_4911),
.Y(n_9221)
);

NAND3xp33_ASAP7_75t_L g9222 ( 
.A(n_9174),
.B(n_5071),
.C(n_5544),
.Y(n_9222)
);

AOI21xp5_ASAP7_75t_L g9223 ( 
.A1(n_9073),
.A2(n_4864),
.B(n_4860),
.Y(n_9223)
);

XNOR2xp5_ASAP7_75t_L g9224 ( 
.A(n_9072),
.B(n_5544),
.Y(n_9224)
);

OAI21xp33_ASAP7_75t_L g9225 ( 
.A1(n_9119),
.A2(n_4085),
.B(n_3977),
.Y(n_9225)
);

INVx2_ASAP7_75t_L g9226 ( 
.A(n_9135),
.Y(n_9226)
);

NOR2xp67_ASAP7_75t_L g9227 ( 
.A(n_9115),
.B(n_4426),
.Y(n_9227)
);

NAND2xp5_ASAP7_75t_SL g9228 ( 
.A(n_9107),
.B(n_4638),
.Y(n_9228)
);

INVx1_ASAP7_75t_L g9229 ( 
.A(n_9133),
.Y(n_9229)
);

NAND2xp5_ASAP7_75t_L g9230 ( 
.A(n_9146),
.B(n_5272),
.Y(n_9230)
);

INVx1_ASAP7_75t_L g9231 ( 
.A(n_9130),
.Y(n_9231)
);

OAI31xp33_ASAP7_75t_SL g9232 ( 
.A1(n_9094),
.A2(n_4971),
.A3(n_5022),
.B(n_4395),
.Y(n_9232)
);

AOI21xp5_ASAP7_75t_L g9233 ( 
.A1(n_9080),
.A2(n_4864),
.B(n_4860),
.Y(n_9233)
);

O2A1O1Ixp5_ASAP7_75t_L g9234 ( 
.A1(n_9138),
.A2(n_4438),
.B(n_4426),
.C(n_4638),
.Y(n_9234)
);

NAND2xp5_ASAP7_75t_L g9235 ( 
.A(n_9149),
.B(n_5157),
.Y(n_9235)
);

INVxp67_ASAP7_75t_SL g9236 ( 
.A(n_9083),
.Y(n_9236)
);

NOR3x1_ASAP7_75t_L g9237 ( 
.A(n_9148),
.B(n_4152),
.C(n_4115),
.Y(n_9237)
);

NAND3xp33_ASAP7_75t_L g9238 ( 
.A(n_9091),
.B(n_5696),
.C(n_5072),
.Y(n_9238)
);

NAND2xp5_ASAP7_75t_L g9239 ( 
.A(n_9125),
.B(n_5168),
.Y(n_9239)
);

INVxp67_ASAP7_75t_L g9240 ( 
.A(n_9092),
.Y(n_9240)
);

AOI21xp5_ASAP7_75t_SL g9241 ( 
.A1(n_9166),
.A2(n_5696),
.B(n_4303),
.Y(n_9241)
);

INVxp67_ASAP7_75t_L g9242 ( 
.A(n_9140),
.Y(n_9242)
);

NAND2xp33_ASAP7_75t_SL g9243 ( 
.A(n_9098),
.B(n_4401),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_9139),
.Y(n_9244)
);

NAND2xp5_ASAP7_75t_L g9245 ( 
.A(n_9143),
.B(n_9097),
.Y(n_9245)
);

NAND3xp33_ASAP7_75t_L g9246 ( 
.A(n_9087),
.B(n_4659),
.C(n_4490),
.Y(n_9246)
);

NOR4xp25_ASAP7_75t_L g9247 ( 
.A(n_9173),
.B(n_5106),
.C(n_4835),
.D(n_4434),
.Y(n_9247)
);

NAND2xp5_ASAP7_75t_L g9248 ( 
.A(n_9143),
.B(n_5260),
.Y(n_9248)
);

INVxp33_ASAP7_75t_SL g9249 ( 
.A(n_9178),
.Y(n_9249)
);

OAI21xp33_ASAP7_75t_SL g9250 ( 
.A1(n_9145),
.A2(n_4395),
.B(n_4426),
.Y(n_9250)
);

NOR2xp33_ASAP7_75t_L g9251 ( 
.A(n_9123),
.B(n_5260),
.Y(n_9251)
);

OAI21xp33_ASAP7_75t_SL g9252 ( 
.A1(n_9175),
.A2(n_4438),
.B(n_4873),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_9096),
.Y(n_9253)
);

BUFx2_ASAP7_75t_L g9254 ( 
.A(n_9169),
.Y(n_9254)
);

AOI211xp5_ASAP7_75t_L g9255 ( 
.A1(n_9163),
.A2(n_5263),
.B(n_4280),
.C(n_4401),
.Y(n_9255)
);

BUFx2_ASAP7_75t_L g9256 ( 
.A(n_9158),
.Y(n_9256)
);

OAI221xp5_ASAP7_75t_L g9257 ( 
.A1(n_9159),
.A2(n_5043),
.B1(n_4207),
.B2(n_4652),
.C(n_4648),
.Y(n_9257)
);

NAND3xp33_ASAP7_75t_SL g9258 ( 
.A(n_9154),
.B(n_4434),
.C(n_4558),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_9120),
.Y(n_9259)
);

O2A1O1Ixp33_ASAP7_75t_L g9260 ( 
.A1(n_9179),
.A2(n_4160),
.B(n_5043),
.C(n_4223),
.Y(n_9260)
);

NAND2xp5_ASAP7_75t_L g9261 ( 
.A(n_9160),
.B(n_5263),
.Y(n_9261)
);

NAND3xp33_ASAP7_75t_L g9262 ( 
.A(n_9155),
.B(n_4663),
.C(n_4657),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_9134),
.Y(n_9263)
);

OAI211xp5_ASAP7_75t_L g9264 ( 
.A1(n_9182),
.A2(n_4438),
.B(n_4937),
.C(n_4755),
.Y(n_9264)
);

BUFx2_ASAP7_75t_L g9265 ( 
.A(n_9180),
.Y(n_9265)
);

INVx1_ASAP7_75t_L g9266 ( 
.A(n_9136),
.Y(n_9266)
);

OAI211xp5_ASAP7_75t_L g9267 ( 
.A1(n_9099),
.A2(n_4438),
.B(n_4937),
.C(n_4755),
.Y(n_9267)
);

NAND4xp25_ASAP7_75t_L g9268 ( 
.A(n_9142),
.B(n_9126),
.C(n_9105),
.D(n_9184),
.Y(n_9268)
);

NAND2xp5_ASAP7_75t_L g9269 ( 
.A(n_9160),
.B(n_3981),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_9114),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_9122),
.Y(n_9271)
);

NAND2xp5_ASAP7_75t_L g9272 ( 
.A(n_9167),
.B(n_3981),
.Y(n_9272)
);

INVxp67_ASAP7_75t_SL g9273 ( 
.A(n_9121),
.Y(n_9273)
);

NAND2xp5_ASAP7_75t_SL g9274 ( 
.A(n_9109),
.B(n_4638),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_9124),
.Y(n_9275)
);

OAI211xp5_ASAP7_75t_SL g9276 ( 
.A1(n_9104),
.A2(n_4689),
.B(n_4743),
.C(n_4672),
.Y(n_9276)
);

AND4x1_ASAP7_75t_L g9277 ( 
.A(n_9128),
.B(n_4301),
.C(n_4562),
.D(n_4641),
.Y(n_9277)
);

AOI211x1_ASAP7_75t_L g9278 ( 
.A1(n_9101),
.A2(n_4870),
.B(n_4871),
.C(n_4866),
.Y(n_9278)
);

NAND2xp5_ASAP7_75t_L g9279 ( 
.A(n_9176),
.B(n_3981),
.Y(n_9279)
);

NAND2xp5_ASAP7_75t_L g9280 ( 
.A(n_9170),
.B(n_4885),
.Y(n_9280)
);

NAND2xp5_ASAP7_75t_SL g9281 ( 
.A(n_9103),
.B(n_4672),
.Y(n_9281)
);

OAI22xp5_ASAP7_75t_L g9282 ( 
.A1(n_9172),
.A2(n_4792),
.B1(n_4909),
.B2(n_4589),
.Y(n_9282)
);

AND3x4_ASAP7_75t_L g9283 ( 
.A(n_9177),
.B(n_4440),
.C(n_3801),
.Y(n_9283)
);

AOI21xp5_ASAP7_75t_L g9284 ( 
.A1(n_9151),
.A2(n_4870),
.B(n_4866),
.Y(n_9284)
);

NAND2xp5_ASAP7_75t_L g9285 ( 
.A(n_9147),
.B(n_4885),
.Y(n_9285)
);

NAND2xp5_ASAP7_75t_L g9286 ( 
.A(n_9171),
.B(n_3992),
.Y(n_9286)
);

XNOR2xp5_ASAP7_75t_L g9287 ( 
.A(n_9171),
.B(n_9150),
.Y(n_9287)
);

NOR4xp25_ASAP7_75t_SL g9288 ( 
.A(n_9157),
.B(n_4163),
.C(n_4148),
.D(n_4183),
.Y(n_9288)
);

AOI211xp5_ASAP7_75t_SL g9289 ( 
.A1(n_9152),
.A2(n_4689),
.B(n_4743),
.C(n_4672),
.Y(n_9289)
);

INVx2_ASAP7_75t_L g9290 ( 
.A(n_9204),
.Y(n_9290)
);

NOR3xp33_ASAP7_75t_L g9291 ( 
.A(n_9196),
.B(n_9137),
.C(n_9153),
.Y(n_9291)
);

NOR2xp33_ASAP7_75t_SL g9292 ( 
.A(n_9236),
.B(n_9164),
.Y(n_9292)
);

OAI21xp5_ASAP7_75t_L g9293 ( 
.A1(n_9191),
.A2(n_9161),
.B(n_9162),
.Y(n_9293)
);

NAND2xp5_ASAP7_75t_L g9294 ( 
.A(n_9240),
.B(n_9165),
.Y(n_9294)
);

NOR3xp33_ASAP7_75t_L g9295 ( 
.A(n_9187),
.B(n_9183),
.C(n_4534),
.Y(n_9295)
);

NAND3xp33_ASAP7_75t_L g9296 ( 
.A(n_9197),
.B(n_4530),
.C(n_4863),
.Y(n_9296)
);

NAND4xp25_ASAP7_75t_L g9297 ( 
.A(n_9218),
.B(n_9199),
.C(n_9186),
.D(n_9216),
.Y(n_9297)
);

NOR3x1_ASAP7_75t_L g9298 ( 
.A(n_9265),
.B(n_9254),
.C(n_9256),
.Y(n_9298)
);

NOR3x1_ASAP7_75t_L g9299 ( 
.A(n_9201),
.B(n_4152),
.C(n_4115),
.Y(n_9299)
);

NAND2xp5_ASAP7_75t_L g9300 ( 
.A(n_9198),
.B(n_3992),
.Y(n_9300)
);

INVx2_ASAP7_75t_SL g9301 ( 
.A(n_9226),
.Y(n_9301)
);

NAND2xp5_ASAP7_75t_L g9302 ( 
.A(n_9242),
.B(n_3992),
.Y(n_9302)
);

INVx2_ASAP7_75t_SL g9303 ( 
.A(n_9190),
.Y(n_9303)
);

NOR3xp33_ASAP7_75t_L g9304 ( 
.A(n_9192),
.B(n_4280),
.C(n_4441),
.Y(n_9304)
);

NOR2xp33_ASAP7_75t_L g9305 ( 
.A(n_9249),
.B(n_9189),
.Y(n_9305)
);

NAND4xp25_ASAP7_75t_L g9306 ( 
.A(n_9195),
.B(n_4394),
.C(n_4894),
.D(n_4875),
.Y(n_9306)
);

AOI211xp5_ASAP7_75t_L g9307 ( 
.A1(n_9193),
.A2(n_4441),
.B(n_3945),
.C(n_3900),
.Y(n_9307)
);

INVxp67_ASAP7_75t_L g9308 ( 
.A(n_9194),
.Y(n_9308)
);

NOR2xp33_ASAP7_75t_L g9309 ( 
.A(n_9212),
.B(n_3693),
.Y(n_9309)
);

NAND2xp5_ASAP7_75t_L g9310 ( 
.A(n_9200),
.B(n_3992),
.Y(n_9310)
);

HB1xp67_ASAP7_75t_L g9311 ( 
.A(n_9209),
.Y(n_9311)
);

NOR3xp33_ASAP7_75t_L g9312 ( 
.A(n_9245),
.B(n_4267),
.C(n_4274),
.Y(n_9312)
);

NAND2xp5_ASAP7_75t_L g9313 ( 
.A(n_9273),
.B(n_3992),
.Y(n_9313)
);

INVx1_ASAP7_75t_L g9314 ( 
.A(n_9210),
.Y(n_9314)
);

NAND3xp33_ASAP7_75t_SL g9315 ( 
.A(n_9229),
.B(n_9203),
.C(n_9231),
.Y(n_9315)
);

NAND2xp5_ASAP7_75t_L g9316 ( 
.A(n_9211),
.B(n_3992),
.Y(n_9316)
);

O2A1O1Ixp5_ASAP7_75t_L g9317 ( 
.A1(n_9188),
.A2(n_4743),
.B(n_4757),
.C(n_4689),
.Y(n_9317)
);

NAND3xp33_ASAP7_75t_SL g9318 ( 
.A(n_9244),
.B(n_9207),
.C(n_9202),
.Y(n_9318)
);

HB1xp67_ASAP7_75t_L g9319 ( 
.A(n_9253),
.Y(n_9319)
);

HB1xp67_ASAP7_75t_L g9320 ( 
.A(n_9214),
.Y(n_9320)
);

NOR2x1_ASAP7_75t_L g9321 ( 
.A(n_9185),
.B(n_4207),
.Y(n_9321)
);

NOR2x1_ASAP7_75t_L g9322 ( 
.A(n_9268),
.B(n_4292),
.Y(n_9322)
);

NAND2xp5_ASAP7_75t_L g9323 ( 
.A(n_9224),
.B(n_3992),
.Y(n_9323)
);

INVx1_ASAP7_75t_L g9324 ( 
.A(n_9221),
.Y(n_9324)
);

NOR2xp33_ASAP7_75t_L g9325 ( 
.A(n_9268),
.B(n_3710),
.Y(n_9325)
);

AND2x2_ASAP7_75t_L g9326 ( 
.A(n_9237),
.B(n_4557),
.Y(n_9326)
);

NAND2xp5_ASAP7_75t_SL g9327 ( 
.A(n_9243),
.B(n_4689),
.Y(n_9327)
);

NAND3xp33_ASAP7_75t_L g9328 ( 
.A(n_9275),
.B(n_5090),
.C(n_5084),
.Y(n_9328)
);

NOR2xp33_ASAP7_75t_SL g9329 ( 
.A(n_9263),
.B(n_3717),
.Y(n_9329)
);

NAND2xp5_ASAP7_75t_L g9330 ( 
.A(n_9227),
.B(n_4208),
.Y(n_9330)
);

NOR2xp33_ASAP7_75t_SL g9331 ( 
.A(n_9266),
.B(n_3717),
.Y(n_9331)
);

AND2x2_ASAP7_75t_L g9332 ( 
.A(n_9288),
.B(n_4557),
.Y(n_9332)
);

INVx1_ASAP7_75t_L g9333 ( 
.A(n_9271),
.Y(n_9333)
);

OAI221xp5_ASAP7_75t_L g9334 ( 
.A1(n_9250),
.A2(n_4626),
.B1(n_4584),
.B2(n_4792),
.C(n_4589),
.Y(n_9334)
);

NAND2xp5_ASAP7_75t_SL g9335 ( 
.A(n_9259),
.B(n_4743),
.Y(n_9335)
);

NOR3x1_ASAP7_75t_L g9336 ( 
.A(n_9228),
.B(n_4152),
.C(n_4115),
.Y(n_9336)
);

NAND2xp5_ASAP7_75t_L g9337 ( 
.A(n_9270),
.B(n_4208),
.Y(n_9337)
);

OR3x1_ASAP7_75t_L g9338 ( 
.A(n_9276),
.B(n_3882),
.C(n_4871),
.Y(n_9338)
);

INVx1_ASAP7_75t_L g9339 ( 
.A(n_9287),
.Y(n_9339)
);

INVx1_ASAP7_75t_L g9340 ( 
.A(n_9230),
.Y(n_9340)
);

OAI21xp33_ASAP7_75t_L g9341 ( 
.A1(n_9251),
.A2(n_4221),
.B(n_4153),
.Y(n_9341)
);

NAND3xp33_ASAP7_75t_L g9342 ( 
.A(n_9248),
.B(n_5055),
.C(n_4996),
.Y(n_9342)
);

AOI21xp5_ASAP7_75t_L g9343 ( 
.A1(n_9206),
.A2(n_4873),
.B(n_4872),
.Y(n_9343)
);

NAND2x1_ASAP7_75t_L g9344 ( 
.A(n_9241),
.B(n_4589),
.Y(n_9344)
);

OAI21xp33_ASAP7_75t_SL g9345 ( 
.A1(n_9232),
.A2(n_5102),
.B(n_4874),
.Y(n_9345)
);

NOR4xp25_ASAP7_75t_L g9346 ( 
.A(n_9239),
.B(n_4267),
.C(n_4874),
.D(n_4872),
.Y(n_9346)
);

AOI21xp5_ASAP7_75t_L g9347 ( 
.A1(n_9274),
.A2(n_9223),
.B(n_9235),
.Y(n_9347)
);

NOR4xp25_ASAP7_75t_L g9348 ( 
.A(n_9252),
.B(n_5079),
.C(n_5083),
.D(n_5076),
.Y(n_9348)
);

NOR2x1_ASAP7_75t_SL g9349 ( 
.A(n_9264),
.B(n_4585),
.Y(n_9349)
);

OAI211xp5_ASAP7_75t_L g9350 ( 
.A1(n_9288),
.A2(n_4937),
.B(n_5033),
.C(n_4755),
.Y(n_9350)
);

INVxp67_ASAP7_75t_L g9351 ( 
.A(n_9272),
.Y(n_9351)
);

NAND3xp33_ASAP7_75t_SL g9352 ( 
.A(n_9234),
.B(n_4626),
.C(n_4584),
.Y(n_9352)
);

NAND4xp75_ASAP7_75t_L g9353 ( 
.A(n_9205),
.B(n_4254),
.C(n_4301),
.D(n_4153),
.Y(n_9353)
);

NAND3xp33_ASAP7_75t_SL g9354 ( 
.A(n_9267),
.B(n_4626),
.C(n_4584),
.Y(n_9354)
);

NOR3xp33_ASAP7_75t_L g9355 ( 
.A(n_9279),
.B(n_4336),
.C(n_4274),
.Y(n_9355)
);

AOI21xp33_ASAP7_75t_L g9356 ( 
.A1(n_9286),
.A2(n_5055),
.B(n_4996),
.Y(n_9356)
);

NOR2xp67_ASAP7_75t_L g9357 ( 
.A(n_9261),
.B(n_4292),
.Y(n_9357)
);

NAND2xp5_ASAP7_75t_L g9358 ( 
.A(n_9278),
.B(n_4208),
.Y(n_9358)
);

NAND2xp5_ASAP7_75t_L g9359 ( 
.A(n_9233),
.B(n_4208),
.Y(n_9359)
);

INVxp67_ASAP7_75t_L g9360 ( 
.A(n_9269),
.Y(n_9360)
);

INVx2_ASAP7_75t_SL g9361 ( 
.A(n_9281),
.Y(n_9361)
);

NOR3x1_ASAP7_75t_L g9362 ( 
.A(n_9246),
.B(n_4221),
.C(n_4153),
.Y(n_9362)
);

NAND2xp5_ASAP7_75t_L g9363 ( 
.A(n_9247),
.B(n_4996),
.Y(n_9363)
);

NAND3xp33_ASAP7_75t_L g9364 ( 
.A(n_9289),
.B(n_9280),
.C(n_9220),
.Y(n_9364)
);

INVxp67_ASAP7_75t_SL g9365 ( 
.A(n_9262),
.Y(n_9365)
);

NAND4xp75_ASAP7_75t_L g9366 ( 
.A(n_9285),
.B(n_4254),
.C(n_4415),
.D(n_4221),
.Y(n_9366)
);

INVx1_ASAP7_75t_L g9367 ( 
.A(n_9283),
.Y(n_9367)
);

OAI221xp5_ASAP7_75t_SL g9368 ( 
.A1(n_9225),
.A2(n_4394),
.B1(n_4507),
.B2(n_5035),
.C(n_4928),
.Y(n_9368)
);

INVx2_ASAP7_75t_L g9369 ( 
.A(n_9219),
.Y(n_9369)
);

AND2x2_ASAP7_75t_L g9370 ( 
.A(n_9217),
.B(n_4585),
.Y(n_9370)
);

NOR3xp33_ASAP7_75t_L g9371 ( 
.A(n_9238),
.B(n_9258),
.C(n_9260),
.Y(n_9371)
);

AND2x2_ASAP7_75t_L g9372 ( 
.A(n_9215),
.B(n_4712),
.Y(n_9372)
);

NAND2xp33_ASAP7_75t_L g9373 ( 
.A(n_9282),
.B(n_9284),
.Y(n_9373)
);

INVx1_ASAP7_75t_L g9374 ( 
.A(n_9208),
.Y(n_9374)
);

NAND3xp33_ASAP7_75t_SL g9375 ( 
.A(n_9255),
.B(n_9213),
.C(n_9257),
.Y(n_9375)
);

NAND4xp25_ASAP7_75t_L g9376 ( 
.A(n_9222),
.B(n_4903),
.C(n_4457),
.D(n_4499),
.Y(n_9376)
);

NOR2xp33_ASAP7_75t_L g9377 ( 
.A(n_9277),
.B(n_5055),
.Y(n_9377)
);

AND3x4_ASAP7_75t_L g9378 ( 
.A(n_9207),
.B(n_4440),
.C(n_5074),
.Y(n_9378)
);

NOR2xp33_ASAP7_75t_L g9379 ( 
.A(n_9236),
.B(n_5057),
.Y(n_9379)
);

AOI21xp5_ASAP7_75t_L g9380 ( 
.A1(n_9187),
.A2(n_4878),
.B(n_4877),
.Y(n_9380)
);

NAND2xp5_ASAP7_75t_L g9381 ( 
.A(n_9236),
.B(n_5057),
.Y(n_9381)
);

AND2x2_ASAP7_75t_L g9382 ( 
.A(n_9204),
.B(n_4712),
.Y(n_9382)
);

NAND5xp2_ASAP7_75t_L g9383 ( 
.A(n_9236),
.B(n_4719),
.C(n_4781),
.D(n_4735),
.E(n_4678),
.Y(n_9383)
);

AOI221x1_ASAP7_75t_L g9384 ( 
.A1(n_9187),
.A2(n_5088),
.B1(n_5092),
.B2(n_5083),
.C(n_5079),
.Y(n_9384)
);

NAND2x1_ASAP7_75t_L g9385 ( 
.A(n_9265),
.B(n_4792),
.Y(n_9385)
);

NAND2xp5_ASAP7_75t_L g9386 ( 
.A(n_9236),
.B(n_5057),
.Y(n_9386)
);

NAND2xp5_ASAP7_75t_SL g9387 ( 
.A(n_9204),
.B(n_4757),
.Y(n_9387)
);

NAND3xp33_ASAP7_75t_L g9388 ( 
.A(n_9236),
.B(n_5099),
.C(n_5090),
.Y(n_9388)
);

INVxp67_ASAP7_75t_L g9389 ( 
.A(n_9236),
.Y(n_9389)
);

INVx1_ASAP7_75t_L g9390 ( 
.A(n_9187),
.Y(n_9390)
);

OAI22xp33_ASAP7_75t_L g9391 ( 
.A1(n_9197),
.A2(n_4988),
.B1(n_4909),
.B2(n_3907),
.Y(n_9391)
);

NOR2xp33_ASAP7_75t_SL g9392 ( 
.A(n_9236),
.B(n_4292),
.Y(n_9392)
);

NOR3xp33_ASAP7_75t_SL g9393 ( 
.A(n_9236),
.B(n_4429),
.C(n_4296),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_9187),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_9187),
.Y(n_9395)
);

NAND2xp5_ASAP7_75t_L g9396 ( 
.A(n_9389),
.B(n_9311),
.Y(n_9396)
);

INVxp67_ASAP7_75t_L g9397 ( 
.A(n_9305),
.Y(n_9397)
);

INVxp67_ASAP7_75t_SL g9398 ( 
.A(n_9298),
.Y(n_9398)
);

INVx1_ASAP7_75t_L g9399 ( 
.A(n_9319),
.Y(n_9399)
);

XOR2x2_ASAP7_75t_L g9400 ( 
.A(n_9385),
.B(n_4361),
.Y(n_9400)
);

INVxp67_ASAP7_75t_L g9401 ( 
.A(n_9292),
.Y(n_9401)
);

INVxp67_ASAP7_75t_SL g9402 ( 
.A(n_9290),
.Y(n_9402)
);

OAI22xp5_ASAP7_75t_L g9403 ( 
.A1(n_9303),
.A2(n_4988),
.B1(n_4909),
.B2(n_4757),
.Y(n_9403)
);

OAI211xp5_ASAP7_75t_L g9404 ( 
.A1(n_9297),
.A2(n_4937),
.B(n_5033),
.C(n_4755),
.Y(n_9404)
);

AOI322xp5_ASAP7_75t_L g9405 ( 
.A1(n_9318),
.A2(n_4639),
.A3(n_4934),
.B1(n_4947),
.B2(n_4800),
.C1(n_5063),
.C2(n_5061),
.Y(n_9405)
);

INVx1_ASAP7_75t_L g9406 ( 
.A(n_9301),
.Y(n_9406)
);

INVx1_ASAP7_75t_L g9407 ( 
.A(n_9314),
.Y(n_9407)
);

CKINVDCx20_ASAP7_75t_R g9408 ( 
.A(n_9395),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_9344),
.Y(n_9409)
);

OAI21xp33_ASAP7_75t_L g9410 ( 
.A1(n_9392),
.A2(n_4415),
.B(n_4440),
.Y(n_9410)
);

AOI22xp33_ASAP7_75t_L g9411 ( 
.A1(n_9339),
.A2(n_9315),
.B1(n_9291),
.B2(n_9308),
.Y(n_9411)
);

XNOR2x1_ASAP7_75t_L g9412 ( 
.A(n_9390),
.B(n_4507),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_9394),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_9320),
.Y(n_9414)
);

NAND2xp5_ASAP7_75t_SL g9415 ( 
.A(n_9333),
.B(n_4757),
.Y(n_9415)
);

INVx2_ASAP7_75t_L g9416 ( 
.A(n_9332),
.Y(n_9416)
);

NAND2xp5_ASAP7_75t_SL g9417 ( 
.A(n_9324),
.B(n_9322),
.Y(n_9417)
);

OAI21xp5_ASAP7_75t_L g9418 ( 
.A1(n_9294),
.A2(n_4191),
.B(n_4474),
.Y(n_9418)
);

AOI21xp33_ASAP7_75t_L g9419 ( 
.A1(n_9340),
.A2(n_5082),
.B(n_5077),
.Y(n_9419)
);

NAND2xp5_ASAP7_75t_L g9420 ( 
.A(n_9377),
.B(n_5077),
.Y(n_9420)
);

INVx1_ASAP7_75t_L g9421 ( 
.A(n_9363),
.Y(n_9421)
);

INVx1_ASAP7_75t_SL g9422 ( 
.A(n_9381),
.Y(n_9422)
);

AND2x2_ASAP7_75t_L g9423 ( 
.A(n_9382),
.B(n_4800),
.Y(n_9423)
);

NOR3x1_ASAP7_75t_L g9424 ( 
.A(n_9293),
.B(n_4415),
.C(n_4148),
.Y(n_9424)
);

NOR2x1_ASAP7_75t_L g9425 ( 
.A(n_9367),
.B(n_4292),
.Y(n_9425)
);

NOR2xp33_ASAP7_75t_L g9426 ( 
.A(n_9374),
.B(n_5077),
.Y(n_9426)
);

AOI22xp33_ASAP7_75t_L g9427 ( 
.A1(n_9365),
.A2(n_5090),
.B1(n_5099),
.B2(n_5082),
.Y(n_9427)
);

AOI221xp5_ASAP7_75t_SL g9428 ( 
.A1(n_9373),
.A2(n_4878),
.B1(n_4883),
.B2(n_4879),
.C(n_4877),
.Y(n_9428)
);

INVxp67_ASAP7_75t_SL g9429 ( 
.A(n_9361),
.Y(n_9429)
);

NAND2xp5_ASAP7_75t_L g9430 ( 
.A(n_9379),
.B(n_5082),
.Y(n_9430)
);

XOR2x2_ASAP7_75t_L g9431 ( 
.A(n_9378),
.B(n_4361),
.Y(n_9431)
);

NOR3x1_ASAP7_75t_L g9432 ( 
.A(n_9387),
.B(n_4163),
.C(n_4183),
.Y(n_9432)
);

NAND2xp5_ASAP7_75t_L g9433 ( 
.A(n_9357),
.B(n_5084),
.Y(n_9433)
);

NAND2x1p5_ASAP7_75t_L g9434 ( 
.A(n_9369),
.B(n_4297),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_9386),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_9300),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_9321),
.Y(n_9437)
);

O2A1O1Ixp33_ASAP7_75t_L g9438 ( 
.A1(n_9360),
.A2(n_4692),
.B(n_4719),
.C(n_4678),
.Y(n_9438)
);

NAND2x1_ASAP7_75t_SL g9439 ( 
.A(n_9325),
.B(n_4851),
.Y(n_9439)
);

NOR2xp33_ASAP7_75t_L g9440 ( 
.A(n_9364),
.B(n_5084),
.Y(n_9440)
);

AOI22xp5_ASAP7_75t_L g9441 ( 
.A1(n_9295),
.A2(n_4988),
.B1(n_4510),
.B2(n_4941),
.Y(n_9441)
);

AOI22xp33_ASAP7_75t_L g9442 ( 
.A1(n_9371),
.A2(n_5099),
.B1(n_5108),
.B2(n_3907),
.Y(n_9442)
);

XNOR2xp5_ASAP7_75t_L g9443 ( 
.A(n_9375),
.B(n_4507),
.Y(n_9443)
);

NAND2xp5_ASAP7_75t_L g9444 ( 
.A(n_9370),
.B(n_5108),
.Y(n_9444)
);

INVx1_ASAP7_75t_L g9445 ( 
.A(n_9313),
.Y(n_9445)
);

NAND3xp33_ASAP7_75t_L g9446 ( 
.A(n_9351),
.B(n_9347),
.C(n_9331),
.Y(n_9446)
);

AOI22xp5_ASAP7_75t_L g9447 ( 
.A1(n_9329),
.A2(n_4988),
.B1(n_4510),
.B2(n_4941),
.Y(n_9447)
);

NAND3xp33_ASAP7_75t_SL g9448 ( 
.A(n_9309),
.B(n_4984),
.C(n_4973),
.Y(n_9448)
);

HB1xp67_ASAP7_75t_L g9449 ( 
.A(n_9335),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_9316),
.Y(n_9450)
);

A2O1A1Ixp33_ASAP7_75t_L g9451 ( 
.A1(n_9317),
.A2(n_9345),
.B(n_9330),
.C(n_9341),
.Y(n_9451)
);

OAI21xp33_ASAP7_75t_SL g9452 ( 
.A1(n_9327),
.A2(n_5051),
.B(n_5050),
.Y(n_9452)
);

NAND2x1_ASAP7_75t_L g9453 ( 
.A(n_9326),
.B(n_4297),
.Y(n_9453)
);

HB1xp67_ASAP7_75t_L g9454 ( 
.A(n_9302),
.Y(n_9454)
);

INVx1_ASAP7_75t_SL g9455 ( 
.A(n_9310),
.Y(n_9455)
);

OAI21xp33_ASAP7_75t_L g9456 ( 
.A1(n_9350),
.A2(n_5087),
.B(n_5058),
.Y(n_9456)
);

INVx2_ASAP7_75t_SL g9457 ( 
.A(n_9337),
.Y(n_9457)
);

INVx2_ASAP7_75t_L g9458 ( 
.A(n_9338),
.Y(n_9458)
);

OAI21xp33_ASAP7_75t_SL g9459 ( 
.A1(n_9353),
.A2(n_5051),
.B(n_5050),
.Y(n_9459)
);

A2O1A1Ixp33_ASAP7_75t_L g9460 ( 
.A1(n_9359),
.A2(n_4916),
.B(n_4942),
.C(n_4883),
.Y(n_9460)
);

NAND2xp5_ASAP7_75t_SL g9461 ( 
.A(n_9391),
.B(n_4851),
.Y(n_9461)
);

INVx1_ASAP7_75t_SL g9462 ( 
.A(n_9323),
.Y(n_9462)
);

OAI22xp5_ASAP7_75t_L g9463 ( 
.A1(n_9366),
.A2(n_5087),
.B1(n_5058),
.B2(n_4941),
.Y(n_9463)
);

INVx1_ASAP7_75t_L g9464 ( 
.A(n_9362),
.Y(n_9464)
);

OAI21xp33_ASAP7_75t_L g9465 ( 
.A1(n_9304),
.A2(n_5087),
.B(n_5058),
.Y(n_9465)
);

INVx1_ASAP7_75t_L g9466 ( 
.A(n_9358),
.Y(n_9466)
);

INVxp67_ASAP7_75t_L g9467 ( 
.A(n_9388),
.Y(n_9467)
);

NAND2x1p5_ASAP7_75t_L g9468 ( 
.A(n_9299),
.B(n_4297),
.Y(n_9468)
);

INVxp67_ASAP7_75t_L g9469 ( 
.A(n_9349),
.Y(n_9469)
);

XNOR2x1_ASAP7_75t_L g9470 ( 
.A(n_9372),
.B(n_4507),
.Y(n_9470)
);

INVx1_ASAP7_75t_L g9471 ( 
.A(n_9336),
.Y(n_9471)
);

AOI221xp5_ASAP7_75t_SL g9472 ( 
.A1(n_9380),
.A2(n_4884),
.B1(n_4895),
.B2(n_4888),
.C(n_4879),
.Y(n_9472)
);

AOI221xp5_ASAP7_75t_L g9473 ( 
.A1(n_9348),
.A2(n_3900),
.B1(n_3931),
.B2(n_3929),
.C(n_3907),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_9355),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_9402),
.Y(n_9475)
);

AOI22xp5_ASAP7_75t_L g9476 ( 
.A1(n_9399),
.A2(n_9296),
.B1(n_9312),
.B2(n_9354),
.Y(n_9476)
);

AOI221xp5_ASAP7_75t_L g9477 ( 
.A1(n_9401),
.A2(n_9346),
.B1(n_9356),
.B2(n_9343),
.C(n_9352),
.Y(n_9477)
);

INVx1_ASAP7_75t_L g9478 ( 
.A(n_9396),
.Y(n_9478)
);

AOI221xp5_ASAP7_75t_L g9479 ( 
.A1(n_9397),
.A2(n_9328),
.B1(n_9306),
.B2(n_9342),
.C(n_9368),
.Y(n_9479)
);

AOI22xp5_ASAP7_75t_L g9480 ( 
.A1(n_9414),
.A2(n_9342),
.B1(n_9393),
.B2(n_9376),
.Y(n_9480)
);

AOI31xp33_ASAP7_75t_L g9481 ( 
.A1(n_9429),
.A2(n_9307),
.A3(n_9334),
.B(n_9383),
.Y(n_9481)
);

NOR2xp33_ASAP7_75t_SL g9482 ( 
.A(n_9398),
.B(n_9307),
.Y(n_9482)
);

INVx2_ASAP7_75t_L g9483 ( 
.A(n_9408),
.Y(n_9483)
);

NAND2xp5_ASAP7_75t_L g9484 ( 
.A(n_9411),
.B(n_9384),
.Y(n_9484)
);

INVx1_ASAP7_75t_L g9485 ( 
.A(n_9413),
.Y(n_9485)
);

INVx1_ASAP7_75t_L g9486 ( 
.A(n_9407),
.Y(n_9486)
);

NAND4xp25_ASAP7_75t_L g9487 ( 
.A(n_9446),
.B(n_5008),
.C(n_4230),
.D(n_4311),
.Y(n_9487)
);

AOI22xp5_ASAP7_75t_L g9488 ( 
.A1(n_9416),
.A2(n_4851),
.B1(n_5007),
.B2(n_4941),
.Y(n_9488)
);

NOR2xp33_ASAP7_75t_L g9489 ( 
.A(n_9469),
.B(n_5108),
.Y(n_9489)
);

NAND2xp5_ASAP7_75t_L g9490 ( 
.A(n_9421),
.B(n_4675),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_9406),
.Y(n_9491)
);

HB1xp67_ASAP7_75t_L g9492 ( 
.A(n_9409),
.Y(n_9492)
);

BUFx2_ASAP7_75t_L g9493 ( 
.A(n_9439),
.Y(n_9493)
);

NAND2xp5_ASAP7_75t_L g9494 ( 
.A(n_9422),
.B(n_4675),
.Y(n_9494)
);

AO22x2_ASAP7_75t_L g9495 ( 
.A1(n_9458),
.A2(n_4182),
.B1(n_4888),
.B2(n_4884),
.Y(n_9495)
);

INVx2_ASAP7_75t_L g9496 ( 
.A(n_9468),
.Y(n_9496)
);

NOR2x1_ASAP7_75t_L g9497 ( 
.A(n_9417),
.B(n_4297),
.Y(n_9497)
);

INVx1_ASAP7_75t_L g9498 ( 
.A(n_9412),
.Y(n_9498)
);

INVx1_ASAP7_75t_L g9499 ( 
.A(n_9444),
.Y(n_9499)
);

INVx1_ASAP7_75t_L g9500 ( 
.A(n_9437),
.Y(n_9500)
);

NOR2xp33_ASAP7_75t_L g9501 ( 
.A(n_9453),
.B(n_4427),
.Y(n_9501)
);

AOI22xp5_ASAP7_75t_L g9502 ( 
.A1(n_9464),
.A2(n_4851),
.B1(n_5087),
.B2(n_5058),
.Y(n_9502)
);

NOR4xp25_ASAP7_75t_L g9503 ( 
.A(n_9462),
.B(n_5007),
.C(n_4905),
.D(n_4906),
.Y(n_9503)
);

INVx1_ASAP7_75t_L g9504 ( 
.A(n_9434),
.Y(n_9504)
);

NOR2x1_ASAP7_75t_L g9505 ( 
.A(n_9435),
.B(n_5007),
.Y(n_9505)
);

AOI31xp33_ASAP7_75t_L g9506 ( 
.A1(n_9449),
.A2(n_4678),
.A3(n_4719),
.B(n_4692),
.Y(n_9506)
);

INVx1_ASAP7_75t_L g9507 ( 
.A(n_9420),
.Y(n_9507)
);

INVx1_ASAP7_75t_L g9508 ( 
.A(n_9443),
.Y(n_9508)
);

AOI22xp5_ASAP7_75t_L g9509 ( 
.A1(n_9467),
.A2(n_5007),
.B1(n_4510),
.B2(n_3983),
.Y(n_9509)
);

AOI22xp5_ASAP7_75t_L g9510 ( 
.A1(n_9440),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9510)
);

INVxp67_ASAP7_75t_SL g9511 ( 
.A(n_9454),
.Y(n_9511)
);

AO211x2_ASAP7_75t_L g9512 ( 
.A1(n_9471),
.A2(n_4336),
.B(n_4230),
.C(n_4895),
.Y(n_9512)
);

INVx1_ASAP7_75t_L g9513 ( 
.A(n_9433),
.Y(n_9513)
);

INVx1_ASAP7_75t_L g9514 ( 
.A(n_9426),
.Y(n_9514)
);

AO22x2_ASAP7_75t_L g9515 ( 
.A1(n_9455),
.A2(n_4182),
.B1(n_4906),
.B2(n_4905),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_9424),
.Y(n_9516)
);

INVx1_ASAP7_75t_L g9517 ( 
.A(n_9415),
.Y(n_9517)
);

NAND2xp5_ASAP7_75t_L g9518 ( 
.A(n_9457),
.B(n_4694),
.Y(n_9518)
);

AO22x1_ASAP7_75t_L g9519 ( 
.A1(n_9425),
.A2(n_3868),
.B1(n_3870),
.B2(n_4337),
.Y(n_9519)
);

AOI22xp5_ASAP7_75t_L g9520 ( 
.A1(n_9436),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9520)
);

NOR4xp25_ASAP7_75t_L g9521 ( 
.A(n_9466),
.B(n_4916),
.C(n_4923),
.D(n_4912),
.Y(n_9521)
);

AO22x2_ASAP7_75t_L g9522 ( 
.A1(n_9445),
.A2(n_9450),
.B1(n_9474),
.B2(n_9404),
.Y(n_9522)
);

AOI22xp5_ASAP7_75t_L g9523 ( 
.A1(n_9459),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9523)
);

AO22x1_ASAP7_75t_L g9524 ( 
.A1(n_9432),
.A2(n_3868),
.B1(n_3870),
.B2(n_4337),
.Y(n_9524)
);

NOR4xp25_ASAP7_75t_L g9525 ( 
.A(n_9451),
.B(n_4923),
.C(n_4925),
.D(n_4912),
.Y(n_9525)
);

NOR4xp25_ASAP7_75t_L g9526 ( 
.A(n_9459),
.B(n_4931),
.C(n_4938),
.D(n_4925),
.Y(n_9526)
);

NOR3xp33_ASAP7_75t_L g9527 ( 
.A(n_9430),
.B(n_4408),
.C(n_4474),
.Y(n_9527)
);

NOR2x1_ASAP7_75t_L g9528 ( 
.A(n_9460),
.B(n_4931),
.Y(n_9528)
);

INVx1_ASAP7_75t_L g9529 ( 
.A(n_9431),
.Y(n_9529)
);

INVx1_ASAP7_75t_L g9530 ( 
.A(n_9400),
.Y(n_9530)
);

INVx2_ASAP7_75t_L g9531 ( 
.A(n_9470),
.Y(n_9531)
);

OAI22xp5_ASAP7_75t_L g9532 ( 
.A1(n_9441),
.A2(n_4942),
.B1(n_4948),
.B2(n_4938),
.Y(n_9532)
);

INVx1_ASAP7_75t_L g9533 ( 
.A(n_9452),
.Y(n_9533)
);

AOI22xp5_ASAP7_75t_L g9534 ( 
.A1(n_9423),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9534)
);

AOI22xp5_ASAP7_75t_L g9535 ( 
.A1(n_9442),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9535)
);

NOR4xp25_ASAP7_75t_L g9536 ( 
.A(n_9452),
.B(n_4952),
.C(n_4954),
.D(n_4948),
.Y(n_9536)
);

NOR2x1_ASAP7_75t_L g9537 ( 
.A(n_9461),
.B(n_4952),
.Y(n_9537)
);

AOI22xp5_ASAP7_75t_L g9538 ( 
.A1(n_9418),
.A2(n_4510),
.B1(n_3983),
.B2(n_4033),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_9465),
.Y(n_9539)
);

NAND3xp33_ASAP7_75t_SL g9540 ( 
.A(n_9483),
.B(n_9447),
.C(n_9456),
.Y(n_9540)
);

OAI21xp5_ASAP7_75t_L g9541 ( 
.A1(n_9511),
.A2(n_9419),
.B(n_9448),
.Y(n_9541)
);

NOR3xp33_ASAP7_75t_L g9542 ( 
.A(n_9478),
.B(n_9403),
.C(n_9410),
.Y(n_9542)
);

INVxp67_ASAP7_75t_L g9543 ( 
.A(n_9492),
.Y(n_9543)
);

INVx1_ASAP7_75t_L g9544 ( 
.A(n_9493),
.Y(n_9544)
);

NAND2xp5_ASAP7_75t_SL g9545 ( 
.A(n_9475),
.B(n_9428),
.Y(n_9545)
);

INVx1_ASAP7_75t_SL g9546 ( 
.A(n_9485),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_9486),
.Y(n_9547)
);

INVx1_ASAP7_75t_L g9548 ( 
.A(n_9484),
.Y(n_9548)
);

NAND3xp33_ASAP7_75t_L g9549 ( 
.A(n_9482),
.B(n_9427),
.C(n_9472),
.Y(n_9549)
);

INVxp67_ASAP7_75t_SL g9550 ( 
.A(n_9491),
.Y(n_9550)
);

NAND2xp5_ASAP7_75t_L g9551 ( 
.A(n_9500),
.B(n_9473),
.Y(n_9551)
);

NAND3xp33_ASAP7_75t_L g9552 ( 
.A(n_9504),
.B(n_9405),
.C(n_9438),
.Y(n_9552)
);

NOR2xp67_ASAP7_75t_L g9553 ( 
.A(n_9480),
.B(n_9463),
.Y(n_9553)
);

NAND2xp5_ASAP7_75t_L g9554 ( 
.A(n_9496),
.B(n_4694),
.Y(n_9554)
);

O2A1O1Ixp33_ASAP7_75t_SL g9555 ( 
.A1(n_9516),
.A2(n_5065),
.B(n_5076),
.C(n_5053),
.Y(n_9555)
);

AOI21xp33_ASAP7_75t_L g9556 ( 
.A1(n_9513),
.A2(n_9499),
.B(n_9507),
.Y(n_9556)
);

NOR2x1_ASAP7_75t_L g9557 ( 
.A(n_9533),
.B(n_5074),
.Y(n_9557)
);

OR2x2_ASAP7_75t_L g9558 ( 
.A(n_9494),
.B(n_4427),
.Y(n_9558)
);

OR2x2_ASAP7_75t_L g9559 ( 
.A(n_9514),
.B(n_4015),
.Y(n_9559)
);

NOR3xp33_ASAP7_75t_L g9560 ( 
.A(n_9508),
.B(n_3879),
.C(n_3848),
.Y(n_9560)
);

NAND2xp5_ASAP7_75t_SL g9561 ( 
.A(n_9477),
.B(n_3900),
.Y(n_9561)
);

NAND2xp5_ASAP7_75t_SL g9562 ( 
.A(n_9479),
.B(n_9476),
.Y(n_9562)
);

NAND3xp33_ASAP7_75t_L g9563 ( 
.A(n_9530),
.B(n_3907),
.C(n_3900),
.Y(n_9563)
);

NAND2xp5_ASAP7_75t_L g9564 ( 
.A(n_9531),
.B(n_4710),
.Y(n_9564)
);

AND2x2_ASAP7_75t_L g9565 ( 
.A(n_9497),
.B(n_5101),
.Y(n_9565)
);

NOR2x1_ASAP7_75t_L g9566 ( 
.A(n_9517),
.B(n_5101),
.Y(n_9566)
);

AOI21xp33_ASAP7_75t_L g9567 ( 
.A1(n_9498),
.A2(n_9529),
.B(n_9522),
.Y(n_9567)
);

NAND2xp5_ASAP7_75t_L g9568 ( 
.A(n_9522),
.B(n_4710),
.Y(n_9568)
);

AND2x2_ASAP7_75t_L g9569 ( 
.A(n_9501),
.B(n_5101),
.Y(n_9569)
);

NAND2xp5_ASAP7_75t_L g9570 ( 
.A(n_9505),
.B(n_4796),
.Y(n_9570)
);

INVxp67_ASAP7_75t_L g9571 ( 
.A(n_9489),
.Y(n_9571)
);

NAND3xp33_ASAP7_75t_L g9572 ( 
.A(n_9539),
.B(n_3907),
.C(n_3900),
.Y(n_9572)
);

AND3x1_ASAP7_75t_L g9573 ( 
.A(n_9525),
.B(n_4145),
.C(n_4136),
.Y(n_9573)
);

NAND2x1p5_ASAP7_75t_L g9574 ( 
.A(n_9537),
.B(n_3912),
.Y(n_9574)
);

NAND2xp33_ASAP7_75t_L g9575 ( 
.A(n_9528),
.B(n_4937),
.Y(n_9575)
);

NOR2x1p5_ASAP7_75t_L g9576 ( 
.A(n_9518),
.B(n_4136),
.Y(n_9576)
);

NOR2xp33_ASAP7_75t_L g9577 ( 
.A(n_9481),
.B(n_9490),
.Y(n_9577)
);

NAND2xp5_ASAP7_75t_L g9578 ( 
.A(n_9503),
.B(n_4796),
.Y(n_9578)
);

NAND2xp5_ASAP7_75t_L g9579 ( 
.A(n_9526),
.B(n_4807),
.Y(n_9579)
);

INVx1_ASAP7_75t_SL g9580 ( 
.A(n_9524),
.Y(n_9580)
);

NAND3xp33_ASAP7_75t_L g9581 ( 
.A(n_9487),
.B(n_3907),
.C(n_3900),
.Y(n_9581)
);

NAND2xp5_ASAP7_75t_SL g9582 ( 
.A(n_9488),
.B(n_3907),
.Y(n_9582)
);

NOR2xp33_ASAP7_75t_L g9583 ( 
.A(n_9532),
.B(n_4807),
.Y(n_9583)
);

NAND2xp5_ASAP7_75t_SL g9584 ( 
.A(n_9520),
.B(n_3929),
.Y(n_9584)
);

BUFx3_ASAP7_75t_L g9585 ( 
.A(n_9515),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_9512),
.Y(n_9586)
);

INVx1_ASAP7_75t_L g9587 ( 
.A(n_9515),
.Y(n_9587)
);

NAND2xp5_ASAP7_75t_SL g9588 ( 
.A(n_9509),
.B(n_3929),
.Y(n_9588)
);

AOI22xp5_ASAP7_75t_L g9589 ( 
.A1(n_9538),
.A2(n_4033),
.B1(n_4045),
.B2(n_3976),
.Y(n_9589)
);

AND2x2_ASAP7_75t_L g9590 ( 
.A(n_9536),
.B(n_5101),
.Y(n_9590)
);

INVx1_ASAP7_75t_L g9591 ( 
.A(n_9521),
.Y(n_9591)
);

NAND2xp5_ASAP7_75t_SL g9592 ( 
.A(n_9523),
.B(n_3929),
.Y(n_9592)
);

OR2x2_ASAP7_75t_L g9593 ( 
.A(n_9543),
.B(n_9519),
.Y(n_9593)
);

NOR3xp33_ASAP7_75t_L g9594 ( 
.A(n_9567),
.B(n_9527),
.C(n_9506),
.Y(n_9594)
);

NAND4xp75_ASAP7_75t_L g9595 ( 
.A(n_9544),
.B(n_9502),
.C(n_9510),
.D(n_9534),
.Y(n_9595)
);

NOR2x1_ASAP7_75t_L g9596 ( 
.A(n_9547),
.B(n_9495),
.Y(n_9596)
);

AOI221xp5_ASAP7_75t_L g9597 ( 
.A1(n_9550),
.A2(n_9495),
.B1(n_9535),
.B2(n_3929),
.C(n_3931),
.Y(n_9597)
);

NOR3xp33_ASAP7_75t_L g9598 ( 
.A(n_9556),
.B(n_3879),
.C(n_3848),
.Y(n_9598)
);

NAND4xp75_ASAP7_75t_L g9599 ( 
.A(n_9562),
.B(n_4956),
.C(n_4957),
.D(n_4954),
.Y(n_9599)
);

NOR2x1_ASAP7_75t_SL g9600 ( 
.A(n_9545),
.B(n_3803),
.Y(n_9600)
);

BUFx6f_ASAP7_75t_L g9601 ( 
.A(n_9548),
.Y(n_9601)
);

NOR3xp33_ASAP7_75t_L g9602 ( 
.A(n_9546),
.B(n_3879),
.C(n_3848),
.Y(n_9602)
);

NOR3x1_ASAP7_75t_L g9603 ( 
.A(n_9541),
.B(n_4286),
.C(n_4186),
.Y(n_9603)
);

NAND3xp33_ASAP7_75t_SL g9604 ( 
.A(n_9577),
.B(n_4311),
.C(n_4692),
.Y(n_9604)
);

AND3x4_ASAP7_75t_L g9605 ( 
.A(n_9542),
.B(n_3755),
.C(n_4118),
.Y(n_9605)
);

NAND3x1_ASAP7_75t_SL g9606 ( 
.A(n_9557),
.B(n_3755),
.C(n_3832),
.Y(n_9606)
);

INVx2_ASAP7_75t_SL g9607 ( 
.A(n_9568),
.Y(n_9607)
);

NOR3xp33_ASAP7_75t_L g9608 ( 
.A(n_9571),
.B(n_9551),
.C(n_9553),
.Y(n_9608)
);

NAND2xp5_ASAP7_75t_SL g9609 ( 
.A(n_9586),
.B(n_3929),
.Y(n_9609)
);

NAND3xp33_ASAP7_75t_L g9610 ( 
.A(n_9591),
.B(n_3931),
.C(n_3929),
.Y(n_9610)
);

NAND4xp25_ASAP7_75t_L g9611 ( 
.A(n_9552),
.B(n_4444),
.C(n_4269),
.D(n_4276),
.Y(n_9611)
);

AND3x4_ASAP7_75t_L g9612 ( 
.A(n_9566),
.B(n_4119),
.C(n_4118),
.Y(n_9612)
);

AND2x4_ASAP7_75t_SL g9613 ( 
.A(n_9565),
.B(n_3915),
.Y(n_9613)
);

AND2x4_ASAP7_75t_L g9614 ( 
.A(n_9549),
.B(n_4186),
.Y(n_9614)
);

NOR2x1_ASAP7_75t_L g9615 ( 
.A(n_9585),
.B(n_4956),
.Y(n_9615)
);

NAND3xp33_ASAP7_75t_L g9616 ( 
.A(n_9587),
.B(n_3931),
.C(n_3976),
.Y(n_9616)
);

NAND3xp33_ASAP7_75t_SL g9617 ( 
.A(n_9580),
.B(n_9564),
.C(n_9561),
.Y(n_9617)
);

NAND2xp5_ASAP7_75t_L g9618 ( 
.A(n_9559),
.B(n_4814),
.Y(n_9618)
);

NOR2xp33_ASAP7_75t_L g9619 ( 
.A(n_9540),
.B(n_9554),
.Y(n_9619)
);

INVx2_ASAP7_75t_SL g9620 ( 
.A(n_9576),
.Y(n_9620)
);

NOR2x1_ASAP7_75t_L g9621 ( 
.A(n_9575),
.B(n_4957),
.Y(n_9621)
);

NOR4xp25_ASAP7_75t_L g9622 ( 
.A(n_9563),
.B(n_4965),
.C(n_4966),
.D(n_4959),
.Y(n_9622)
);

OR2x2_ASAP7_75t_L g9623 ( 
.A(n_9558),
.B(n_4015),
.Y(n_9623)
);

NAND2xp5_ASAP7_75t_L g9624 ( 
.A(n_9570),
.B(n_9574),
.Y(n_9624)
);

NAND3x1_ASAP7_75t_L g9625 ( 
.A(n_9590),
.B(n_4145),
.C(n_4136),
.Y(n_9625)
);

NOR3xp33_ASAP7_75t_L g9626 ( 
.A(n_9578),
.B(n_3879),
.C(n_3848),
.Y(n_9626)
);

NOR2x1p5_ASAP7_75t_L g9627 ( 
.A(n_9579),
.B(n_9569),
.Y(n_9627)
);

NAND4xp25_ASAP7_75t_L g9628 ( 
.A(n_9560),
.B(n_4255),
.C(n_4281),
.D(n_4283),
.Y(n_9628)
);

AND4x1_ASAP7_75t_L g9629 ( 
.A(n_9572),
.B(n_9581),
.C(n_9583),
.D(n_9573),
.Y(n_9629)
);

NAND3xp33_ASAP7_75t_L g9630 ( 
.A(n_9573),
.B(n_9592),
.C(n_9584),
.Y(n_9630)
);

NOR3xp33_ASAP7_75t_L g9631 ( 
.A(n_9582),
.B(n_3879),
.C(n_3848),
.Y(n_9631)
);

INVx1_ASAP7_75t_SL g9632 ( 
.A(n_9588),
.Y(n_9632)
);

NAND3xp33_ASAP7_75t_L g9633 ( 
.A(n_9555),
.B(n_3931),
.C(n_3976),
.Y(n_9633)
);

NAND4xp25_ASAP7_75t_L g9634 ( 
.A(n_9589),
.B(n_4231),
.C(n_4360),
.D(n_4316),
.Y(n_9634)
);

OR2x2_ASAP7_75t_L g9635 ( 
.A(n_9543),
.B(n_4021),
.Y(n_9635)
);

NOR2x1_ASAP7_75t_L g9636 ( 
.A(n_9544),
.B(n_4959),
.Y(n_9636)
);

NOR3x1_ASAP7_75t_L g9637 ( 
.A(n_9550),
.B(n_4437),
.C(n_4286),
.Y(n_9637)
);

INVx1_ASAP7_75t_L g9638 ( 
.A(n_9550),
.Y(n_9638)
);

AND5x1_ASAP7_75t_L g9639 ( 
.A(n_9577),
.B(n_4364),
.C(n_4258),
.D(n_4383),
.E(n_4245),
.Y(n_9639)
);

INVx1_ASAP7_75t_L g9640 ( 
.A(n_9601),
.Y(n_9640)
);

INVx1_ASAP7_75t_L g9641 ( 
.A(n_9601),
.Y(n_9641)
);

INVx2_ASAP7_75t_L g9642 ( 
.A(n_9601),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_9638),
.Y(n_9643)
);

NOR3xp33_ASAP7_75t_L g9644 ( 
.A(n_9608),
.B(n_3899),
.C(n_3884),
.Y(n_9644)
);

AND2x4_ASAP7_75t_L g9645 ( 
.A(n_9627),
.B(n_4437),
.Y(n_9645)
);

OAI221xp5_ASAP7_75t_SL g9646 ( 
.A1(n_9594),
.A2(n_4299),
.B1(n_4293),
.B2(n_4966),
.C(n_4965),
.Y(n_9646)
);

AND2x2_ASAP7_75t_L g9647 ( 
.A(n_9603),
.B(n_4968),
.Y(n_9647)
);

OR2x2_ASAP7_75t_L g9648 ( 
.A(n_9635),
.B(n_4053),
.Y(n_9648)
);

AND2x4_ASAP7_75t_L g9649 ( 
.A(n_9614),
.B(n_4136),
.Y(n_9649)
);

NOR3xp33_ASAP7_75t_L g9650 ( 
.A(n_9607),
.B(n_3899),
.C(n_3884),
.Y(n_9650)
);

OAI311xp33_ASAP7_75t_L g9651 ( 
.A1(n_9593),
.A2(n_4144),
.A3(n_4104),
.B1(n_4021),
.C1(n_4968),
.Y(n_9651)
);

NOR3xp33_ASAP7_75t_L g9652 ( 
.A(n_9619),
.B(n_3899),
.C(n_3884),
.Y(n_9652)
);

OA22x2_ASAP7_75t_L g9653 ( 
.A1(n_9614),
.A2(n_4975),
.B1(n_4985),
.B2(n_4970),
.Y(n_9653)
);

NAND2xp33_ASAP7_75t_SL g9654 ( 
.A(n_9620),
.B(n_3906),
.Y(n_9654)
);

OAI211xp5_ASAP7_75t_L g9655 ( 
.A1(n_9596),
.A2(n_5044),
.B(n_5033),
.C(n_5092),
.Y(n_9655)
);

AOI22xp33_ASAP7_75t_SL g9656 ( 
.A1(n_9600),
.A2(n_4034),
.B1(n_4095),
.B2(n_3931),
.Y(n_9656)
);

AND2x4_ASAP7_75t_L g9657 ( 
.A(n_9613),
.B(n_9636),
.Y(n_9657)
);

NOR2x1_ASAP7_75t_L g9658 ( 
.A(n_9617),
.B(n_4970),
.Y(n_9658)
);

NOR2x1_ASAP7_75t_L g9659 ( 
.A(n_9624),
.B(n_4975),
.Y(n_9659)
);

NAND3xp33_ASAP7_75t_SL g9660 ( 
.A(n_9632),
.B(n_4781),
.C(n_4735),
.Y(n_9660)
);

INVx2_ASAP7_75t_L g9661 ( 
.A(n_9615),
.Y(n_9661)
);

AOI21xp5_ASAP7_75t_L g9662 ( 
.A1(n_9609),
.A2(n_4986),
.B(n_4985),
.Y(n_9662)
);

OR2x2_ASAP7_75t_L g9663 ( 
.A(n_9623),
.B(n_4053),
.Y(n_9663)
);

NOR3xp33_ASAP7_75t_L g9664 ( 
.A(n_9595),
.B(n_3899),
.C(n_3884),
.Y(n_9664)
);

NOR2xp33_ASAP7_75t_L g9665 ( 
.A(n_9629),
.B(n_4021),
.Y(n_9665)
);

NOR3xp33_ASAP7_75t_L g9666 ( 
.A(n_9630),
.B(n_9606),
.C(n_9616),
.Y(n_9666)
);

HB1xp67_ASAP7_75t_L g9667 ( 
.A(n_9610),
.Y(n_9667)
);

OAI22xp33_ASAP7_75t_L g9668 ( 
.A1(n_9597),
.A2(n_3931),
.B1(n_5032),
.B2(n_5020),
.Y(n_9668)
);

INVx2_ASAP7_75t_L g9669 ( 
.A(n_9625),
.Y(n_9669)
);

NOR2xp33_ASAP7_75t_L g9670 ( 
.A(n_9618),
.B(n_9612),
.Y(n_9670)
);

AOI221x1_ASAP7_75t_L g9671 ( 
.A1(n_9626),
.A2(n_4997),
.B1(n_4998),
.B2(n_4994),
.C(n_4986),
.Y(n_9671)
);

NOR2xp33_ASAP7_75t_L g9672 ( 
.A(n_9621),
.B(n_4104),
.Y(n_9672)
);

NOR3x2_ASAP7_75t_L g9673 ( 
.A(n_9599),
.B(n_4144),
.C(n_4104),
.Y(n_9673)
);

NAND4xp25_ASAP7_75t_L g9674 ( 
.A(n_9637),
.B(n_4231),
.C(n_4316),
.D(n_4299),
.Y(n_9674)
);

OR2x2_ASAP7_75t_L g9675 ( 
.A(n_9642),
.B(n_9631),
.Y(n_9675)
);

INVx2_ASAP7_75t_L g9676 ( 
.A(n_9640),
.Y(n_9676)
);

AOI21xp5_ASAP7_75t_L g9677 ( 
.A1(n_9641),
.A2(n_9605),
.B(n_9598),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_9661),
.Y(n_9678)
);

OR4x2_ASAP7_75t_L g9679 ( 
.A(n_9643),
.B(n_9604),
.C(n_9639),
.D(n_9602),
.Y(n_9679)
);

NAND4xp25_ASAP7_75t_L g9680 ( 
.A(n_9670),
.B(n_9666),
.C(n_9665),
.D(n_9657),
.Y(n_9680)
);

INVx3_ASAP7_75t_L g9681 ( 
.A(n_9645),
.Y(n_9681)
);

NAND2x1_ASAP7_75t_L g9682 ( 
.A(n_9658),
.B(n_9633),
.Y(n_9682)
);

AND3x2_ASAP7_75t_L g9683 ( 
.A(n_9667),
.B(n_9622),
.C(n_9611),
.Y(n_9683)
);

INVx1_ASAP7_75t_L g9684 ( 
.A(n_9669),
.Y(n_9684)
);

NOR4xp25_ASAP7_75t_L g9685 ( 
.A(n_9655),
.B(n_9647),
.C(n_9668),
.D(n_9651),
.Y(n_9685)
);

NOR2x1_ASAP7_75t_L g9686 ( 
.A(n_9659),
.B(n_9628),
.Y(n_9686)
);

NAND2xp5_ASAP7_75t_L g9687 ( 
.A(n_9649),
.B(n_9634),
.Y(n_9687)
);

INVx1_ASAP7_75t_L g9688 ( 
.A(n_9672),
.Y(n_9688)
);

AND2x4_ASAP7_75t_L g9689 ( 
.A(n_9644),
.B(n_3827),
.Y(n_9689)
);

NOR3xp33_ASAP7_75t_L g9690 ( 
.A(n_9654),
.B(n_3899),
.C(n_3884),
.Y(n_9690)
);

NAND2xp5_ASAP7_75t_L g9691 ( 
.A(n_9664),
.B(n_5020),
.Y(n_9691)
);

NAND4xp75_ASAP7_75t_L g9692 ( 
.A(n_9671),
.B(n_4296),
.C(n_4997),
.D(n_4994),
.Y(n_9692)
);

AND2x2_ASAP7_75t_SL g9693 ( 
.A(n_9652),
.B(n_3797),
.Y(n_9693)
);

INVx1_ASAP7_75t_L g9694 ( 
.A(n_9653),
.Y(n_9694)
);

INVx2_ASAP7_75t_L g9695 ( 
.A(n_9673),
.Y(n_9695)
);

AOI22xp5_ASAP7_75t_L g9696 ( 
.A1(n_9650),
.A2(n_9656),
.B1(n_9674),
.B2(n_9660),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_9663),
.Y(n_9697)
);

OR2x2_ASAP7_75t_L g9698 ( 
.A(n_9648),
.B(n_4053),
.Y(n_9698)
);

NOR2xp67_ASAP7_75t_L g9699 ( 
.A(n_9662),
.B(n_3720),
.Y(n_9699)
);

AND3x4_ASAP7_75t_L g9700 ( 
.A(n_9646),
.B(n_3608),
.C(n_3601),
.Y(n_9700)
);

XOR2xp5_ASAP7_75t_L g9701 ( 
.A(n_9680),
.B(n_3762),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_9676),
.Y(n_9702)
);

INVx2_ASAP7_75t_L g9703 ( 
.A(n_9679),
.Y(n_9703)
);

NAND3xp33_ASAP7_75t_L g9704 ( 
.A(n_9678),
.B(n_9684),
.C(n_9688),
.Y(n_9704)
);

INVx1_ASAP7_75t_L g9705 ( 
.A(n_9681),
.Y(n_9705)
);

XNOR2xp5_ASAP7_75t_L g9706 ( 
.A(n_9683),
.B(n_3762),
.Y(n_9706)
);

INVx1_ASAP7_75t_L g9707 ( 
.A(n_9686),
.Y(n_9707)
);

INVx1_ASAP7_75t_L g9708 ( 
.A(n_9695),
.Y(n_9708)
);

AOI21xp5_ASAP7_75t_L g9709 ( 
.A1(n_9677),
.A2(n_5044),
.B(n_5033),
.Y(n_9709)
);

HB1xp67_ASAP7_75t_L g9710 ( 
.A(n_9697),
.Y(n_9710)
);

NAND2xp5_ASAP7_75t_L g9711 ( 
.A(n_9685),
.B(n_5095),
.Y(n_9711)
);

OAI22xp5_ASAP7_75t_L g9712 ( 
.A1(n_9696),
.A2(n_5095),
.B1(n_4999),
.B2(n_5003),
.Y(n_9712)
);

OA22x2_ASAP7_75t_L g9713 ( 
.A1(n_9694),
.A2(n_4999),
.B1(n_5003),
.B2(n_4998),
.Y(n_9713)
);

XOR2x1_ASAP7_75t_L g9714 ( 
.A(n_9675),
.B(n_4735),
.Y(n_9714)
);

AOI22xp5_ASAP7_75t_L g9715 ( 
.A1(n_9700),
.A2(n_3818),
.B1(n_3826),
.B2(n_3803),
.Y(n_9715)
);

INVx2_ASAP7_75t_L g9716 ( 
.A(n_9682),
.Y(n_9716)
);

XNOR2xp5_ASAP7_75t_L g9717 ( 
.A(n_9687),
.B(n_3762),
.Y(n_9717)
);

AOI222xp33_ASAP7_75t_L g9718 ( 
.A1(n_9699),
.A2(n_5041),
.B1(n_5037),
.B2(n_5042),
.C1(n_5039),
.C2(n_5032),
.Y(n_9718)
);

OAI22xp5_ASAP7_75t_L g9719 ( 
.A1(n_9693),
.A2(n_5039),
.B1(n_5041),
.B2(n_5037),
.Y(n_9719)
);

XOR2xp5_ASAP7_75t_L g9720 ( 
.A(n_9689),
.B(n_3762),
.Y(n_9720)
);

BUFx6f_ASAP7_75t_L g9721 ( 
.A(n_9691),
.Y(n_9721)
);

NAND5xp2_ASAP7_75t_L g9722 ( 
.A(n_9690),
.B(n_4853),
.C(n_4806),
.D(n_4781),
.E(n_4310),
.Y(n_9722)
);

OAI22x1_ASAP7_75t_SL g9723 ( 
.A1(n_9692),
.A2(n_3653),
.B1(n_3656),
.B2(n_3634),
.Y(n_9723)
);

INVx2_ASAP7_75t_L g9724 ( 
.A(n_9703),
.Y(n_9724)
);

INVx1_ASAP7_75t_L g9725 ( 
.A(n_9710),
.Y(n_9725)
);

OAI22xp5_ASAP7_75t_L g9726 ( 
.A1(n_9704),
.A2(n_9698),
.B1(n_3909),
.B2(n_3832),
.Y(n_9726)
);

AOI22x1_ASAP7_75t_L g9727 ( 
.A1(n_9702),
.A2(n_3818),
.B1(n_3826),
.B2(n_3803),
.Y(n_9727)
);

AOI22xp5_ASAP7_75t_L g9728 ( 
.A1(n_9707),
.A2(n_5044),
.B1(n_5033),
.B2(n_3826),
.Y(n_9728)
);

OAI22xp5_ASAP7_75t_L g9729 ( 
.A1(n_9705),
.A2(n_3909),
.B1(n_5088),
.B2(n_5065),
.Y(n_9729)
);

OAI22xp5_ASAP7_75t_L g9730 ( 
.A1(n_9716),
.A2(n_5017),
.B1(n_5019),
.B2(n_5016),
.Y(n_9730)
);

INVx1_ASAP7_75t_L g9731 ( 
.A(n_9708),
.Y(n_9731)
);

AO22x2_ASAP7_75t_L g9732 ( 
.A1(n_9701),
.A2(n_4330),
.B1(n_5015),
.B2(n_5006),
.Y(n_9732)
);

AND2x2_ASAP7_75t_L g9733 ( 
.A(n_9721),
.B(n_5023),
.Y(n_9733)
);

INVx2_ASAP7_75t_L g9734 ( 
.A(n_9721),
.Y(n_9734)
);

XNOR2xp5_ASAP7_75t_L g9735 ( 
.A(n_9706),
.B(n_4806),
.Y(n_9735)
);

INVx1_ASAP7_75t_SL g9736 ( 
.A(n_9711),
.Y(n_9736)
);

OA22x2_ASAP7_75t_L g9737 ( 
.A1(n_9717),
.A2(n_5015),
.B1(n_5016),
.B2(n_5006),
.Y(n_9737)
);

INVx2_ASAP7_75t_L g9738 ( 
.A(n_9720),
.Y(n_9738)
);

XOR2xp5_ASAP7_75t_L g9739 ( 
.A(n_9709),
.B(n_3797),
.Y(n_9739)
);

AOI22x1_ASAP7_75t_L g9740 ( 
.A1(n_9718),
.A2(n_3828),
.B1(n_3849),
.B2(n_3818),
.Y(n_9740)
);

XOR2xp5_ASAP7_75t_L g9741 ( 
.A(n_9723),
.B(n_3797),
.Y(n_9741)
);

INVx1_ASAP7_75t_L g9742 ( 
.A(n_9713),
.Y(n_9742)
);

INVx1_ASAP7_75t_L g9743 ( 
.A(n_9714),
.Y(n_9743)
);

CKINVDCx20_ASAP7_75t_R g9744 ( 
.A(n_9725),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_9724),
.Y(n_9745)
);

NAND2xp5_ASAP7_75t_L g9746 ( 
.A(n_9731),
.B(n_9715),
.Y(n_9746)
);

AOI22xp5_ASAP7_75t_L g9747 ( 
.A1(n_9734),
.A2(n_9719),
.B1(n_9712),
.B2(n_9722),
.Y(n_9747)
);

INVx2_ASAP7_75t_L g9748 ( 
.A(n_9743),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_9736),
.Y(n_9749)
);

BUFx2_ASAP7_75t_L g9750 ( 
.A(n_9738),
.Y(n_9750)
);

CKINVDCx20_ASAP7_75t_R g9751 ( 
.A(n_9742),
.Y(n_9751)
);

CKINVDCx20_ASAP7_75t_R g9752 ( 
.A(n_9726),
.Y(n_9752)
);

AND2x2_ASAP7_75t_L g9753 ( 
.A(n_9733),
.B(n_4814),
.Y(n_9753)
);

AOI22xp33_ASAP7_75t_L g9754 ( 
.A1(n_9741),
.A2(n_5044),
.B1(n_4045),
.B2(n_4125),
.Y(n_9754)
);

HB1xp67_ASAP7_75t_L g9755 ( 
.A(n_9735),
.Y(n_9755)
);

OAI22xp5_ASAP7_75t_SL g9756 ( 
.A1(n_9739),
.A2(n_3738),
.B1(n_3746),
.B2(n_3720),
.Y(n_9756)
);

OAI21xp5_ASAP7_75t_L g9757 ( 
.A1(n_9740),
.A2(n_4408),
.B(n_4497),
.Y(n_9757)
);

INVxp67_ASAP7_75t_SL g9758 ( 
.A(n_9745),
.Y(n_9758)
);

INVx2_ASAP7_75t_L g9759 ( 
.A(n_9751),
.Y(n_9759)
);

INVx1_ASAP7_75t_L g9760 ( 
.A(n_9744),
.Y(n_9760)
);

INVx1_ASAP7_75t_L g9761 ( 
.A(n_9750),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_9749),
.Y(n_9762)
);

INVx1_ASAP7_75t_L g9763 ( 
.A(n_9748),
.Y(n_9763)
);

HB1xp67_ASAP7_75t_L g9764 ( 
.A(n_9755),
.Y(n_9764)
);

INVx1_ASAP7_75t_L g9765 ( 
.A(n_9746),
.Y(n_9765)
);

INVxp67_ASAP7_75t_SL g9766 ( 
.A(n_9752),
.Y(n_9766)
);

INVx1_ASAP7_75t_L g9767 ( 
.A(n_9747),
.Y(n_9767)
);

INVx2_ASAP7_75t_L g9768 ( 
.A(n_9753),
.Y(n_9768)
);

INVx1_ASAP7_75t_L g9769 ( 
.A(n_9756),
.Y(n_9769)
);

AOI22xp5_ASAP7_75t_L g9770 ( 
.A1(n_9761),
.A2(n_9728),
.B1(n_9754),
.B2(n_9737),
.Y(n_9770)
);

AOI22xp33_ASAP7_75t_L g9771 ( 
.A1(n_9759),
.A2(n_9727),
.B1(n_9732),
.B2(n_9757),
.Y(n_9771)
);

INVxp67_ASAP7_75t_SL g9772 ( 
.A(n_9764),
.Y(n_9772)
);

INVx2_ASAP7_75t_L g9773 ( 
.A(n_9760),
.Y(n_9773)
);

INVx1_ASAP7_75t_L g9774 ( 
.A(n_9766),
.Y(n_9774)
);

INVx1_ASAP7_75t_L g9775 ( 
.A(n_9772),
.Y(n_9775)
);

AOI21xp33_ASAP7_75t_L g9776 ( 
.A1(n_9774),
.A2(n_9758),
.B(n_9763),
.Y(n_9776)
);

INVx2_ASAP7_75t_L g9777 ( 
.A(n_9773),
.Y(n_9777)
);

INVx1_ASAP7_75t_L g9778 ( 
.A(n_9770),
.Y(n_9778)
);

INVx1_ASAP7_75t_L g9779 ( 
.A(n_9775),
.Y(n_9779)
);

CKINVDCx16_ASAP7_75t_R g9780 ( 
.A(n_9777),
.Y(n_9780)
);

NAND2xp5_ASAP7_75t_L g9781 ( 
.A(n_9780),
.B(n_9762),
.Y(n_9781)
);

OAI21x1_ASAP7_75t_L g9782 ( 
.A1(n_9781),
.A2(n_9765),
.B(n_9779),
.Y(n_9782)
);

AOI21xp5_ASAP7_75t_L g9783 ( 
.A1(n_9782),
.A2(n_9776),
.B(n_9778),
.Y(n_9783)
);

OAI21xp5_ASAP7_75t_L g9784 ( 
.A1(n_9783),
.A2(n_9767),
.B(n_9768),
.Y(n_9784)
);

AOI22xp5_ASAP7_75t_L g9785 ( 
.A1(n_9783),
.A2(n_9769),
.B1(n_9771),
.B2(n_9732),
.Y(n_9785)
);

AOI22xp33_ASAP7_75t_L g9786 ( 
.A1(n_9784),
.A2(n_9729),
.B1(n_9730),
.B2(n_5044),
.Y(n_9786)
);

AOI21xp33_ASAP7_75t_SL g9787 ( 
.A1(n_9786),
.A2(n_9785),
.B(n_3906),
.Y(n_9787)
);

AOI211xp5_ASAP7_75t_L g9788 ( 
.A1(n_9787),
.A2(n_3906),
.B(n_3797),
.C(n_3672),
.Y(n_9788)
);


endmodule