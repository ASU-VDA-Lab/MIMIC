module real_jpeg_9815_n_17 (n_5, n_4, n_8, n_0, n_12, n_299, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_299;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_211;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_295;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_1),
.A2(n_49),
.B(n_59),
.C(n_127),
.D(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_49),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_1),
.B(n_47),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_1),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_83),
.B(n_146),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_1),
.A2(n_32),
.B(n_43),
.C(n_180),
.D(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_1),
.B(n_115),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_1),
.A2(n_29),
.B(n_33),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_27),
.B1(n_35),
.B2(n_161),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_55),
.B1(n_64),
.B2(n_66),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_4),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_64),
.B1(n_66),
.B2(n_92),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_5),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_164),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_154),
.B1(n_190),
.B2(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_64),
.B1(n_66),
.B2(n_141),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_141),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_141),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_11),
.A2(n_38),
.B1(n_64),
.B2(n_66),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_52),
.B1(n_64),
.B2(n_66),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_14),
.A2(n_27),
.B1(n_35),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_64),
.B1(n_66),
.B2(n_113),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_113),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_113),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_16),
.A2(n_36),
.B1(n_64),
.B2(n_66),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_16),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_26),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_26),
.A2(n_31),
.B1(n_112),
.B2(n_245),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_27),
.A2(n_28),
.B(n_161),
.C(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_34),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_31),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_31),
.A2(n_90),
.B(n_245),
.Y(n_244)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_44),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_70),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_42),
.A2(n_53),
.B1(n_199),
.B2(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_42),
.A2(n_233),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_47),
.B1(n_51),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_43),
.A2(n_47),
.B1(n_74),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_43),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_48),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_49),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_53),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_53),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_53),
.A2(n_200),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_68),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_67),
.B1(n_77),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_67),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_58),
.A2(n_67),
.B1(n_140),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_58),
.A2(n_178),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_58),
.A2(n_67),
.B1(n_107),
.B2(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_63),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_59),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_60),
.B(n_66),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_64),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_84),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_66),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_67),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_67),
.A2(n_142),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_81),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_88),
.B1(n_89),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_280),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_83),
.A2(n_84),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_83),
.A2(n_84),
.B1(n_105),
.B2(n_223),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_84),
.A2(n_153),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_161),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_93),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_95),
.Y(n_285)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_101),
.A2(n_102),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_110),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_103),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_104),
.B(n_106),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_108),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_114),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_273),
.A3(n_286),
.B1(n_292),
.B2(n_297),
.C(n_299),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_239),
.C(n_269),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_212),
.B(n_238),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_193),
.B(n_211),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_172),
.B(n_192),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_149),
.B(n_171),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_139),
.C(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_158),
.B(n_170),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_165),
.B(n_169),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_174),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_191),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_184),
.C(n_191),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_207),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_208),
.C(n_209),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_206),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_214),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_227),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_226),
.C(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_221),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_240),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_255),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_255),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_251),
.C(n_254),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_267),
.B2(n_268),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_259),
.C(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_262),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_274),
.B(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.C(n_281),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);


endmodule