module real_jpeg_12605_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_45),
.B1(n_49),
.B2(n_66),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_45),
.B1(n_49),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_7),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_37),
.B1(n_45),
.B2(n_49),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_26),
.B(n_32),
.C(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_13),
.B(n_27),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_27),
.B(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_13),
.B(n_60),
.C(n_77),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_72),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_59),
.B1(n_63),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_13),
.B(n_55),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_14),
.A2(n_42),
.B1(n_60),
.B2(n_61),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_45),
.B1(n_49),
.B2(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_15),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_27),
.A2(n_30),
.B(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_SL g141 ( 
.A(n_28),
.B(n_47),
.C(n_49),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_36),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_43),
.A2(n_44),
.B1(n_101),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_43),
.A2(n_44),
.B1(n_120),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_49),
.B1(n_77),
.B2(n_78),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_45),
.A2(n_48),
.B(n_139),
.C(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_45),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_69),
.B1(n_70),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_89),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_58),
.A2(n_64),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_59),
.A2(n_63),
.B1(n_170),
.B2(n_178),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_59),
.A2(n_172),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_63),
.B(n_72),
.Y(n_176)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_65),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_64),
.B(n_144),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_72),
.B(n_76),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_91),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_86),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B(n_81),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_98),
.B1(n_134),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_84),
.A2(n_98),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_84),
.A2(n_98),
.B1(n_157),
.B2(n_167),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_102),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_97),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_94),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_113),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_202),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_145),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_129),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_136),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_158),
.B(n_201),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_195),
.B(n_200),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_184),
.B(n_194),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_173),
.B(n_183),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_168),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_165),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_179),
.B(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.C(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_199),
.Y(n_200)
);


endmodule