module real_jpeg_26101_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_355, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_355;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_37),
.B1(n_71),
.B2(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_1),
.A2(n_37),
.B1(n_220),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_61),
.B1(n_71),
.B2(n_72),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_3),
.A2(n_71),
.B1(n_72),
.B2(n_117),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_3),
.A2(n_48),
.B1(n_62),
.B2(n_117),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_71),
.B1(n_72),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_134),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_134),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_4),
.A2(n_47),
.B1(n_58),
.B2(n_134),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_6),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_6),
.A2(n_71),
.B1(n_72),
.B2(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_6),
.A2(n_82),
.B1(n_126),
.B2(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx8_ASAP7_75t_SL g56 ( 
.A(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_42),
.B1(n_58),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_42),
.B1(n_71),
.B2(n_72),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_10),
.A2(n_50),
.B1(n_71),
.B2(n_72),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_50),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_11),
.A2(n_67),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_11),
.B(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_129),
.B1(n_153),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_33),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_11),
.B(n_59),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_15),
.Y(n_132)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_15),
.Y(n_146)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_101),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_99),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_19),
.B(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_76),
.B2(n_87),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_63),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_22),
.A2(n_23),
.B1(n_63),
.B2(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_25),
.A2(n_39),
.B(n_234),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_26),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_26),
.A2(n_38),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_27),
.A2(n_29),
.A3(n_33),
.B1(n_169),
.B2(n_178),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_28),
.A2(n_29),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_28),
.B(n_31),
.Y(n_178)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_29),
.A2(n_69),
.B(n_113),
.C(n_119),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_32),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_32),
.A2(n_98),
.B(n_170),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_33),
.B(n_55),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_34),
.B(n_113),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_34),
.A2(n_48),
.A3(n_54),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_39),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_39),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_39),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_39),
.A2(n_85),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_39),
.A2(n_85),
.B1(n_196),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_39),
.A2(n_85),
.B1(n_96),
.B2(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_85),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_43),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_53),
.B(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_47),
.A2(n_113),
.B(n_219),
.Y(n_239)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_48),
.Y(n_220)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_60),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_81),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_51),
.A2(n_59),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_51),
.A2(n_59),
.B1(n_240),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_52),
.A2(n_53),
.B1(n_252),
.B2(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_52),
.A2(n_270),
.B(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_52),
.A2(n_80),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_59),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_63),
.A2(n_64),
.B1(n_95),
.B2(n_340),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_92),
.C(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_74),
.B(n_75),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_65),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_65),
.A2(n_74),
.B1(n_116),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_65),
.A2(n_74),
.B1(n_125),
.B2(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_65),
.A2(n_75),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_65),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_70),
.B(n_113),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_70),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_70),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_70),
.A2(n_114),
.B1(n_259),
.B2(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_71),
.B(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_74),
.B(n_75),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_94),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_338),
.Y(n_345)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_92),
.A2(n_338),
.B1(n_339),
.B2(n_341),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_92),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_94),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_95),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_335),
.A3(n_346),
.B1(n_351),
.B2(n_352),
.C(n_355),
.Y(n_101)
);

AOI311xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_286),
.A3(n_325),
.B(n_329),
.C(n_330),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_242),
.C(n_281),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_213),
.B(n_241),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_189),
.B(n_212),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_162),
.B(n_188),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_139),
.B(n_161),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_120),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_156),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_113),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_114),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_114),
.A2(n_276),
.B(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B(n_135),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_138),
.B1(n_143),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_129),
.A2(n_181),
.B(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_129),
.A2(n_156),
.B(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_130),
.B(n_185),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_130),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_222)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_135),
.B(n_203),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_149),
.B(n_160),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_147),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_154),
.B(n_159),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_176),
.B1(n_186),
.B2(n_187),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_175),
.C(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_179),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_204),
.B2(n_205),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_207),
.C(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_199),
.C(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_209),
.B(n_260),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_215),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_231),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_230),
.C(n_231),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_226),
.Y(n_247)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_222),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_235),
.C(n_238),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_243),
.A2(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_262),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_244),
.B(n_262),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.C(n_255),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_246),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_249),
.C(n_250),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_254),
.B(n_255),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_277),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_264),
.B(n_277),
.C(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_272),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_287),
.A2(n_326),
.B(n_331),
.C(n_334),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_307),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_307),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_300),
.C(n_306),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_289),
.B(n_300),
.CI(n_306),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_299),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_293),
.C(n_297),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_295),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_303),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_305),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_315),
.B(n_319),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_324),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_337),
.B1(n_342),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_322),
.C(n_324),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_344),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_336),
.B(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.C(n_343),
.Y(n_336)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_347),
.B(n_348),
.Y(n_351)
);


endmodule