module fake_jpeg_18695_n_184 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_15),
.B1(n_12),
.B2(n_16),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_26),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_22),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_45),
.B(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_22),
.B(n_30),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_41),
.B1(n_34),
.B2(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_34),
.B1(n_38),
.B2(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_27),
.B1(n_49),
.B2(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_44),
.B1(n_64),
.B2(n_18),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_40),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_77),
.B(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_45),
.B1(n_49),
.B2(n_32),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_59),
.B1(n_61),
.B2(n_56),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_16),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_67),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_96),
.B1(n_44),
.B2(n_14),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_95),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_79),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_65),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_54),
.B(n_57),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_77),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_27),
.C(n_35),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_77),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_14),
.B1(n_11),
.B2(n_16),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_108),
.B1(n_112),
.B2(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_11),
.B1(n_14),
.B2(n_16),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_92),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_125),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_104),
.C(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_129),
.C(n_103),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_95),
.C(n_84),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_111),
.C(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_130),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_96),
.C(n_91),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_91),
.C(n_64),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_12),
.C(n_23),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_102),
.B1(n_97),
.B2(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_140),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_143),
.C(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_112),
.B1(n_110),
.B2(n_106),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_8),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_5),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_135),
.C(n_143),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_123),
.B(n_118),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_148),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_116),
.C(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_124),
.B(n_16),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_21),
.B(n_13),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_16),
.C(n_13),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_13),
.C(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_6),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_4),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_157),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_132),
.B(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_21),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_0),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_163),
.B(n_167),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_165),
.B(n_4),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_13),
.B1(n_21),
.B2(n_2),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_168),
.B(n_0),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_155),
.C(n_13),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_170),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_13),
.B(n_9),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_21),
.C(n_3),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_3),
.C(n_4),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_1),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_1),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_1),
.C(n_2),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_177),
.B(n_1),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);


endmodule