module fake_jpeg_3246_n_64 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_64);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_19),
.Y(n_29)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_21),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_22),
.Y(n_38)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_27),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_25),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_20),
.C(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_48),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_2),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_39),
.B2(n_3),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_55),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

AOI321xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_52),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C(n_6),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_56),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_58),
.B(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_7),
.Y(n_64)
);


endmodule