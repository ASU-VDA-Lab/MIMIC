module fake_jpeg_1583_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_9),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_27),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_20),
.B(n_33),
.C(n_38),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_19),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g93 ( 
.A(n_48),
.B(n_6),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_42),
.B1(n_35),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_2),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_87),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_33),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_18),
.B1(n_38),
.B2(n_40),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_78),
.B1(n_68),
.B2(n_50),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_80)
);

OAI21x1_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_18),
.B1(n_32),
.B2(n_16),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_76),
.B1(n_74),
.B2(n_93),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_59),
.B1(n_7),
.B2(n_13),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_2),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_10),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_50),
.B1(n_68),
.B2(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_103),
.B1(n_108),
.B2(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_58),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_58),
.C(n_52),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_72),
.C(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_59),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_132),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_81),
.B1(n_131),
.B2(n_128),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_74),
.B(n_113),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_97),
.C(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_74),
.B1(n_72),
.B2(n_75),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_113),
.B1(n_117),
.B2(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_73),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_112),
.Y(n_142)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_97),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.C(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_149),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_130),
.B(n_119),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_112),
.C(n_100),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_124),
.C(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_75),
.B1(n_98),
.B2(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_120),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_123),
.B(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_153),
.A2(n_136),
.B1(n_148),
.B2(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_167),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_134),
.B1(n_146),
.B2(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_142),
.B1(n_145),
.B2(n_118),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_150),
.C(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_150),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_174),
.B1(n_159),
.B2(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_157),
.Y(n_174)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_152),
.B1(n_168),
.B2(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_169),
.C(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_174),
.C(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_177),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_175),
.B(n_81),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_81),
.Y(n_188)
);


endmodule