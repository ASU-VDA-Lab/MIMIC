module fake_netlist_5_2419_n_2005 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2005);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2005;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_28),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_4),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_112),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_104),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_60),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_28),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_54),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_27),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_54),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_128),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_93),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_108),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_122),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_63),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_132),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_77),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_36),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_48),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_115),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_64),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_152),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_47),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_56),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_177),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_78),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_185),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_163),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_9),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_10),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_63),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_19),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_56),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_90),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_69),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_12),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_186),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_191),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_193),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_116),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_120),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_196),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_159),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_158),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_165),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_117),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_73),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_118),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_89),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_102),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_27),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_150),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_111),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_67),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_153),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_110),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_130),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_178),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_84),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_26),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_92),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_164),
.Y(n_309)
);

BUFx8_ASAP7_75t_SL g310 ( 
.A(n_85),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_81),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_144),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_124),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_169),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_30),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_1),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_45),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_95),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_12),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_98),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_141),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_137),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_97),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_145),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_121),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_136),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_174),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_8),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_29),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_26),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_107),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_103),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_15),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_25),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_74),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_53),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_66),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_171),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_16),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_43),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_140),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_64),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_59),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_42),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_25),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_13),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_187),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_147),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_99),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_192),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_183),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_46),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_24),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_49),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_94),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_79),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_20),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_65),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_105),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_135),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_5),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_129),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_60),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_131),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_55),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_39),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_119),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_134),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_51),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_100),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_167),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_86),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_65),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_38),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_109),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_19),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_11),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_18),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_170),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_133),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_197),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_38),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_62),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_46),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_13),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_55),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_76),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_160),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_24),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_57),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_30),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_285),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_285),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_378),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_263),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_391),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_391),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_201),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_204),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_202),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_207),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_204),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_275),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_284),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_216),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_271),
.B(n_194),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_R g415 ( 
.A(n_206),
.B(n_2),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_271),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_206),
.B(n_312),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_287),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_219),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_313),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_285),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_312),
.B(n_2),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_285),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_216),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_223),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_285),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_220),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_231),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_310),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_229),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_242),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_229),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_246),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_200),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_306),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_3),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_233),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_233),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_249),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_364),
.B(n_3),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_203),
.B(n_5),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_255),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_256),
.Y(n_446)
);

BUFx6f_ASAP7_75t_SL g447 ( 
.A(n_228),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_257),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_257),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_258),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_306),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_268),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_341),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_259),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_264),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_274),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_278),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_285),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_280),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_293),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_293),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_341),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_295),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_384),
.B(n_6),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_199),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_205),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_295),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_208),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_298),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_200),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_298),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_234),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_209),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_214),
.B(n_6),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_299),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_212),
.B(n_10),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_214),
.B(n_11),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_299),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_210),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_314),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_212),
.B(n_16),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_314),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_321),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_211),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_213),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_321),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_234),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_329),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_221),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_329),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_296),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_234),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_291),
.B(n_17),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_215),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_217),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_301),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_307),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_416),
.B(n_230),
.Y(n_500)
);

INVx6_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_481),
.A2(n_241),
.B(n_210),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_422),
.B(n_243),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_474),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_459),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_400),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_R g521 ( 
.A(n_401),
.B(n_316),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_414),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_414),
.B(n_271),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_230),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_273),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_438),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_417),
.B(n_228),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_398),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_273),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_244),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_430),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_431),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_441),
.B(n_244),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_449),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_226),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_461),
.B(n_273),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_464),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_469),
.B(n_227),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_232),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_477),
.A2(n_482),
.B(n_480),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_485),
.B(n_286),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_488),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_490),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_492),
.B(n_286),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_452),
.A2(n_238),
.B1(n_237),
.B2(n_239),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_408),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_437),
.B(n_286),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_495),
.B(n_354),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_403),
.B(n_354),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_465),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_571),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_534),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_512),
.B(n_404),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_467),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_408),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_505),
.B(n_409),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

HB1xp67_ASAP7_75t_SL g587 ( 
.A(n_542),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_519),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_519),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_456),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_570),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_572),
.B(n_409),
.Y(n_593)
);

BUFx8_ASAP7_75t_SL g594 ( 
.A(n_538),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_291),
.B1(n_315),
.B2(n_283),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_570),
.B(n_419),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_571),
.B(n_466),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_419),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_523),
.B(n_570),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_523),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_516),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_570),
.B(n_425),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_523),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_532),
.B(n_425),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_570),
.B(n_429),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_523),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_527),
.Y(n_611)
);

INVx4_ASAP7_75t_SL g612 ( 
.A(n_501),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_527),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_523),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_523),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_562),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_572),
.B(n_429),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_516),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_533),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_533),
.Y(n_622)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_501),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_572),
.B(n_433),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

CKINVDCx6p67_ASAP7_75t_R g627 ( 
.A(n_567),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_535),
.B(n_531),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_544),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_538),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_548),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_531),
.B(n_468),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_541),
.B(n_433),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_544),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_562),
.B(n_402),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_549),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_534),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_520),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_541),
.B(n_415),
.C(n_241),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_579),
.B(n_470),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_517),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_579),
.B(n_241),
.C(n_210),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_503),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_574),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_503),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_570),
.B(n_435),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_530),
.B(n_300),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_574),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_517),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_503),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_517),
.Y(n_657)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_500),
.A2(n_340),
.B(n_335),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_576),
.B(n_475),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_570),
.B(n_354),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_517),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_507),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_507),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_507),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_503),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_576),
.B(n_486),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_532),
.B(n_435),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_507),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_520),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_572),
.B(n_446),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_574),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_574),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_570),
.B(n_446),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_540),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_578),
.B(n_450),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_502),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_530),
.B(n_450),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_503),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_515),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_574),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_515),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_576),
.A2(n_315),
.B1(n_283),
.B2(n_394),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_520),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_530),
.B(n_335),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_530),
.B(n_455),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_548),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_578),
.B(n_455),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_530),
.B(n_457),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_501),
.A2(n_355),
.B1(n_361),
.B2(n_340),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_501),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_530),
.B(n_300),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_574),
.B(n_457),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_503),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_402),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_578),
.B(n_458),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_550),
.B(n_458),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_500),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_577),
.A2(n_374),
.B1(n_266),
.B2(n_243),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_506),
.Y(n_708)
);

BUFx4f_ASAP7_75t_L g709 ( 
.A(n_558),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_577),
.A2(n_283),
.B1(n_356),
.B2(n_330),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_506),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_557),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_506),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_540),
.B(n_569),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_557),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_511),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_569),
.B(n_405),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_561),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_561),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_550),
.B(n_460),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_577),
.A2(n_487),
.B1(n_497),
.B2(n_496),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_300),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_552),
.B(n_355),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_561),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_558),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_575),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_578),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_558),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_540),
.B(n_460),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_511),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_573),
.B(n_493),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_628),
.B(n_555),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_555),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_603),
.B(n_556),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_588),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_706),
.B(n_556),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_580),
.B(n_596),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_721),
.B(n_566),
.C(n_405),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_603),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_613),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_588),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_637),
.B(n_611),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_643),
.A2(n_221),
.B(n_224),
.C(n_222),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_580),
.B(n_573),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_615),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_705),
.B(n_493),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_599),
.B(n_573),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_603),
.A2(n_412),
.B1(n_418),
.B2(n_411),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_714),
.B(n_552),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_611),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_606),
.B(n_609),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_727),
.B(n_590),
.Y(n_752)
);

OAI21xp33_ASAP7_75t_L g753 ( 
.A1(n_634),
.A2(n_568),
.B(n_575),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_662),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_652),
.B(n_548),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_589),
.Y(n_756)
);

BUFx6f_ASAP7_75t_SL g757 ( 
.A(n_617),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_725),
.B(n_320),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_649),
.A2(n_525),
.B(n_524),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_725),
.A2(n_222),
.B1(n_225),
.B2(n_224),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_662),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_676),
.B(n_525),
.Y(n_762)
);

NOR3xp33_ASAP7_75t_L g763 ( 
.A(n_583),
.B(n_667),
.C(n_659),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_615),
.B(n_235),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_727),
.B(n_568),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_663),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_615),
.B(n_536),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_615),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_720),
.B(n_498),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_635),
.A2(n_521),
.B1(n_454),
.B2(n_463),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_617),
.Y(n_771)
);

NOR2x1p5_ASAP7_75t_L g772 ( 
.A(n_627),
.B(n_567),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_683),
.A2(n_420),
.B1(n_327),
.B2(n_320),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_615),
.B(n_536),
.Y(n_774)
);

NOR2x1p5_ASAP7_75t_L g775 ( 
.A(n_627),
.B(n_567),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_691),
.A2(n_521),
.B1(n_552),
.B2(n_560),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_637),
.B(n_498),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_589),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_663),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_695),
.A2(n_560),
.B1(n_552),
.B2(n_499),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_664),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_728),
.A2(n_289),
.B1(n_383),
.B2(n_247),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_643),
.A2(n_350),
.B(n_395),
.C(n_383),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_714),
.B(n_558),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_633),
.B(n_552),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_646),
.A2(n_374),
.B1(n_266),
.B2(n_568),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_728),
.B(n_320),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_590),
.B(n_575),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_702),
.B(n_499),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_R g790 ( 
.A(n_632),
.B(n_587),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_700),
.A2(n_552),
.B1(n_560),
.B2(n_373),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_649),
.B(n_558),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_633),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_654),
.B(n_558),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_598),
.B(n_536),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_697),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_709),
.A2(n_327),
.B1(n_393),
.B2(n_375),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_702),
.B(n_565),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_664),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_633),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_654),
.B(n_560),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_600),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_669),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_672),
.B(n_560),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_642),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_598),
.B(n_536),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_618),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_669),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_598),
.B(n_536),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_560),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_598),
.B(n_536),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_673),
.B(n_686),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_645),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_597),
.B(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_592),
.B(n_536),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_592),
.B(n_536),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_673),
.B(n_536),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_SL g818 ( 
.A(n_581),
.B(n_566),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_645),
.Y(n_819)
);

INVxp33_ASAP7_75t_L g820 ( 
.A(n_644),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_686),
.B(n_522),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_584),
.B(n_436),
.C(n_432),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_597),
.B(n_564),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_717),
.B(n_447),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_618),
.B(n_522),
.Y(n_826)
);

AND2x4_ASAP7_75t_SL g827 ( 
.A(n_722),
.B(n_228),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_621),
.B(n_522),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_645),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_717),
.B(n_447),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_621),
.B(n_522),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_655),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_709),
.A2(n_366),
.B1(n_289),
.B2(n_382),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_655),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_622),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_622),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_731),
.B(n_447),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_592),
.B(n_524),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_731),
.B(n_677),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_608),
.B(n_729),
.C(n_668),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_722),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_709),
.A2(n_366),
.B1(n_382),
.B2(n_317),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_647),
.A2(n_317),
.B1(n_225),
.B2(n_395),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_585),
.A2(n_376),
.B1(n_564),
.B2(n_253),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_641),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_592),
.B(n_524),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_591),
.B(n_564),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_655),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_629),
.B(n_524),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_608),
.B(n_547),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_629),
.B(n_526),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_601),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_668),
.B(n_218),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_600),
.B(n_526),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_526),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_604),
.A2(n_504),
.B(n_526),
.Y(n_856)
);

AND2x6_ASAP7_75t_SL g857 ( 
.A(n_722),
.B(n_247),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_631),
.B(n_528),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_586),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_586),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_600),
.B(n_604),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_604),
.B(n_327),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_636),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_641),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_729),
.B(n_619),
.C(n_593),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_636),
.B(n_528),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_639),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_601),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_640),
.B(n_292),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_639),
.B(n_528),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_650),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_605),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_722),
.B(n_315),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_650),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_604),
.A2(n_504),
.B(n_547),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_605),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_675),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_653),
.B(n_236),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_602),
.B(n_303),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_625),
.B(n_671),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_690),
.A2(n_311),
.B1(n_392),
.B2(n_386),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_675),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_678),
.B(n_528),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_678),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_620),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_694),
.B(n_698),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_694),
.B(n_529),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_620),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_698),
.B(n_529),
.Y(n_889)
);

BUFx6f_ASAP7_75t_SL g890 ( 
.A(n_722),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_602),
.B(n_262),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_704),
.B(n_529),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_582),
.Y(n_893)
);

AND2x4_ASAP7_75t_SL g894 ( 
.A(n_690),
.B(n_723),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_607),
.B(n_610),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_679),
.B(n_322),
.Y(n_896)
);

BUFx6f_ASAP7_75t_SL g897 ( 
.A(n_594),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_642),
.Y(n_898)
);

AO221x1_ASAP7_75t_L g899 ( 
.A1(n_707),
.A2(n_357),
.B1(n_260),
.B2(n_261),
.C(n_269),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_693),
.B(n_331),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_SL g901 ( 
.A(n_623),
.B(n_624),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_732),
.B(n_736),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_833),
.A2(n_610),
.B1(n_614),
.B2(n_607),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_790),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_763),
.A2(n_690),
.B1(n_699),
.B2(n_653),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_735),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_737),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_741),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_733),
.B(n_704),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_850),
.B(n_712),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_756),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_751),
.A2(n_630),
.B(n_624),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_739),
.B(n_653),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_747),
.B(n_712),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_812),
.A2(n_630),
.B(n_624),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_755),
.A2(n_630),
.B(n_624),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_788),
.B(n_715),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_743),
.A2(n_696),
.B(n_703),
.C(n_715),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_801),
.A2(n_665),
.B(n_630),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_805),
.Y(n_920)
);

OAI22x1_ASAP7_75t_L g921 ( 
.A1(n_770),
.A2(n_670),
.B1(n_689),
.B2(n_582),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_804),
.A2(n_665),
.B(n_610),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_758),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_810),
.A2(n_665),
.B(n_610),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_739),
.B(n_665),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_833),
.A2(n_647),
.B1(n_658),
.B2(n_653),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_762),
.A2(n_614),
.B(n_607),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_823),
.B(n_718),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_746),
.B(n_718),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_792),
.A2(n_614),
.B(n_607),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_794),
.A2(n_616),
.B(n_614),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_746),
.B(n_719),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_739),
.B(n_616),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_752),
.B(n_814),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_842),
.A2(n_595),
.B(n_724),
.C(n_719),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_815),
.A2(n_616),
.B(n_623),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_815),
.A2(n_616),
.B(n_623),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_820),
.B(n_724),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_769),
.B(n_690),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_778),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_769),
.B(n_641),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_869),
.B(n_387),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_842),
.A2(n_688),
.B(n_710),
.C(n_723),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_760),
.A2(n_658),
.B1(n_699),
.B2(n_653),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_816),
.A2(n_623),
.B(n_660),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_816),
.A2(n_623),
.B(n_660),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_880),
.A2(n_653),
.B1(n_699),
.B2(n_723),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_734),
.A2(n_660),
.B(n_680),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_744),
.B(n_692),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_807),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_784),
.A2(n_699),
.B(n_653),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_820),
.B(n_692),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_835),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_734),
.A2(n_660),
.B(n_680),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_839),
.B(n_692),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_836),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_841),
.B(n_660),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_863),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_840),
.A2(n_697),
.B1(n_623),
.B2(n_723),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_SL g960 ( 
.A1(n_797),
.A2(n_375),
.B(n_361),
.C(n_393),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_682),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_760),
.A2(n_658),
.B1(n_699),
.B2(n_696),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_867),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_765),
.B(n_753),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_875),
.A2(n_699),
.B(n_708),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_871),
.B(n_874),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_877),
.B(n_682),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_802),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_745),
.A2(n_730),
.B(n_716),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_882),
.B(n_884),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_749),
.B(n_685),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_768),
.A2(n_730),
.B(n_716),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_817),
.A2(n_730),
.B(n_716),
.Y(n_973)
);

BUFx8_ASAP7_75t_L g974 ( 
.A(n_897),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_856),
.A2(n_699),
.B(n_708),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_838),
.A2(n_730),
.B(n_716),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_739),
.B(n_612),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_749),
.B(n_685),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_782),
.A2(n_350),
.B(n_370),
.C(n_333),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_898),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_SL g981 ( 
.A(n_897),
.B(n_228),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_825),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_739),
.B(n_612),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_893),
.B(n_687),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_838),
.A2(n_648),
.B(n_626),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_846),
.A2(n_648),
.B(n_626),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_886),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_739),
.B(n_612),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_798),
.B(n_687),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_846),
.A2(n_648),
.B(n_626),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_798),
.B(n_711),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_802),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_861),
.A2(n_713),
.B(n_711),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_743),
.A2(n_713),
.B(n_393),
.C(n_537),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_853),
.B(n_697),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_861),
.A2(n_648),
.B(n_626),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_826),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_754),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_853),
.B(n_697),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_880),
.B(n_651),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_847),
.B(n_303),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_789),
.B(n_750),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_783),
.A2(n_537),
.B(n_529),
.C(n_539),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_757),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_782),
.B(n_651),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_821),
.A2(n_656),
.B(n_651),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_761),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_793),
.B(n_651),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_894),
.A2(n_666),
.B(n_656),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_783),
.A2(n_554),
.B(n_537),
.C(n_539),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_894),
.A2(n_666),
.B(n_656),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_793),
.B(n_656),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_852),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_895),
.A2(n_674),
.B(n_666),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_865),
.A2(n_318),
.B1(n_385),
.B2(n_380),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_776),
.A2(n_308),
.B1(n_377),
.B2(n_372),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_868),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_895),
.A2(n_674),
.B(n_666),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_828),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_800),
.B(n_674),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_795),
.A2(n_681),
.B(n_674),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_800),
.B(n_681),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_802),
.B(n_612),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_802),
.B(n_612),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_795),
.A2(n_684),
.B(n_681),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_806),
.A2(n_684),
.B(n_681),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_845),
.B(n_684),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_806),
.A2(n_701),
.B(n_684),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_845),
.B(n_701),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_748),
.B(n_303),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_899),
.A2(n_330),
.B1(n_394),
.B2(n_356),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_809),
.A2(n_701),
.B(n_504),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_809),
.A2(n_701),
.B(n_657),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_864),
.B(n_661),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_811),
.A2(n_657),
.B(n_638),
.Y(n_1035)
);

NOR2x1p5_ASAP7_75t_SL g1036 ( 
.A(n_813),
.B(n_638),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_661),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_811),
.A2(n_509),
.B(n_508),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_789),
.B(n_537),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_758),
.B(n_539),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_543),
.B(n_539),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_740),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_854),
.A2(n_545),
.B(n_543),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_785),
.B(n_245),
.Y(n_1044)
);

NOR2x1p5_ASAP7_75t_L g1045 ( 
.A(n_742),
.B(n_319),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_771),
.B(n_303),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_891),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_785),
.A2(n_563),
.B(n_559),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_878),
.A2(n_563),
.B(n_559),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_896),
.A2(n_336),
.B(n_396),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_758),
.B(n_543),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_767),
.A2(n_563),
.B(n_559),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_831),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_767),
.A2(n_563),
.B(n_559),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_758),
.B(n_543),
.Y(n_1055)
);

CKINVDCx10_ASAP7_75t_R g1056 ( 
.A(n_757),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_849),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_773),
.A2(n_554),
.B(n_553),
.C(n_546),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_851),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_758),
.B(n_787),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_787),
.B(n_545),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_855),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_837),
.B(n_248),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_893),
.B(n_332),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_777),
.B(n_337),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_858),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_787),
.B(n_545),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_774),
.A2(n_554),
.B(n_553),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_787),
.B(n_545),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_780),
.A2(n_277),
.B1(n_369),
.B2(n_367),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_837),
.B(n_824),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_787),
.B(n_546),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_791),
.A2(n_276),
.B1(n_365),
.B2(n_360),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_774),
.A2(n_554),
.B(n_553),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_759),
.A2(n_553),
.B(n_546),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_843),
.A2(n_356),
.B1(n_394),
.B2(n_319),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_866),
.A2(n_508),
.B(n_509),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_772),
.B(n_260),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_879),
.B(n_339),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_764),
.A2(n_546),
.B(n_510),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_841),
.B(n_250),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_870),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_896),
.B(n_508),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_900),
.B(n_509),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_900),
.B(n_342),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_766),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_775),
.B(n_261),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_796),
.A2(n_887),
.B(n_883),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_824),
.B(n_830),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_830),
.B(n_510),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_844),
.B(n_510),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_889),
.B(n_514),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_796),
.A2(n_518),
.B(n_514),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_968),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_907),
.B(n_902),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_968),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_934),
.B(n_822),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_987),
.B(n_786),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_906),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_SL g1100 ( 
.A(n_923),
.B(n_319),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_SL g1101 ( 
.A1(n_904),
.A2(n_818),
.B1(n_873),
.B2(n_843),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_920),
.B(n_873),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1085),
.A2(n_827),
.B(n_738),
.C(n_841),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_912),
.A2(n_901),
.B(n_892),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_968),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_909),
.B(n_859),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1085),
.A2(n_890),
.B1(n_873),
.B2(n_827),
.Y(n_1107)
);

OAI22x1_ASAP7_75t_L g1108 ( 
.A1(n_1045),
.A2(n_857),
.B1(n_786),
.B2(n_881),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_980),
.A2(n_1065),
.B1(n_1047),
.B2(n_920),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1002),
.B(n_790),
.Y(n_1110)
);

BUFx8_ASAP7_75t_L g1111 ( 
.A(n_1042),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_SL g1112 ( 
.A(n_1065),
.B(n_343),
.C(n_347),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1050),
.A2(n_862),
.B(n_370),
.C(n_363),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_929),
.B(n_860),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_989),
.B(n_872),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1013),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_948),
.A2(n_862),
.B(n_888),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_932),
.B(n_876),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_908),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_950),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_SL g1121 ( 
.A1(n_1089),
.A2(n_885),
.B(n_819),
.C(n_848),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_938),
.B(n_779),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_939),
.A2(n_890),
.B1(n_808),
.B2(n_803),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_SL g1124 ( 
.A(n_942),
.B(n_251),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_938),
.B(n_781),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_944),
.A2(n_363),
.B1(n_333),
.B2(n_345),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_913),
.A2(n_834),
.B(n_832),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_910),
.B(n_799),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_995),
.A2(n_829),
.B1(n_330),
.B2(n_252),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_925),
.A2(n_518),
.B(n_514),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1017),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_968),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_953),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_982),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_952),
.B(n_254),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1032),
.A2(n_931),
.B(n_930),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_961),
.A2(n_269),
.B(n_345),
.C(n_357),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_992),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1017),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_963),
.B(n_70),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_925),
.A2(n_518),
.B(n_514),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_992),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_L g1143 ( 
.A1(n_1090),
.A2(n_518),
.B(n_514),
.C(n_358),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1066),
.B(n_518),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1082),
.B(n_511),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_916),
.A2(n_309),
.B(n_353),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_944),
.A2(n_348),
.B1(n_389),
.B2(n_388),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_992),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_1081),
.B(n_265),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_952),
.B(n_267),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_270),
.Y(n_1152)
);

OR2x6_ASAP7_75t_SL g1153 ( 
.A(n_1015),
.B(n_349),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_928),
.B(n_272),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_L g1155 ( 
.A(n_923),
.B(n_279),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1007),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_917),
.B(n_281),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_955),
.B(n_288),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_919),
.A2(n_325),
.B(n_352),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_915),
.A2(n_975),
.B(n_965),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1086),
.Y(n_1161)
);

CKINVDCx14_ASAP7_75t_R g1162 ( 
.A(n_1046),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_992),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_951),
.A2(n_334),
.B(n_294),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1079),
.B(n_359),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_949),
.A2(n_324),
.B(n_351),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1030),
.A2(n_362),
.B(n_368),
.C(n_371),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_911),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1004),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1071),
.A2(n_326),
.B1(n_297),
.B2(n_346),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_974),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_984),
.B(n_323),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_957),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_997),
.B(n_1019),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_926),
.A2(n_379),
.B1(n_328),
.B2(n_344),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_984),
.B(n_338),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_940),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_957),
.B(n_511),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_SL g1179 ( 
.A(n_981),
.B(n_290),
.C(n_302),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1053),
.B(n_511),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1078),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_957),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_964),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_956),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1001),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_974),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1039),
.A2(n_21),
.B(n_22),
.C(n_31),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_926),
.A2(n_962),
.B1(n_943),
.B2(n_914),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_941),
.B(n_305),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_958),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_999),
.B(n_304),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1057),
.B(n_511),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1059),
.B(n_511),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_511),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_SL g1195 ( 
.A(n_923),
.B(n_511),
.Y(n_1195)
);

AND2x6_ASAP7_75t_L g1196 ( 
.A(n_947),
.B(n_188),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_922),
.A2(n_179),
.B(n_173),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_967),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_924),
.A2(n_168),
.B(n_166),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_935),
.A2(n_156),
.B(n_155),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_971),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_966),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_970),
.B(n_1083),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1064),
.B(n_21),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1084),
.A2(n_154),
.B(n_151),
.C(n_146),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_978),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1077),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1044),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_1044),
.A2(n_143),
.B(n_125),
.C(n_114),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_943),
.B(n_33),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1060),
.A2(n_113),
.B(n_101),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_921),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1000),
.B(n_34),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1034),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1078),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_918),
.A2(n_35),
.B(n_37),
.C(n_40),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1063),
.B(n_96),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_962),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1037),
.Y(n_1219)
);

NAND2xp33_ASAP7_75t_R g1220 ( 
.A(n_1064),
.B(n_87),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_935),
.B(n_41),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1003),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1004),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1087),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_933),
.B(n_44),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_923),
.A2(n_83),
.B(n_72),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_979),
.B(n_44),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_1087),
.B(n_71),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1023),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1023),
.Y(n_1230)
);

NOR3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1070),
.B(n_47),
.C(n_48),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1056),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_979),
.A2(n_1091),
.B(n_1073),
.C(n_1016),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1031),
.B(n_50),
.Y(n_1234)
);

OA22x2_ASAP7_75t_L g1235 ( 
.A1(n_905),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1235)
);

NOR3xp33_ASAP7_75t_SL g1236 ( 
.A(n_933),
.B(n_53),
.C(n_57),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1008),
.B(n_58),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1031),
.A2(n_1076),
.B1(n_1005),
.B2(n_1040),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1076),
.A2(n_62),
.B(n_58),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1010),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1048),
.A2(n_61),
.B(n_1088),
.C(n_927),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_959),
.B(n_61),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_903),
.A2(n_1067),
.B1(n_1072),
.B2(n_1069),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_960),
.A2(n_994),
.B(n_1058),
.C(n_1051),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1055),
.A2(n_1061),
.B1(n_1027),
.B2(n_1012),
.Y(n_1245)
);

NOR2xp67_ASAP7_75t_L g1246 ( 
.A(n_1041),
.B(n_1043),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1020),
.A2(n_1022),
.B1(n_1029),
.B2(n_954),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1036),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_945),
.A2(n_946),
.B(n_996),
.C(n_973),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_993),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_SL g1251 ( 
.A(n_1024),
.B(n_988),
.C(n_977),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1038),
.B(n_1092),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1014),
.B(n_1018),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1024),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_977),
.A2(n_988),
.B1(n_983),
.B2(n_1011),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_983),
.B(n_1009),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1052),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_960),
.A2(n_1054),
.B(n_1074),
.C(n_1068),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1095),
.B(n_1006),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_L g1260 ( 
.A(n_1171),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1204),
.A2(n_1075),
.B(n_1049),
.C(n_990),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1188),
.A2(n_1035),
.B(n_1033),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1200),
.A2(n_1080),
.B(n_1021),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1202),
.B(n_985),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1233),
.A2(n_986),
.B(n_976),
.C(n_1093),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1203),
.B(n_1028),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1173),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1139),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1186),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1116),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1101),
.A2(n_1025),
.B1(n_1026),
.B2(n_936),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_SL g1274 ( 
.A(n_1178),
.B(n_969),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1258),
.A2(n_972),
.B(n_937),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1185),
.B(n_1098),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1218),
.B(n_1239),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1097),
.B(n_1185),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_SL g1279 ( 
.A1(n_1212),
.A2(n_1218),
.B(n_1126),
.C(n_1200),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

INVx3_ASAP7_75t_SL g1281 ( 
.A(n_1232),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_R g1282 ( 
.A(n_1134),
.B(n_1169),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1241),
.A2(n_1160),
.A3(n_1249),
.B(n_1188),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1255),
.A2(n_1127),
.B(n_1253),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1255),
.A2(n_1247),
.B(n_1141),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1174),
.B(n_1198),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1174),
.B(n_1206),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1124),
.A2(n_1162),
.B1(n_1109),
.B2(n_1110),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1247),
.A2(n_1130),
.B(n_1245),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1131),
.B(n_1165),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1119),
.B(n_1120),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1173),
.B(n_1182),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1103),
.A2(n_1243),
.B(n_1115),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1102),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1102),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1210),
.A2(n_1221),
.B(n_1126),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1182),
.B(n_1096),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_L g1298 ( 
.A1(n_1148),
.A2(n_1108),
.B1(n_1167),
.B2(n_1175),
.C(n_1113),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1124),
.B(n_1196),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1238),
.A2(n_1148),
.A3(n_1243),
.B1(n_1175),
.B2(n_1245),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1115),
.A2(n_1256),
.B(n_1106),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1096),
.B(n_1094),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1225),
.A2(n_1164),
.B(n_1237),
.C(n_1112),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1256),
.A2(n_1106),
.B(n_1252),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1133),
.B(n_1215),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1242),
.A2(n_1234),
.B1(n_1227),
.B2(n_1164),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1244),
.A2(n_1143),
.B(n_1250),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1256),
.A2(n_1155),
.B(n_1191),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1216),
.A2(n_1187),
.B(n_1231),
.C(n_1183),
.Y(n_1309)
);

AOI221xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1208),
.A2(n_1137),
.B1(n_1213),
.B2(n_1122),
.C(n_1125),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1209),
.A2(n_1201),
.B(n_1123),
.C(n_1152),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1145),
.A2(n_1180),
.B(n_1192),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1190),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1220),
.A2(n_1153),
.B1(n_1235),
.B2(n_1228),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1235),
.A2(n_1107),
.B1(n_1236),
.B2(n_1190),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1190),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1214),
.B(n_1219),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1180),
.A2(n_1193),
.B(n_1192),
.Y(n_1318)
);

OAI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1154),
.A2(n_1157),
.B1(n_1172),
.B2(n_1224),
.C(n_1215),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1179),
.A2(n_1170),
.B(n_1140),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1215),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1222),
.A2(n_1240),
.B(n_1205),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1114),
.A2(n_1118),
.B(n_1189),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_1151),
.Y(n_1324)
);

OAI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1150),
.A2(n_1129),
.B(n_1158),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1224),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1146),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1156),
.Y(n_1328)
);

AND2x2_ASAP7_75t_SL g1329 ( 
.A(n_1223),
.B(n_1140),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1178),
.A2(n_1251),
.B1(n_1257),
.B2(n_1228),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1224),
.B(n_1228),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1194),
.A2(n_1197),
.B(n_1199),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1166),
.A2(n_1211),
.B(n_1217),
.C(n_1135),
.Y(n_1333)
);

AO21x2_ASAP7_75t_L g1334 ( 
.A1(n_1121),
.A2(n_1246),
.B(n_1147),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1161),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1111),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1128),
.B(n_1196),
.Y(n_1337)
);

AOI221x1_ASAP7_75t_L g1338 ( 
.A1(n_1159),
.A2(n_1194),
.B1(n_1226),
.B2(n_1248),
.C(n_1254),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1254),
.A2(n_1144),
.B(n_1230),
.C(n_1229),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1105),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1144),
.A2(n_1163),
.B(n_1132),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1195),
.A2(n_1248),
.B(n_1163),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1138),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1132),
.A2(n_1149),
.B(n_1142),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1196),
.A2(n_1100),
.B(n_1230),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1196),
.A2(n_1229),
.B(n_1230),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1229),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1138),
.A2(n_1142),
.B(n_1149),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1142),
.A2(n_1181),
.B(n_1111),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1181),
.A2(n_1136),
.B(n_1117),
.Y(n_1350)
);

NOR4xp25_ASAP7_75t_L g1351 ( 
.A(n_1218),
.B(n_1187),
.C(n_1216),
.D(n_1183),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1204),
.A2(n_763),
.B1(n_1085),
.B2(n_628),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1204),
.A2(n_1085),
.B(n_763),
.C(n_628),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1200),
.A2(n_1216),
.B(n_1210),
.C(n_1103),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1101),
.A2(n_566),
.B1(n_538),
.B2(n_1162),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1099),
.B(n_865),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1097),
.B(n_820),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_763),
.B(n_1085),
.C(n_820),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1241),
.A2(n_1160),
.A3(n_1249),
.B(n_1188),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1095),
.B(n_902),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1139),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1203),
.A2(n_902),
.B1(n_842),
.B2(n_833),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1095),
.B(n_902),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1116),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1203),
.A2(n_902),
.B1(n_842),
.B2(n_833),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1241),
.A2(n_1160),
.A3(n_1249),
.B(n_1188),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1204),
.A2(n_1085),
.B(n_763),
.C(n_628),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1160),
.A2(n_1241),
.B(n_1249),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1185),
.B(n_1047),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1094),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1204),
.A2(n_1085),
.B(n_763),
.C(n_628),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1188),
.A2(n_1160),
.B(n_1243),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1168),
.Y(n_1378)
);

AOI211x1_ASAP7_75t_L g1379 ( 
.A1(n_1218),
.A2(n_1098),
.B(n_1239),
.C(n_1200),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1116),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1160),
.A2(n_1247),
.B(n_1207),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1095),
.B(n_902),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1116),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1241),
.A2(n_1160),
.A3(n_1249),
.B(n_1188),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1204),
.B(n_763),
.C(n_1085),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1168),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1204),
.A2(n_1085),
.B(n_763),
.C(n_628),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1168),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_SL g1395 ( 
.A(n_1111),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1203),
.A2(n_902),
.B1(n_842),
.B2(n_833),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1188),
.A2(n_1160),
.B(n_1243),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1185),
.B(n_1047),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1094),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1203),
.A2(n_902),
.B1(n_842),
.B2(n_833),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1188),
.A2(n_1160),
.B(n_1243),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1168),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1095),
.B(n_902),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1168),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1136),
.A2(n_1117),
.B(n_1104),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1188),
.A2(n_1160),
.B(n_1243),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_1232),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1168),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1116),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1188),
.A2(n_1160),
.B(n_1243),
.Y(n_1411)
);

AOI221x1_ASAP7_75t_L g1412 ( 
.A1(n_1204),
.A2(n_763),
.B1(n_1216),
.B2(n_1200),
.C(n_1218),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1203),
.A2(n_902),
.B1(n_842),
.B2(n_833),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1160),
.A2(n_603),
.B(n_751),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1111),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1111),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1168),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1270),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1277),
.A2(n_1299),
.B1(n_1388),
.B2(n_1364),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1388),
.A2(n_1352),
.B1(n_1277),
.B2(n_1298),
.Y(n_1420)
);

BUFx4_ASAP7_75t_SL g1421 ( 
.A(n_1336),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1281),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1314),
.A2(n_1296),
.B1(n_1299),
.B2(n_1377),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1286),
.B(n_1287),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1395),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1383),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1373),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1417),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1361),
.B(n_1365),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1353),
.A2(n_1391),
.B1(n_1375),
.B2(n_1371),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1291),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1412),
.A2(n_1369),
.B1(n_1413),
.B2(n_1396),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1410),
.Y(n_1433)
);

BUFx10_ASAP7_75t_L g1434 ( 
.A(n_1367),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1377),
.A2(n_1397),
.B1(n_1407),
.B2(n_1401),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1397),
.A2(n_1407),
.B1(n_1401),
.B2(n_1411),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1268),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1355),
.A2(n_1288),
.B1(n_1329),
.B2(n_1415),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1411),
.A2(n_1306),
.B1(n_1400),
.B2(n_1325),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1358),
.B(n_1305),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1359),
.A2(n_1303),
.B1(n_1379),
.B2(n_1400),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1269),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1408),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1324),
.A2(n_1320),
.B1(n_1330),
.B2(n_1319),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1280),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1306),
.A2(n_1315),
.B1(n_1382),
.B2(n_1403),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1315),
.A2(n_1330),
.B1(n_1276),
.B2(n_1300),
.Y(n_1447)
);

BUFx4_ASAP7_75t_SL g1448 ( 
.A(n_1416),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1380),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1290),
.A2(n_1398),
.B1(n_1337),
.B2(n_1362),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1293),
.A2(n_1357),
.B1(n_1304),
.B2(n_1405),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1294),
.A2(n_1317),
.B1(n_1339),
.B2(n_1311),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1295),
.B(n_1378),
.Y(n_1453)
);

OAI22x1_ASAP7_75t_L g1454 ( 
.A1(n_1345),
.A2(n_1292),
.B1(n_1313),
.B2(n_1331),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1283),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1408),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1390),
.A2(n_1393),
.B1(n_1409),
.B2(n_1402),
.Y(n_1457)
);

BUFx8_ASAP7_75t_L g1458 ( 
.A(n_1326),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1301),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1260),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1374),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1372),
.A2(n_1266),
.B1(n_1327),
.B2(n_1328),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1335),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1347),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1260),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1320),
.A2(n_1310),
.B1(n_1267),
.B2(n_1354),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1272),
.A2(n_1267),
.B1(n_1321),
.B2(n_1309),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1297),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1264),
.A2(n_1349),
.B1(n_1279),
.B2(n_1259),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1343),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1372),
.A2(n_1307),
.B1(n_1366),
.B2(n_1404),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1399),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1399),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_R g1475 ( 
.A1(n_1282),
.A2(n_1349),
.B1(n_1300),
.B2(n_1351),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1307),
.A2(n_1414),
.B1(n_1389),
.B2(n_1376),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1341),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1310),
.B(n_1323),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1399),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1308),
.A2(n_1345),
.B1(n_1351),
.B2(n_1333),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1340),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1363),
.A2(n_1368),
.B1(n_1262),
.B2(n_1300),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1343),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1340),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1346),
.B(n_1350),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1302),
.Y(n_1486)
);

BUFx8_ASAP7_75t_SL g1487 ( 
.A(n_1381),
.Y(n_1487)
);

INVx6_ASAP7_75t_L g1488 ( 
.A(n_1348),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1283),
.B(n_1360),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1334),
.A2(n_1322),
.B1(n_1262),
.B2(n_1342),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1322),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_L g1492 ( 
.A(n_1344),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_SL g1493 ( 
.A(n_1274),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1312),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1338),
.A2(n_1263),
.B1(n_1360),
.B2(n_1370),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1285),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1318),
.A2(n_1289),
.B1(n_1334),
.B2(n_1284),
.Y(n_1497)
);

CKINVDCx14_ASAP7_75t_R g1498 ( 
.A(n_1360),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1370),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1370),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1332),
.A2(n_1275),
.B1(n_1406),
.B2(n_1273),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1261),
.A2(n_1265),
.B1(n_1387),
.B2(n_1384),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1356),
.A2(n_1385),
.B1(n_1386),
.B2(n_1392),
.Y(n_1503)
);

INVx5_ASAP7_75t_L g1504 ( 
.A(n_1387),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1394),
.A2(n_1388),
.B1(n_763),
.B2(n_1352),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1271),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1271),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1286),
.B(n_934),
.Y(n_1509)
);

BUFx8_ASAP7_75t_L g1510 ( 
.A(n_1278),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1283),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1373),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1271),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1271),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1271),
.Y(n_1516)
);

INVx6_ASAP7_75t_L g1517 ( 
.A(n_1271),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1417),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1270),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1277),
.A2(n_1299),
.B1(n_942),
.B2(n_1218),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1286),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1417),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_1270),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1352),
.A2(n_1388),
.B1(n_1353),
.B2(n_1375),
.Y(n_1526)
);

INVx6_ASAP7_75t_L g1527 ( 
.A(n_1271),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1417),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1283),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1281),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1286),
.B(n_934),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1532)
);

BUFx8_ASAP7_75t_L g1533 ( 
.A(n_1278),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1271),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1283),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1271),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1271),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1395),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1373),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1270),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1271),
.Y(n_1542)
);

CKINVDCx14_ASAP7_75t_R g1543 ( 
.A(n_1336),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1388),
.A2(n_763),
.B1(n_1352),
.B2(n_1204),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1352),
.A2(n_1388),
.B1(n_1353),
.B2(n_1375),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1271),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1277),
.A2(n_1299),
.B1(n_942),
.B2(n_1218),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1271),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1417),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1537),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1501),
.A2(n_1503),
.B(n_1497),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1424),
.B(n_1522),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1455),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1501),
.A2(n_1503),
.B(n_1497),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1455),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1491),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1489),
.B(n_1511),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1494),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1496),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1472),
.A2(n_1476),
.B(n_1482),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1529),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1529),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1498),
.B(n_1439),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1535),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1502),
.A2(n_1485),
.B(n_1472),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1459),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1459),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1522),
.B(n_1427),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1454),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1498),
.B(n_1439),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1442),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1496),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1435),
.A2(n_1436),
.B(n_1430),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1485),
.A2(n_1477),
.B(n_1476),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1496),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1496),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_SL g1578 ( 
.A1(n_1466),
.A2(n_1444),
.B(n_1526),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1490),
.A2(n_1500),
.B(n_1482),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1499),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1440),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1419),
.B(n_1447),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1445),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1428),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1504),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1437),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1478),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1480),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1441),
.Y(n_1589)
);

AO31x2_ASAP7_75t_L g1590 ( 
.A1(n_1545),
.A2(n_1452),
.A3(n_1468),
.B(n_1432),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1518),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1451),
.A2(n_1462),
.B(n_1435),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1523),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1528),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1436),
.A2(n_1495),
.B(n_1432),
.Y(n_1595)
);

INVx8_ASAP7_75t_L g1596 ( 
.A(n_1473),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1419),
.B(n_1447),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1483),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1451),
.A2(n_1462),
.B(n_1505),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1505),
.A2(n_1423),
.B(n_1446),
.Y(n_1600)
);

AO21x1_ASAP7_75t_SL g1601 ( 
.A1(n_1423),
.A2(n_1420),
.B(n_1446),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1492),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1549),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1450),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1426),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1457),
.A2(n_1420),
.B(n_1469),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1495),
.A2(n_1470),
.B(n_1464),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1487),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1426),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1426),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1506),
.A2(n_1512),
.B(n_1521),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1463),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1470),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1513),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1493),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1431),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1488),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1520),
.B(n_1547),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1488),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1520),
.B(n_1547),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1540),
.B(n_1429),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1467),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1475),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_R g1624 ( 
.A(n_1422),
.B(n_1530),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1506),
.B(n_1512),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1510),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1471),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1481),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1510),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1509),
.B(n_1531),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1492),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1521),
.A2(n_1532),
.B(n_1544),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1525),
.B(n_1532),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1525),
.B(n_1544),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1453),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1484),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1486),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1533),
.B(n_1548),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1533),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1461),
.A2(n_1479),
.B(n_1474),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1625),
.A2(n_1633),
.B1(n_1634),
.B2(n_1611),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1608),
.A2(n_1438),
.B1(n_1543),
.B2(n_1539),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1580),
.B(n_1449),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1595),
.B(n_1599),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1584),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1580),
.B(n_1514),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1578),
.A2(n_1465),
.B(n_1460),
.C(n_1543),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_R g1649 ( 
.A(n_1611),
.B(n_1425),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_SL g1650 ( 
.A1(n_1623),
.A2(n_1421),
.B(n_1448),
.C(n_1458),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1581),
.B(n_1515),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1613),
.A2(n_1434),
.B(n_1458),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1574),
.A2(n_1546),
.B(n_1542),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1578),
.A2(n_1508),
.B1(n_1507),
.B2(n_1448),
.C(n_1421),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1552),
.B(n_1622),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1556),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1517),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1569),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1608),
.A2(n_1517),
.B1(n_1433),
.B2(n_1538),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1625),
.B(n_1516),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1626),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1550),
.B(n_1516),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1564),
.B(n_1516),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1564),
.B(n_1571),
.Y(n_1664)
);

OA21x2_ASAP7_75t_L g1665 ( 
.A1(n_1613),
.A2(n_1434),
.B(n_1433),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1571),
.B(n_1538),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1633),
.A2(n_1443),
.B1(n_1456),
.B2(n_1524),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1618),
.A2(n_1527),
.B1(n_1538),
.B2(n_1418),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1611),
.A2(n_1527),
.B(n_1524),
.C(n_1519),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1602),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1588),
.B(n_1541),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1561),
.B(n_1570),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1604),
.B(n_1589),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1611),
.B(n_1618),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1630),
.B(n_1636),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1584),
.B(n_1586),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1558),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1599),
.B(n_1592),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1557),
.B(n_1630),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1605),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1636),
.B(n_1621),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1632),
.A2(n_1600),
.B(n_1620),
.C(n_1597),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1614),
.B(n_1587),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1592),
.B(n_1566),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1620),
.A2(n_1582),
.B(n_1597),
.C(n_1572),
.Y(n_1685)
);

A2O1A1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1632),
.A2(n_1600),
.B(n_1582),
.C(n_1566),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1606),
.A2(n_1631),
.B(n_1617),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1591),
.B(n_1593),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1587),
.B(n_1627),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1579),
.B(n_1575),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1559),
.B(n_1573),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1573),
.B(n_1576),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1626),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1583),
.B(n_1612),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1628),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1629),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1561),
.B(n_1607),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1567),
.A2(n_1568),
.B(n_1561),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1590),
.B(n_1594),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1551),
.A2(n_1554),
.B(n_1585),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1606),
.A2(n_1631),
.B(n_1617),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1601),
.A2(n_1561),
.B1(n_1640),
.B2(n_1629),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1685),
.A2(n_1640),
.B(n_1598),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1658),
.B(n_1607),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1672),
.B(n_1579),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1646),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1664),
.B(n_1607),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1553),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1692),
.B(n_1576),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1674),
.A2(n_1649),
.B1(n_1645),
.B2(n_1698),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1679),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1692),
.B(n_1577),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1665),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1649),
.A2(n_1602),
.B1(n_1601),
.B2(n_1635),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1718)
);

INVxp33_ASAP7_75t_L g1719 ( 
.A(n_1662),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1700),
.B(n_1590),
.Y(n_1720)
);

NOR2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1694),
.B(n_1602),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1678),
.B(n_1553),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1684),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1645),
.B(n_1555),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1645),
.B(n_1560),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1699),
.B(n_1562),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1675),
.B(n_1590),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1656),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1642),
.A2(n_1590),
.B1(n_1615),
.B2(n_1619),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1688),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1676),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1686),
.B(n_1563),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_1698),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1710),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1712),
.A2(n_1703),
.B1(n_1671),
.B2(n_1660),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1710),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1704),
.B(n_1682),
.C(n_1703),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1717),
.A2(n_1682),
.B1(n_1697),
.B2(n_1661),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1726),
.Y(n_1741)
);

AND2x4_ASAP7_75t_SL g1742 ( 
.A(n_1717),
.B(n_1670),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1712),
.A2(n_1671),
.B1(n_1660),
.B2(n_1668),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1704),
.A2(n_1673),
.B1(n_1643),
.B2(n_1654),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1710),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1707),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1729),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1726),
.Y(n_1748)
);

CKINVDCx14_ASAP7_75t_R g1749 ( 
.A(n_1735),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1726),
.Y(n_1750)
);

INVx5_ASAP7_75t_SL g1751 ( 
.A(n_1711),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1735),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1734),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1723),
.B(n_1693),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1719),
.B(n_1667),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1711),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1701),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1711),
.Y(n_1759)
);

AOI211x1_ASAP7_75t_L g1760 ( 
.A1(n_1734),
.A2(n_1653),
.B(n_1683),
.C(n_1681),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1706),
.B(n_1701),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1708),
.B(n_1690),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1707),
.Y(n_1764)
);

OAI33xp33_ASAP7_75t_L g1765 ( 
.A1(n_1705),
.A2(n_1689),
.A3(n_1659),
.B1(n_1651),
.B2(n_1603),
.B3(n_1695),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1690),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1708),
.B(n_1690),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1705),
.B(n_1691),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1565),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1730),
.A2(n_1652),
.B1(n_1666),
.B2(n_1663),
.Y(n_1770)
);

AND2x2_ASAP7_75t_SL g1771 ( 
.A(n_1730),
.B(n_1652),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_L g1772 ( 
.A(n_1727),
.B(n_1669),
.C(n_1673),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1728),
.A2(n_1648),
.B(n_1702),
.C(n_1687),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.B(n_1652),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1716),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1728),
.B(n_1657),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1723),
.B(n_1732),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1761),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1769),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1769),
.Y(n_1782)
);

NOR2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1727),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1736),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1758),
.B(n_1720),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1736),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1738),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1738),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1745),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1768),
.B(n_1720),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1759),
.B(n_1755),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1709),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1753),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1746),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1756),
.B(n_1624),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1745),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1759),
.B(n_1722),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1776),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1760),
.B(n_1731),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1722),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_1733),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1747),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1760),
.B(n_1754),
.Y(n_1805)
);

OA21x2_ASAP7_75t_L g1806 ( 
.A1(n_1741),
.A2(n_1714),
.B(n_1716),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1747),
.Y(n_1807)
);

AOI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1740),
.A2(n_1725),
.B(n_1724),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1754),
.B(n_1772),
.Y(n_1809)
);

INVx4_ASAP7_75t_L g1810 ( 
.A(n_1742),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1772),
.B(n_1731),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1755),
.B(n_1733),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1761),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1763),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1806),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1810),
.B(n_1763),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1806),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1785),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1784),
.B(n_1752),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1785),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1810),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1784),
.B(n_1752),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1787),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1803),
.B(n_1767),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1787),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1809),
.B(n_1775),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1806),
.Y(n_1828)
);

NOR2x1p5_ASAP7_75t_SL g1829 ( 
.A(n_1778),
.B(n_1761),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1789),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1790),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1801),
.B(n_1749),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1803),
.B(n_1812),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1795),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1790),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1806),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1792),
.B(n_1764),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1778),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1796),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1812),
.B(n_1767),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1808),
.A2(n_1650),
.B(n_1740),
.C(n_1744),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1792),
.B(n_1775),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1805),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1813),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1813),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1791),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1798),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1793),
.B(n_1741),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1798),
.Y(n_1851)
);

INVxp33_ASAP7_75t_L g1852 ( 
.A(n_1797),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1804),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1793),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1804),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1793),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1800),
.B(n_1762),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1807),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1781),
.B(n_1762),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1819),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1841),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1833),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1816),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1819),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1852),
.B(n_1624),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1821),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1834),
.B(n_1802),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1816),
.Y(n_1868)
);

AOI211x1_ASAP7_75t_SL g1869 ( 
.A1(n_1827),
.A2(n_1773),
.B(n_1739),
.C(n_1783),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1835),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1827),
.B(n_1786),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1834),
.B(n_1802),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1821),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1814),
.B(n_1786),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1825),
.B(n_1793),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1835),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1854),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1824),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1838),
.B(n_1782),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1825),
.B(n_1779),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1842),
.B(n_1779),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1845),
.B(n_1782),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1842),
.B(n_1822),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1824),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1816),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1826),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1822),
.B(n_1744),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1826),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1830),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1843),
.B(n_1777),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1830),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1831),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1843),
.B(n_1777),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1896)
);

INVx3_ASAP7_75t_SL g1897 ( 
.A(n_1850),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1870),
.B(n_1820),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_L g1899 ( 
.A1(n_1888),
.A2(n_1737),
.B(n_1771),
.Y(n_1899)
);

AOI321xp33_ASAP7_75t_L g1900 ( 
.A1(n_1891),
.A2(n_1743),
.A3(n_1770),
.B1(n_1837),
.B2(n_1828),
.C(n_1818),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1877),
.A2(n_1771),
.B1(n_1817),
.B2(n_1854),
.Y(n_1901)
);

AOI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1862),
.A2(n_1856),
.B(n_1823),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1897),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1861),
.B(n_1820),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1860),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1869),
.B(n_1817),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1883),
.A2(n_1856),
.B(n_1823),
.Y(n_1907)
);

AOI21xp33_ASAP7_75t_L g1908 ( 
.A1(n_1878),
.A2(n_1832),
.B(n_1831),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1884),
.B(n_1857),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1884),
.B(n_1838),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1894),
.A2(n_1771),
.B1(n_1897),
.B2(n_1871),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1860),
.Y(n_1912)
);

AOI21xp33_ASAP7_75t_L g1913 ( 
.A1(n_1878),
.A2(n_1836),
.B(n_1832),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1867),
.B(n_1859),
.Y(n_1914)
);

AO21x1_ASAP7_75t_L g1915 ( 
.A1(n_1863),
.A2(n_1828),
.B(n_1818),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1897),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1864),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1865),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1874),
.B(n_1661),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1871),
.B(n_1874),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1864),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1867),
.B(n_1859),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1876),
.B(n_1844),
.Y(n_1923)
);

OAI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1876),
.A2(n_1850),
.B(n_1829),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1906),
.A2(n_1863),
.B(n_1868),
.C(n_1886),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_SL g1926 ( 
.A1(n_1903),
.A2(n_1886),
.B(n_1868),
.C(n_1893),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1919),
.B(n_1872),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1916),
.B(n_1872),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1918),
.B(n_1850),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1916),
.B(n_1895),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1899),
.A2(n_1896),
.B1(n_1895),
.B2(n_1875),
.Y(n_1931)
);

OAI21xp33_ASAP7_75t_L g1932 ( 
.A1(n_1910),
.A2(n_1896),
.B(n_1880),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1900),
.B(n_1650),
.C(n_1892),
.D(n_1890),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1904),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1911),
.A2(n_1880),
.B1(n_1892),
.B2(n_1890),
.C(n_1889),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1918),
.B(n_1875),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1898),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1920),
.B(n_1697),
.Y(n_1938)
);

AOI21xp33_ASAP7_75t_SL g1939 ( 
.A1(n_1902),
.A2(n_1844),
.B(n_1639),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1923),
.B(n_1909),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1907),
.B(n_1881),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1911),
.A2(n_1901),
.B1(n_1922),
.B2(n_1914),
.Y(n_1942)
);

AO21x1_ASAP7_75t_L g1943 ( 
.A1(n_1908),
.A2(n_1873),
.B(n_1866),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1924),
.A2(n_1850),
.B1(n_1881),
.B2(n_1882),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1905),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1933),
.A2(n_1928),
.B1(n_1938),
.B2(n_1943),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1934),
.Y(n_1947)
);

NOR2xp67_ASAP7_75t_L g1948 ( 
.A(n_1936),
.B(n_1912),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1928),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1937),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1940),
.Y(n_1951)
);

AOI322xp5_ASAP7_75t_L g1952 ( 
.A1(n_1942),
.A2(n_1913),
.A3(n_1921),
.B1(n_1917),
.B2(n_1818),
.C1(n_1828),
.C2(n_1837),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1944),
.B(n_1931),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1929),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1930),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1945),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1941),
.A2(n_1882),
.B1(n_1751),
.B2(n_1799),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1932),
.B(n_1866),
.Y(n_1958)
);

AOI322xp5_ASAP7_75t_L g1959 ( 
.A1(n_1946),
.A2(n_1927),
.A3(n_1933),
.B1(n_1926),
.B2(n_1837),
.C1(n_1873),
.C2(n_1879),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1949),
.B(n_1939),
.Y(n_1960)
);

NOR2x1_ASAP7_75t_L g1961 ( 
.A(n_1948),
.B(n_1925),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1954),
.B(n_1935),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1947),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1951),
.B(n_1915),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1953),
.B(n_1879),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1953),
.A2(n_1893),
.B1(n_1889),
.B2(n_1887),
.C(n_1885),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1955),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1958),
.B(n_1885),
.Y(n_1968)
);

AOI211xp5_ASAP7_75t_L g1969 ( 
.A1(n_1950),
.A2(n_1887),
.B(n_1641),
.C(n_1765),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1958),
.B1(n_1956),
.B2(n_1957),
.C(n_1952),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1962),
.A2(n_1748),
.B1(n_1750),
.B2(n_1858),
.C(n_1851),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1959),
.B(n_1836),
.Y(n_1972)
);

AOI31xp33_ASAP7_75t_L g1973 ( 
.A1(n_1961),
.A2(n_1644),
.A3(n_1647),
.B(n_1680),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_L g1974 ( 
.A(n_1960),
.B(n_1721),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1965),
.A2(n_1748),
.B1(n_1750),
.B2(n_1855),
.Y(n_1975)
);

OAI221xp5_ASAP7_75t_L g1976 ( 
.A1(n_1970),
.A2(n_1967),
.B1(n_1966),
.B2(n_1963),
.C(n_1969),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1974),
.A2(n_1968),
.B1(n_1858),
.B2(n_1855),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1972),
.A2(n_1851),
.B1(n_1849),
.B2(n_1840),
.C(n_1839),
.Y(n_1978)
);

AOI222xp33_ASAP7_75t_L g1979 ( 
.A1(n_1971),
.A2(n_1829),
.B1(n_1849),
.B2(n_1840),
.C1(n_1847),
.C2(n_1846),
.Y(n_1979)
);

NAND3xp33_ASAP7_75t_L g1980 ( 
.A(n_1973),
.B(n_1846),
.C(n_1839),
.Y(n_1980)
);

AOI222xp33_ASAP7_75t_L g1981 ( 
.A1(n_1975),
.A2(n_1847),
.B1(n_1846),
.B2(n_1839),
.C1(n_1848),
.C2(n_1853),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1973),
.B(n_1847),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1977),
.B(n_1982),
.Y(n_1983)
);

XNOR2xp5_ASAP7_75t_L g1984 ( 
.A(n_1976),
.B(n_1641),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1980),
.Y(n_1985)
);

NAND4xp75_ASAP7_75t_L g1986 ( 
.A(n_1978),
.B(n_1979),
.C(n_1981),
.D(n_1774),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1976),
.B(n_1848),
.Y(n_1987)
);

OAI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1976),
.A2(n_1848),
.B1(n_1853),
.B2(n_1615),
.Y(n_1988)
);

NOR2x1_ASAP7_75t_L g1989 ( 
.A(n_1983),
.B(n_1638),
.Y(n_1989)
);

OR3x2_ASAP7_75t_L g1990 ( 
.A(n_1987),
.B(n_1596),
.C(n_1637),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1985),
.B(n_1788),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1984),
.A2(n_1853),
.B1(n_1638),
.B2(n_1799),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1991),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1993),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1994),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1994),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1995),
.A2(n_1990),
.B1(n_1992),
.B2(n_1986),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1996),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1998),
.Y(n_1999)
);

AO22x2_ASAP7_75t_L g2000 ( 
.A1(n_1997),
.A2(n_1989),
.B1(n_1988),
.B2(n_1638),
.Y(n_2000)
);

AOI21xp33_ASAP7_75t_L g2001 ( 
.A1(n_1999),
.A2(n_1596),
.B(n_1638),
.Y(n_2001)
);

AOI21xp33_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_2000),
.B(n_1596),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_2002),
.Y(n_2003)
);

OAI221xp5_ASAP7_75t_R g2004 ( 
.A1(n_2003),
.A2(n_1596),
.B1(n_1799),
.B2(n_1610),
.C(n_1609),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_2004),
.A2(n_1596),
.B1(n_1799),
.B2(n_1794),
.Y(n_2005)
);


endmodule