module real_jpeg_1824_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_286;
wire n_166;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_24),
.B1(n_28),
.B2(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_36),
.B1(n_68),
.B2(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_2),
.A2(n_36),
.B1(n_48),
.B2(n_53),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_30),
.B1(n_33),
.B2(n_140),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_3),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_3),
.A2(n_24),
.B1(n_28),
.B2(n_140),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_48),
.B1(n_53),
.B2(n_140),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_68),
.B1(n_69),
.B2(n_140),
.Y(n_229)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_22),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_4),
.B(n_28),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_33),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_67),
.C(n_69),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_4),
.A2(n_48),
.B1(n_53),
.B2(n_133),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_46),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_103),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_65),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_4),
.A2(n_28),
.B(n_182),
.Y(n_248)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_24),
.B1(n_28),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_32),
.B1(n_48),
.B2(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_32),
.B1(n_68),
.B2(n_69),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_30),
.B1(n_33),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_48),
.B1(n_53),
.B2(n_61),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_8),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_8),
.A2(n_24),
.B1(n_28),
.B2(n_61),
.Y(n_159)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_30),
.B1(n_33),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_24),
.B1(n_28),
.B2(n_94),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_11),
.A2(n_48),
.B1(n_53),
.B2(n_94),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_94),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_30),
.B1(n_33),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_12),
.A2(n_24),
.B1(n_28),
.B2(n_92),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_12),
.A2(n_48),
.B1(n_53),
.B2(n_92),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_92),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_14),
.A2(n_30),
.B1(n_33),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_14),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_14),
.A2(n_48),
.B1(n_53),
.B2(n_63),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_14),
.A2(n_24),
.B1(n_28),
.B2(n_63),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_336),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_81),
.B(n_333),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_20),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_21),
.A2(n_38),
.B(n_93),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_35),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_22),
.A2(n_29),
.B(n_37),
.Y(n_336)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_23),
.A2(n_38),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_23),
.A2(n_38),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_23),
.A2(n_38),
.B1(n_91),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_23),
.A2(n_38),
.B1(n_139),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_23),
.A2(n_34),
.B(n_60),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_24),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_24),
.A2(n_27),
.B(n_132),
.C(n_134),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_24),
.B(n_50),
.C(n_53),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_26),
.B(n_28),
.C(n_30),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_29),
.Y(n_290)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_30),
.B(n_133),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_38),
.A2(n_62),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_38),
.A2(n_80),
.B(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_40),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_77),
.C(n_78),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_41),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_59),
.C(n_64),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_42),
.A2(n_64),
.B1(n_312),
.B2(n_323),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_42),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_43),
.A2(n_57),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_47),
.B(n_57),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_57),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_46),
.B(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_46),
.A2(n_56),
.B1(n_137),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_46),
.A2(n_56),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_47),
.A2(n_54),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_47),
.A2(n_57),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_47),
.A2(n_57),
.B1(n_168),
.B2(n_248),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_53),
.B1(n_67),
.B2(n_72),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_48),
.A2(n_51),
.B(n_181),
.C(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_48),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_57),
.A2(n_96),
.B(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_59),
.B(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_64),
.A2(n_309),
.B1(n_310),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_64),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_64),
.B(n_309),
.C(n_313),
.Y(n_318)
);

OAI21x1_ASAP7_75t_R g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_75),
.Y(n_64)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_65),
.B(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_65),
.A2(n_73),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_65),
.A2(n_73),
.B1(n_215),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_66),
.B(n_76),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_66)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_69),
.B(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_73),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_76),
.A2(n_122),
.B(n_150),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_77),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_327),
.B(n_332),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_301),
.B(n_324),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_278),
.B(n_300),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_162),
.B(n_277),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_141),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_86),
.B(n_141),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_113),
.C(n_124),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_87),
.B(n_113),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_97),
.B2(n_98),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_95),
.C(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_99),
.B(n_108),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_106),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_102),
.B(n_117),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_100),
.A2(n_106),
.B(n_117),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_100),
.A2(n_102),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_101),
.A2(n_116),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_101),
.A2(n_103),
.B1(n_133),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_101),
.A2(n_103),
.B1(n_229),
.B2(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_102),
.A2(n_119),
.B(n_130),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_110),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_109),
.A2(n_122),
.B1(n_177),
.B2(n_250),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_111),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_123),
.B(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_124),
.B(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.C(n_138),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_125),
.A2(n_126),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_135),
.B(n_138),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_161),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_153),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_145),
.B(n_153),
.C(n_161),
.Y(n_299)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_147),
.B(n_149),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_147),
.A2(n_151),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_147),
.A2(n_286),
.B(n_288),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_160),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_159),
.Y(n_296)
);

AOI321xp33_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_258),
.A3(n_269),
.B1(n_275),
.B2(n_276),
.C(n_339),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_204),
.B(n_257),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_185),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_165),
.B(n_185),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.C(n_179),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_166),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_171),
.C(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_175),
.B(n_179),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_178),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_184),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_197),
.B2(n_198),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_199),
.C(n_202),
.Y(n_270)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_188),
.B(n_192),
.C(n_196),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_252),
.B(n_256),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_242),
.B(n_251),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_223),
.B(n_241),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_235),
.B(n_240),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_234),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_233),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.C(n_268),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_263),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_271),
.Y(n_275)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_299),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_299),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_284),
.C(n_292),
.Y(n_303)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_291),
.B2(n_292),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_295),
.B(n_298),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_297),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_305),
.CI(n_306),
.CON(n_304),
.SN(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_305),
.C(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_315),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_304),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_304),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_313),
.A2(n_314),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_318),
.C(n_320),
.Y(n_328)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_317),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule