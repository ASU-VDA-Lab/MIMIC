module fake_jpeg_31505_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_22),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_30),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_4),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_34),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_58),
.Y(n_68)
);

AND2x4_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_45),
.B1(n_52),
.B2(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_72),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_52),
.B(n_13),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_14),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_76),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_65),
.B1(n_74),
.B2(n_68),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_67),
.B(n_70),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_21),
.B(n_23),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_24),
.Y(n_88)
);


endmodule