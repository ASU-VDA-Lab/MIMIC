module real_jpeg_25090_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_26),
.B1(n_34),
.B2(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_1),
.A2(n_49),
.B1(n_61),
.B2(n_66),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_1),
.A2(n_49),
.B1(n_70),
.B2(n_136),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_61),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_84),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_26),
.B1(n_34),
.B2(n_84),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_58),
.B1(n_61),
.B2(n_66),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_58),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_5),
.A2(n_26),
.B1(n_34),
.B2(n_58),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_111),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_7),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_7),
.A2(n_61),
.B1(n_66),
.B2(n_162),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_162),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_7),
.A2(n_26),
.B1(n_34),
.B2(n_162),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_39),
.B1(n_61),
.B2(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_39),
.B1(n_70),
.B2(n_109),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_8),
.A2(n_26),
.B1(n_34),
.B2(n_39),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_57),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_61),
.B1(n_66),
.B2(n_72),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_72),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_11),
.A2(n_26),
.B1(n_34),
.B2(n_72),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_12),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_12),
.A2(n_61),
.B1(n_66),
.B2(n_108),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_108),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_12),
.A2(n_26),
.B1(n_34),
.B2(n_108),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_13),
.B(n_135),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_13),
.B(n_60),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_13),
.B(n_40),
.C(n_80),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_13),
.A2(n_61),
.B1(n_66),
.B2(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_13),
.B(n_126),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_214),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_13),
.B(n_26),
.C(n_45),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_13),
.A2(n_25),
.B(n_274),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_15),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_15),
.A2(n_35),
.B1(n_61),
.B2(n_66),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_15),
.A2(n_35),
.B1(n_57),
.B2(n_135),
.Y(n_351)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_16),
.B(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_16),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_347),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_138),
.A3(n_152),
.B(n_331),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_115),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_21),
.B(n_115),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_22),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_23),
.A2(n_24),
.B(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_24),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_33),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_96),
.B1(n_97),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_25),
.A2(n_190),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_25),
.B(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_25),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_27),
.Y(n_191)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_32),
.B(n_214),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_34),
.B(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_42),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_40),
.B(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_43),
.A2(n_50),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_43),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_43),
.A2(n_50),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_47),
.A2(n_87),
.B1(n_102),
.B2(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_173),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_47),
.A2(n_210),
.B(n_247),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_47),
.B(n_214),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_50),
.B(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_67),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_59),
.B1(n_112),
.B2(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_74)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_69),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_59),
.A2(n_112),
.B1(n_134),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_59),
.A2(n_67),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_60),
.A2(n_73),
.B1(n_107),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_60),
.A2(n_73),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_60),
.A2(n_73),
.B1(n_342),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_66),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_61),
.B(n_65),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_61),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_64),
.A2(n_66),
.A3(n_109),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_73),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_73),
.A2(n_114),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_78),
.A2(n_79),
.B1(n_128),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_78),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_78),
.A2(n_182),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_104),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_79),
.A2(n_166),
.B(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_87),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_87),
.A2(n_262),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_91),
.A2(n_92),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.C(n_105),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_93),
.A2(n_94),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_103),
.B(n_105),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_112),
.B(n_113),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_109),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_137),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_126),
.B1(n_181),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_125),
.A2(n_126),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_126),
.B(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_130),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_130),
.B(n_145),
.C(n_149),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_133),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_137),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_133),
.B(n_141),
.C(n_144),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_139),
.A2(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_140),
.B(n_151),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_146),
.Y(n_341)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_150),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_324),
.B(n_330),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_199),
.B(n_323),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_192),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_155),
.B(n_192),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_174),
.C(n_176),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_156),
.A2(n_157),
.B1(n_174),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_168),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_164),
.C(n_168),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_172),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_174),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_176),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_183),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_179),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_183),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_187),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_188),
.A2(n_285),
.B1(n_287),
.B2(n_289),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_194),
.B(n_195),
.C(n_198),
.Y(n_329)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_232),
.B(n_317),
.C(n_322),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_226),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_216),
.C(n_217),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_202),
.A2(n_203),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_208),
.C(n_212),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_216),
.B(n_217),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_227),
.B(n_230),
.C(n_231),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_311),
.B(n_316),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_263),
.B(n_310),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_252),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_237),
.B(n_252),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_245),
.C(n_249),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_245),
.A2(n_249),
.B1(n_250),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_259),
.C(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_304),
.B(n_309),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_282),
.B(n_303),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_276),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_276),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_292),
.B(n_302),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_290),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_288),
.B(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_297),
.B(n_301),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_340),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_352),
.Y(n_353)
);


endmodule