module fake_jpeg_19246_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx16_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_6),
.C(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_0),
.Y(n_14)
);

O2A1O1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_0),
.B(n_5),
.C(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_5),
.B(n_10),
.C(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_20),
.Y(n_26)
);

INVx5_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_26),
.Y(n_28)
);

BUFx24_ASAP7_75t_SL g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_21),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.C(n_11),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_15),
.B(n_16),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_18),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_12),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_30),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_37),
.Y(n_40)
);


endmodule