module fake_jpeg_31603_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_44),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_42),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_8),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_59),
.B(n_93),
.Y(n_134)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_31),
.B1(n_30),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_66),
.A2(n_72),
.B1(n_83),
.B2(n_19),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_36),
.B1(n_38),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_76),
.B1(n_86),
.B2(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_84),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_30),
.B1(n_34),
.B2(n_29),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_36),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_30),
.B1(n_34),
.B2(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_32),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_36),
.B1(n_28),
.B2(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_11),
.Y(n_108)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_34),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_34),
.B1(n_29),
.B2(n_26),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_45),
.B1(n_41),
.B2(n_25),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_55),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_127),
.C(n_93),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_39),
.CI(n_37),
.CON(n_97),
.SN(n_97)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_58),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_56),
.B1(n_73),
.B2(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_108),
.B(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_41),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_119),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_0),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_37),
.B1(n_19),
.B2(n_25),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_125),
.B1(n_56),
.B2(n_90),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_129),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_79),
.A2(n_37),
.B1(n_43),
.B2(n_19),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_69),
.A2(n_37),
.B(n_43),
.C(n_10),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_128),
.B(n_11),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_37),
.C(n_19),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_19),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_74),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_0),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_85),
.B1(n_81),
.B2(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_148),
.B1(n_150),
.B2(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_57),
.B1(n_73),
.B2(n_88),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_124),
.B1(n_99),
.B2(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_75),
.Y(n_201)
);

AO22x2_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_120),
.B1(n_95),
.B2(n_102),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_99),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_98),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_134),
.B(n_133),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_58),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_107),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_74),
.C(n_88),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_126),
.C(n_101),
.Y(n_176)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_166),
.B(n_133),
.Y(n_170)
);

AO22x1_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_88),
.B1(n_58),
.B2(n_75),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_1),
.B(n_3),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_75),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_200),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_175),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_182),
.B(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_173),
.A2(n_179),
.B1(n_181),
.B2(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_100),
.B1(n_119),
.B2(n_108),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_199),
.B1(n_155),
.B2(n_11),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_176),
.B(n_140),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_135),
.B1(n_148),
.B2(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_96),
.C(n_123),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_194),
.C(n_201),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_141),
.Y(n_185)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_R g186 ( 
.A(n_150),
.B(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_118),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_116),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_106),
.C(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_131),
.B1(n_106),
.B2(n_6),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_137),
.A2(n_151),
.B1(n_160),
.B2(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_160),
.B1(n_145),
.B2(n_161),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_202),
.A2(n_187),
.B1(n_189),
.B2(n_193),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_141),
.B(n_166),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_208),
.B(n_177),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_205),
.B(n_209),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_206),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_139),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_162),
.C(n_144),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_211),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_164),
.B1(n_140),
.B2(n_155),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_224),
.B1(n_14),
.B2(n_4),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_146),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_227),
.C(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_146),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_173),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_15),
.C(n_9),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_9),
.B1(n_14),
.B2(n_6),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_178),
.B1(n_189),
.B2(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_176),
.B(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_15),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_12),
.C(n_14),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_245),
.B(n_228),
.Y(n_265)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_179),
.B1(n_199),
.B2(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_242),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_240),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_171),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_248),
.C(n_252),
.Y(n_260)
);

AOI22x1_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_195),
.B1(n_178),
.B2(n_172),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_241),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_205),
.B1(n_217),
.B2(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_187),
.B1(n_6),
.B2(n_7),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_246),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_13),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_4),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_13),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_225),
.B1(n_209),
.B2(n_223),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_5),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_232),
.C(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_230),
.Y(n_270)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

OAI22x1_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_247),
.B1(n_215),
.B2(n_214),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_273),
.B1(n_277),
.B2(n_242),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_239),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_236),
.A2(n_221),
.B1(n_224),
.B2(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_222),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_235),
.A2(n_245),
.B1(n_247),
.B2(n_256),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_288),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_233),
.B(n_204),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_235),
.B1(n_254),
.B2(n_214),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_275),
.B1(n_266),
.B2(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_238),
.C(n_211),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_260),
.C(n_243),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_258),
.A2(n_214),
.B(n_208),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_240),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_263),
.B1(n_265),
.B2(n_259),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_273),
.B1(n_276),
.B2(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_231),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_300),
.C(n_301),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_302),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_258),
.B(n_271),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_278),
.B(n_287),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_285),
.C(n_243),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_252),
.C(n_239),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_284),
.B(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_299),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_291),
.B(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_313),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_282),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_268),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_300),
.B(n_296),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_295),
.B(n_309),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_250),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_295),
.C(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_316),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_316),
.A3(n_297),
.B1(n_279),
.B2(n_286),
.C1(n_216),
.C2(n_267),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_322),
.C(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_324),
.C(n_317),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_330),
.C(n_248),
.Y(n_336)
);

OAI321xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_216),
.A3(n_218),
.B1(n_229),
.B2(n_255),
.C(n_328),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_218),
.Y(n_338)
);


endmodule