module fake_netlist_1_541_n_45 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_45);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_7), .B(n_4), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_12), .B(n_1), .Y(n_19) );
OAI22xp5_ASAP7_75t_SL g20 ( .A1(n_13), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_15), .B(n_3), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_12), .B(n_14), .Y(n_23) );
OAI21x1_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_17), .B(n_6), .Y(n_24) );
OAI21x1_ASAP7_75t_SL g25 ( .A1(n_18), .A2(n_17), .B(n_6), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_26), .B(n_18), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_20), .B1(n_24), .B2(n_23), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_23), .Y(n_31) );
INVx2_ASAP7_75t_SL g32 ( .A(n_27), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
OR2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_5), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVxp33_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_33), .Y(n_38) );
OR2x2_ASAP7_75t_L g39 ( .A(n_38), .B(n_36), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g40 ( .A(n_38), .B(n_25), .Y(n_40) );
NAND2x1p5_ASAP7_75t_L g41 ( .A(n_37), .B(n_35), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g42 ( .A(n_39), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_41), .Y(n_43) );
NOR2xp33_ASAP7_75t_R g44 ( .A(n_42), .B(n_40), .Y(n_44) );
AOI322xp5_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_43), .A3(n_37), .B1(n_25), .B2(n_36), .C1(n_32), .C2(n_7), .Y(n_45) );
endmodule