module fake_jpeg_28780_n_499 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_499);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_499;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_25),
.A2(n_16),
.B1(n_8),
.B2(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_53),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_110)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_15),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_80),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_60),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_69),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_15),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_93),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_15),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_34),
.B(n_29),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_101),
.B(n_104),
.C(n_116),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_35),
.C(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_27),
.B1(n_22),
.B2(n_45),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_35),
.C(n_36),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_49),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_127),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_34),
.B(n_18),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_125),
.A2(n_157),
.B(n_102),
.C(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_33),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_139),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_46),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_137),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_46),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_91),
.B(n_48),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_60),
.B(n_48),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_71),
.B(n_47),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_60),
.B(n_47),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_52),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_53),
.B1(n_75),
.B2(n_82),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_158),
.B(n_186),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_183),
.B1(n_115),
.B2(n_131),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_189),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_88),
.B1(n_68),
.B2(n_72),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_67),
.B1(n_63),
.B2(n_90),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_164),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_167),
.Y(n_210)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_39),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_170),
.Y(n_245)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_185),
.Y(n_247)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_154),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_180),
.Y(n_237)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_199),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_101),
.A2(n_27),
.B1(n_45),
.B2(n_83),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_132),
.A2(n_66),
.B1(n_19),
.B2(n_52),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_85),
.B1(n_76),
.B2(n_100),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_21),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_168),
.B(n_161),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_108),
.B(n_117),
.C(n_129),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_95),
.C(n_156),
.Y(n_229)
);

NAND2xp33_ASAP7_75t_R g196 ( 
.A(n_143),
.B(n_92),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_198),
.C(n_131),
.Y(n_216)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_200),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_21),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_21),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_205),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_121),
.A2(n_64),
.B1(n_62),
.B2(n_21),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_185),
.B1(n_189),
.B2(n_163),
.Y(n_225)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_18),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_146),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_123),
.B1(n_111),
.B2(n_154),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_150),
.B1(n_155),
.B2(n_124),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_219),
.B1(n_15),
.B2(n_12),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_123),
.C(n_111),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_224),
.C(n_243),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_214),
.B(n_216),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_217),
.A2(n_222),
.B1(n_234),
.B2(n_239),
.Y(n_252)
);

OAI22x1_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_156),
.B1(n_147),
.B2(n_148),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_168),
.A2(n_148),
.B1(n_113),
.B2(n_145),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_86),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_247),
.B1(n_244),
.B2(n_168),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_164),
.C(n_180),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_160),
.B(n_173),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_182),
.A2(n_113),
.B1(n_118),
.B2(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_177),
.A2(n_118),
.B1(n_176),
.B2(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_18),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_18),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_220),
.B(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_258),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_287),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_165),
.B(n_171),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_263),
.B(n_268),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_257),
.A2(n_273),
.B(n_237),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_181),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_264),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_187),
.B1(n_179),
.B2(n_172),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_265),
.B1(n_271),
.B2(n_272),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_178),
.B(n_180),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_217),
.A2(n_170),
.B1(n_166),
.B2(n_169),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_204),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_276),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_197),
.B(n_184),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_210),
.B(n_188),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_269),
.B(n_270),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_219),
.A2(n_200),
.B1(n_208),
.B2(n_206),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_192),
.B1(n_164),
.B2(n_10),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_232),
.A2(n_198),
.B(n_2),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_223),
.A2(n_198),
.B1(n_2),
.B2(n_3),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_284),
.B1(n_237),
.B2(n_211),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_0),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_0),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_213),
.B(n_2),
.C(n_3),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_2),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_3),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_234),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_8),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_288),
.Y(n_311)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_12),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_214),
.A2(n_216),
.B(n_215),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_282),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_297),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_282),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_259),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_300),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_234),
.B1(n_222),
.B2(n_245),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_237),
.B1(n_236),
.B2(n_242),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_306),
.A2(n_319),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_256),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_288),
.Y(n_338)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_261),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_322),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_258),
.A3(n_269),
.B1(n_275),
.B2(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_234),
.Y(n_316)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_317),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_251),
.B(n_286),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_SL g319 ( 
.A(n_282),
.B(n_248),
.C(n_226),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_246),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_280),
.A2(n_211),
.B1(n_221),
.B2(n_250),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_242),
.B(n_241),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_221),
.B(n_226),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_262),
.B1(n_268),
.B2(n_284),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_328),
.A2(n_336),
.B1(n_345),
.B2(n_322),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_252),
.B1(n_271),
.B2(n_265),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_335),
.B1(n_341),
.B2(n_352),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_273),
.B1(n_289),
.B2(n_274),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_333),
.B(n_355),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_257),
.B1(n_264),
.B2(n_281),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_289),
.B1(n_278),
.B2(n_272),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_L g374 ( 
.A1(n_338),
.A2(n_346),
.B(n_311),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_279),
.B(n_277),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_340),
.A2(n_349),
.B(n_293),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_281),
.B1(n_276),
.B2(n_245),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_228),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_335),
.C(n_330),
.Y(n_359)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_301),
.A2(n_250),
.B(n_283),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_325),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_351),
.A2(n_320),
.B(n_297),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_296),
.A2(n_233),
.B1(n_4),
.B2(n_5),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_319),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_318),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_290),
.Y(n_355)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_358),
.A2(n_370),
.B1(n_379),
.B2(n_386),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_313),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_385),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_334),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_363),
.B(n_380),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_294),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_308),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_365),
.B(n_382),
.Y(n_393)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_351),
.B(n_350),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_312),
.Y(n_369)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_327),
.B1(n_339),
.B2(n_348),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_308),
.C(n_297),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_375),
.C(n_381),
.Y(n_395)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_384),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_374),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_354),
.C(n_348),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_327),
.B(n_299),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_328),
.A2(n_310),
.B1(n_315),
.B2(n_298),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_293),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_316),
.C(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_304),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_298),
.B1(n_291),
.B2(n_295),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_375),
.B(n_311),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_410),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_377),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_344),
.Y(n_396)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_332),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_399),
.B(n_412),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_379),
.A2(n_329),
.B1(n_339),
.B2(n_291),
.Y(n_400)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_350),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_402),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_365),
.B(n_331),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_407),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_332),
.C(n_304),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_383),
.C(n_371),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_369),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_386),
.A2(n_299),
.B1(n_345),
.B2(n_355),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_411),
.A2(n_358),
.B1(n_383),
.B2(n_372),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_381),
.B(n_352),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_382),
.C(n_372),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_430),
.C(n_412),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_404),
.A2(n_409),
.B1(n_392),
.B2(n_368),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_421),
.A2(n_399),
.B1(n_398),
.B2(n_388),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_406),
.A2(n_384),
.B1(n_373),
.B2(n_361),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_432),
.Y(n_449)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_370),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_428),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_360),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_367),
.C(n_326),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_393),
.B(n_357),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_393),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_433),
.B(n_445),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_397),
.B(n_404),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_438),
.B(n_448),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_418),
.A2(n_408),
.B1(n_397),
.B2(n_411),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_420),
.B1(n_428),
.B2(n_419),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_425),
.A2(n_389),
.B(n_402),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_403),
.C(n_401),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_429),
.C(n_321),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_394),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_441),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_413),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_420),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_444),
.A2(n_431),
.B1(n_417),
.B2(n_422),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_423),
.Y(n_445)
);

FAx1_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_403),
.CI(n_398),
.CON(n_447),
.SN(n_447)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_3),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_416),
.A2(n_388),
.B(n_376),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_452),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_454),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_464),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_309),
.B1(n_376),
.B2(n_429),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_462),
.B1(n_443),
.B2(n_449),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_303),
.C(n_302),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_439),
.C(n_434),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_441),
.A2(n_303),
.B1(n_356),
.B2(n_233),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_437),
.A2(n_356),
.B1(n_10),
.B2(n_11),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_448),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_11),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_3),
.B(n_4),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_4),
.Y(n_471)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_434),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_471),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_459),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_474),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_460),
.B(n_447),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_435),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_475),
.A2(n_454),
.B(n_447),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_470),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_481),
.B(n_471),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_467),
.C(n_468),
.Y(n_486)
);

OAI21x1_ASAP7_75t_SL g481 ( 
.A1(n_476),
.A2(n_453),
.B(n_458),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_473),
.A2(n_453),
.B(n_463),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_442),
.B(n_450),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_487),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_473),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_488),
.B(n_489),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_435),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_490),
.A2(n_480),
.B(n_482),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_SL g494 ( 
.A(n_493),
.B(n_478),
.C(n_477),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_494),
.A2(n_495),
.B(n_6),
.Y(n_496)
);

OAI311xp33_ASAP7_75t_L g495 ( 
.A1(n_492),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.C1(n_491),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_496),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_6),
.B(n_7),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_6),
.B(n_7),
.Y(n_499)
);


endmodule