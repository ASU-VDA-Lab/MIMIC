module fake_jpeg_30709_n_59 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_3),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_8),
.A3(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_24),
.Y(n_34)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_25),
.B(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_25),
.B1(n_23),
.B2(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_47),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AOI221xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_25),
.B1(n_23),
.B2(n_6),
.C(n_4),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_4),
.B1(n_5),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_35),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_53),
.B1(n_45),
.B2(n_5),
.Y(n_56)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_43),
.C(n_46),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI321xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_56),
.A3(n_55),
.B1(n_54),
.B2(n_52),
.C(n_12),
.Y(n_59)
);


endmodule