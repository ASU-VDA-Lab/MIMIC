module fake_jpeg_22376_n_56 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_56);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_33),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_5),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_6),
.B(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_11),
.B1(n_12),
.B2(n_21),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_17),
.B1(n_20),
.B2(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_44),
.B2(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_38),
.B1(n_41),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_46),
.B1(n_48),
.B2(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_40),
.B(n_39),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_49),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_42),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);


endmodule