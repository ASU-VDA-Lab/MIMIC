module real_jpeg_6409_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_0),
.A2(n_49),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_0),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_0),
.A2(n_243),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_0),
.A2(n_243),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_0),
.A2(n_129),
.B1(n_131),
.B2(n_243),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_1),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_123),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_123),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_1),
.A2(n_123),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_2),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_2),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_2),
.Y(n_290)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_2),
.Y(n_329)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_129),
.B1(n_131),
.B2(n_133),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_4),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_4),
.A2(n_133),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_133),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_63),
.B1(n_166),
.B2(n_170),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_5),
.A2(n_63),
.B1(n_195),
.B2(n_229),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_5),
.A2(n_63),
.B1(n_287),
.B2(n_393),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_256),
.B1(n_259),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_6),
.B(n_273),
.C(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_6),
.B(n_109),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_6),
.B(n_226),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_6),
.B(n_89),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_6),
.B(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_8),
.Y(n_501)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_9),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_10),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_10),
.A2(n_200),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_10),
.A2(n_200),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_10),
.A2(n_200),
.B1(n_353),
.B2(n_355),
.Y(n_352)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_76),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_93),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_93),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_48),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_14),
.A2(n_48),
.B1(n_221),
.B2(n_360),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_14),
.A2(n_48),
.B1(n_91),
.B2(n_194),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_15),
.A2(n_271),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_15),
.A2(n_298),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_15),
.A2(n_298),
.B1(n_367),
.B2(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_15),
.A2(n_49),
.B1(n_146),
.B2(n_298),
.Y(n_455)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_17),
.Y(n_505)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_500),
.B(n_502),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_204),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_203),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_150),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_24),
.B(n_150),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_134),
.B2(n_135),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_64),
.C(n_94),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_27),
.A2(n_136),
.B1(n_137),
.B2(n_149),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_27),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_27),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_46),
.B1(n_55),
.B2(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_28),
.A2(n_55),
.B1(n_57),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_28),
.A2(n_239),
.B(n_244),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_28),
.A2(n_37),
.B1(n_239),
.B2(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_29),
.B(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_29),
.A2(n_430),
.B(n_431),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_37),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_32),
.Y(n_409)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_37),
.B(n_262),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_37)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_38),
.Y(n_411)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_41),
.Y(n_354)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_42),
.Y(n_132)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_42),
.Y(n_169)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_44),
.Y(n_143)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_44),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_47),
.B(n_56),
.Y(n_197)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_55),
.A2(n_198),
.B(n_455),
.Y(n_470)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_56),
.B(n_199),
.Y(n_244)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_64),
.A2(n_65),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_64),
.A2(n_65),
.B1(n_94),
.B2(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_88),
.B(n_90),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_66),
.A2(n_255),
.B(n_263),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_66),
.A2(n_88),
.B1(n_297),
.B2(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_66),
.A2(n_263),
.B(n_340),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_66),
.A2(n_88),
.B1(n_436),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_67),
.A2(n_89),
.B1(n_156),
.B2(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_67),
.A2(n_89),
.B1(n_156),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_67),
.A2(n_89),
.B1(n_193),
.B2(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_67),
.B(n_264),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_69),
.Y(n_229)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_72),
.Y(n_344)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_73),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_78),
.A2(n_297),
.B(n_302),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_84),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_84),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_84),
.Y(n_361)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_85),
.Y(n_310)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_86),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_86),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_88),
.A2(n_302),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_89),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_118),
.B1(n_127),
.B2(n_128),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_96),
.A2(n_127),
.B1(n_128),
.B2(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_96),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_96),
.A2(n_127),
.B1(n_165),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_96),
.A2(n_127),
.B1(n_384),
.B2(n_434),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_102),
.Y(n_350)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_108),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_119),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22x1_ASAP7_75t_L g456 ( 
.A1(n_109),
.A2(n_163),
.B1(n_388),
.B2(n_457),
.Y(n_456)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_111),
.Y(n_370)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_116),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_116),
.Y(n_301)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_116),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g404 ( 
.A1(n_120),
.A2(n_405),
.A3(n_409),
.B1(n_410),
.B2(n_412),
.Y(n_404)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_127),
.B(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_127),
.A2(n_384),
.B(n_387),
.Y(n_383)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_131),
.A2(n_262),
.B(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_171),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_157),
.Y(n_368)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_163),
.A2(n_347),
.B(n_351),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_163),
.B(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_163),
.A2(n_351),
.B(n_473),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_169),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B(n_196),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_192),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_196),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_173),
.A2(n_192),
.B1(n_213),
.B2(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_184),
.B(n_186),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_186),
.B1(n_220),
.B2(n_224),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_174),
.A2(n_282),
.B(n_288),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_174),
.A2(n_262),
.B(n_288),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_174),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_414)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_175),
.B(n_291),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_175),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_175),
.A2(n_359),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_175),
.A2(n_418),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_182),
.Y(n_287)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_182),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_184),
.A2(n_315),
.B(n_319),
.Y(n_314)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_184),
.Y(n_395)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_192),
.Y(n_445)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_245),
.B(n_499),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_206),
.B(n_208),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_214),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_217),
.B(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_230),
.C(n_238),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_218),
.B(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_219),
.B(n_227),
.Y(n_467)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_220),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_226),
.Y(n_452)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_228),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_230),
.B(n_238),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_231),
.Y(n_457)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_241),
.B(n_262),
.Y(n_412)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_242),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_244),
.Y(n_431)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI311xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_439),
.A3(n_475),
.B1(n_493),
.C1(n_494),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_398),
.B(n_438),
.Y(n_248)
);

AO21x1_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_375),
.B(n_397),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_334),
.B(n_374),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_305),
.B(n_333),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_280),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_280),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_268),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_254),
.A2(n_268),
.B1(n_269),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g430 ( 
.A1(n_262),
.A2(n_406),
.B(n_412),
.Y(n_430)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_294),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_295),
.C(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_289),
.Y(n_416)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_292),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_322),
.B(n_332),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_313),
.B(n_321),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_319),
.A2(n_358),
.B(n_362),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_330),
.Y(n_332)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_336),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_356),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_345),
.B2(n_346),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_345),
.C(n_356),
.Y(n_376)
);

INVx3_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_349),
.A2(n_366),
.A3(n_368),
.B1(n_369),
.B2(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_352),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_411),
.Y(n_410)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_365),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_370),
.B(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_376),
.B(n_377),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_382),
.B2(n_396),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_381),
.C(n_396),
.Y(n_399)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_382),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_389),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_390),
.C(n_391),
.Y(n_424)
);

INVx8_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_399),
.B(n_400),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_427),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_413),
.B2(n_414),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_413),
.Y(n_471)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_424),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_425),
.C(n_427),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_432),
.B2(n_437),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_433),
.C(n_435),
.Y(n_484)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_432),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_461),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_440),
.A2(n_461),
.B(n_495),
.C(n_498),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_458),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_441),
.B(n_458),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.C(n_446),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_442),
.B(n_444),
.CI(n_446),
.CON(n_474),
.SN(n_474)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_453),
.C(n_456),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_450),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_453),
.A2(n_454),
.B1(n_456),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_456),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_474),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.C(n_468),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.C(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_472),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_474),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_485),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.C(n_484),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_491),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_490),
.Y(n_496)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx13_ASAP7_75t_L g504 ( 
.A(n_501),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_505),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);


endmodule