module fake_jpeg_2558_n_150 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_5),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_15),
.B1(n_29),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_42),
.B1(n_24),
.B2(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_23),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_75),
.Y(n_99)
);

CKINVDCx11_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_74),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_52),
.C(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_13),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_22),
.B(n_18),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_21),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_2),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_62),
.C(n_54),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_62),
.CI(n_54),
.CON(n_87),
.SN(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_80),
.C(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_67),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_47),
.B1(n_3),
.B2(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_99),
.B(n_94),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_75),
.B(n_72),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_97),
.C(n_91),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_107),
.C(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_99),
.B1(n_87),
.B2(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_124),
.B1(n_122),
.B2(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_87),
.B1(n_95),
.B2(n_92),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_120),
.B(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_131),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_106),
.B1(n_111),
.B2(n_102),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_70),
.A3(n_79),
.B1(n_92),
.B2(n_102),
.C1(n_78),
.C2(n_75),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_138),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_117),
.C(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_125),
.B1(n_131),
.B2(n_117),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_134),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_73),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_136),
.C(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_141),
.B1(n_140),
.B2(n_68),
.C(n_73),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_143),
.Y(n_150)
);


endmodule