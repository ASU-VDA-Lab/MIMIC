module fake_jpeg_24188_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_33),
.B1(n_20),
.B2(n_24),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_63),
.B1(n_80),
.B2(n_56),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_61),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_59),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_25),
.C(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_81),
.B1(n_25),
.B2(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_22),
.B1(n_17),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_75),
.B1(n_43),
.B2(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_31),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_22),
.B1(n_34),
.B2(n_23),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_47),
.B1(n_44),
.B2(n_34),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_23),
.B1(n_31),
.B2(n_19),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_107),
.B1(n_62),
.B2(n_35),
.Y(n_127)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_85),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_102),
.B1(n_103),
.B2(n_110),
.Y(n_132)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_89),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_40),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_111),
.C(n_21),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_25),
.Y(n_95)
);

FAx1_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_21),
.CI(n_30),
.CON(n_138),
.SN(n_138)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_25),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_99),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_40),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_43),
.C(n_48),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_146),
.B(n_99),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_79),
.CI(n_48),
.CON(n_126),
.SN(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_87),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_137),
.B1(n_142),
.B2(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_143),
.Y(n_163)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_71),
.A3(n_48),
.B1(n_42),
.B2(n_53),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_110),
.Y(n_162)
);

AO22x2_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_54),
.B1(n_52),
.B2(n_42),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_91),
.B1(n_118),
.B2(n_113),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_85),
.A2(n_27),
.B1(n_29),
.B2(n_52),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_21),
.B(n_32),
.C(n_77),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_106),
.B1(n_108),
.B2(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_42),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_0),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_86),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_111),
.C(n_90),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_185),
.C(n_146),
.Y(n_202)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_160),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_170),
.B(n_173),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_100),
.A3(n_89),
.B1(n_104),
.B2(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_83),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_171),
.B1(n_183),
.B2(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_91),
.B1(n_114),
.B2(n_88),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_178),
.B1(n_179),
.B2(n_140),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_103),
.B1(n_73),
.B2(n_77),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_30),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_94),
.B(n_30),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_30),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_115),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_26),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_181),
.B(n_184),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_11),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_105),
.B1(n_26),
.B2(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_122),
.C(n_126),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_2),
.B(n_3),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_138),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_215),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_168),
.B(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_199),
.B1(n_209),
.B2(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_157),
.A2(n_126),
.B1(n_123),
.B2(n_146),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_205),
.C(n_206),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_123),
.C(n_150),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_115),
.C(n_147),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_145),
.B(n_147),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_172),
.B(n_160),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_151),
.B(n_26),
.C(n_15),
.D(n_13),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.C(n_178),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_130),
.C(n_145),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_218),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_2),
.B(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_2),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_182),
.B1(n_156),
.B2(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_241),
.B1(n_236),
.B2(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_192),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_227),
.B(n_245),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_235),
.B1(n_237),
.B2(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_205),
.C(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_231),
.C(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_166),
.B1(n_154),
.B2(n_171),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_188),
.B1(n_216),
.B2(n_193),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_158),
.C(n_166),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_241),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_169),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_234),
.B1(n_235),
.B2(n_243),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_164),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_199),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_213),
.B(n_153),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_253),
.C(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_229),
.C(n_232),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_228),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_270),
.B1(n_240),
.B2(n_221),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_210),
.C(n_189),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_210),
.C(n_211),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_247),
.C(n_227),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_239),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_188),
.B1(n_213),
.B2(n_203),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_203),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_226),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_245),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_230),
.A2(n_164),
.B1(n_6),
.B2(n_7),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_246),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

BUFx12_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_220),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_225),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_283),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_238),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_258),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_287),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_251),
.B(n_256),
.C(n_261),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_295),
.B(n_305),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_244),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_269),
.B1(n_264),
.B2(n_253),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_294),
.A2(n_297),
.B1(n_304),
.B2(n_290),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_277),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_270),
.B1(n_251),
.B2(n_252),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_244),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_286),
.Y(n_313)
);

OAI322xp33_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_255),
.A3(n_259),
.B1(n_251),
.B2(n_252),
.C1(n_262),
.C2(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_273),
.C(n_276),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_273),
.C(n_276),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_312),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_274),
.C(n_279),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_272),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_278),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_317),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_282),
.B(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_294),
.C(n_290),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_291),
.B1(n_8),
.B2(n_9),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_5),
.C(n_6),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_12),
.C(n_15),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_327),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_324),
.C(n_327),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_297),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_325),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_306),
.C(n_307),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_331),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_318),
.B1(n_310),
.B2(n_316),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_332),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_311),
.C(n_302),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_322),
.B(n_12),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_12),
.B(n_8),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_333),
.C(n_10),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_337),
.B(n_336),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_329),
.C(n_331),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_340),
.B(n_8),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_10),
.Y(n_345)
);


endmodule