module fake_jpeg_14717_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_17),
.B1(n_31),
.B2(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_51),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_24),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_72),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_40),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_81),
.B1(n_22),
.B2(n_21),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_85),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_84),
.Y(n_104)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_22),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_56),
.Y(n_90)
);

NOR2x1_ASAP7_75t_R g116 ( 
.A(n_90),
.B(n_21),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_56),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_95),
.C(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_65),
.B1(n_55),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_103),
.B1(n_79),
.B2(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_67),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_50),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_46),
.B1(n_57),
.B2(n_63),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_78),
.B1(n_80),
.B2(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_38),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_68),
.Y(n_120)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_1),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_133),
.B1(n_134),
.B2(n_109),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_106),
.B(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_68),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_96),
.B1(n_103),
.B2(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_79),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_20),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_30),
.B1(n_28),
.B2(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_107),
.B1(n_28),
.B2(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_30),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_106),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_133),
.B1(n_118),
.B2(n_135),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_141),
.B(n_151),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_112),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_148),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_97),
.C(n_95),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_136),
.C(n_124),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_97),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_149),
.B(n_162),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_154),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_99),
.B(n_111),
.C(n_104),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_129),
.B1(n_158),
.B2(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_28),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_20),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_1),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_2),
.B(n_3),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_2),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_161),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_174),
.B1(n_185),
.B2(n_2),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_179),
.C(n_182),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_130),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_183),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_157),
.B(n_139),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_147),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_116),
.B(n_130),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_176),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_115),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_132),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_150),
.B1(n_154),
.B2(n_148),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_146),
.C(n_144),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_196),
.C(n_197),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_159),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_158),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_199),
.B1(n_204),
.B2(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_146),
.C(n_152),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_152),
.C(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_193),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_178),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_182),
.C(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_214),
.C(n_4),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_185),
.B1(n_177),
.B2(n_164),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_217),
.B1(n_221),
.B2(n_6),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_174),
.B1(n_171),
.B2(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_171),
.B1(n_173),
.B2(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_200),
.CI(n_203),
.CON(n_224),
.SN(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_191),
.B(n_188),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_220),
.B(n_209),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_208),
.C(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_229),
.C(n_234),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_6),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_8),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_220),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_227),
.CI(n_209),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_228),
.C(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_9),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_230),
.B(n_224),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_226),
.B(n_238),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_252),
.B(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_10),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_235),
.B(n_242),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_258),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_236),
.A3(n_239),
.B1(n_224),
.B2(n_13),
.C1(n_9),
.C2(n_11),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_11),
.B(n_13),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_259),
.B(n_14),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_256),
.C(n_261),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_265),
.B(n_14),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_264),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_14),
.Y(n_270)
);


endmodule