module fake_jpeg_31237_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_52),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_34),
.B1(n_39),
.B2(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_64),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_2),
.C(n_3),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_35),
.B1(n_42),
.B2(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_16),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_55),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_4),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_19),
.B(n_6),
.C(n_7),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_4),
.C(n_8),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_92),
.B1(n_10),
.B2(n_11),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_15),
.B1(n_22),
.B2(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_83),
.C(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_103),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_85),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_102),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_105),
.B1(n_83),
.B2(n_100),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_98),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_86),
.Y(n_110)
);


endmodule