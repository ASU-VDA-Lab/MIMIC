module fake_jpeg_11535_n_443 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_443);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_66),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_20),
.B1(n_42),
.B2(n_49),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_39),
.B1(n_37),
.B2(n_24),
.Y(n_124)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_74),
.B(n_77),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_15),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_26),
.B(n_15),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_26),
.B(n_1),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_30),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_107),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_1),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_50),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_37),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_57),
.A2(n_20),
.B1(n_50),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_116),
.A2(n_124),
.B1(n_136),
.B2(n_160),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_120),
.B(n_113),
.C(n_114),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_62),
.A2(n_50),
.B1(n_18),
.B2(n_40),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_121),
.A2(n_167),
.B(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_125),
.B(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_74),
.B(n_51),
.Y(n_130)
);

NAND2x1p5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_36),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_134),
.B(n_90),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_32),
.B1(n_51),
.B2(n_46),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_139),
.B(n_143),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_77),
.Y(n_143)
);

OA22x2_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_40),
.B1(n_39),
.B2(n_24),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_116),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_46),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_44),
.B1(n_32),
.B2(n_22),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_176),
.B1(n_76),
.B2(n_4),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_59),
.A2(n_55),
.B1(n_31),
.B2(n_27),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_60),
.A2(n_40),
.B1(n_55),
.B2(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_44),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_27),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_23),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_69),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_110),
.A2(n_40),
.B1(n_25),
.B2(n_21),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_180),
.B(n_181),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_85),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_21),
.B(n_92),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_182),
.A2(n_153),
.B(n_128),
.Y(n_257)
);

BUFx6f_ASAP7_75t_SL g183 ( 
.A(n_158),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_127),
.A2(n_99),
.B1(n_70),
.B2(n_72),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_177),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_191),
.B(n_202),
.Y(n_270)
);

OAI21x1_ASAP7_75t_SL g254 ( 
.A1(n_192),
.A2(n_234),
.B(n_153),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_193),
.A2(n_205),
.B(n_217),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_118),
.B(n_2),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_2),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_201),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_198),
.B(n_206),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_81),
.C(n_78),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_199),
.B(n_210),
.C(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_3),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_203),
.B(n_207),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_3),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_131),
.B(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_213),
.Y(n_280)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_214),
.B(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_160),
.B1(n_178),
.B2(n_121),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_223),
.B1(n_220),
.B2(n_212),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_5),
.C(n_7),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_220),
.Y(n_253)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_222),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_167),
.A2(n_8),
.B1(n_10),
.B2(n_144),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_227),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_147),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_225),
.B(n_231),
.Y(n_271)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_228),
.A2(n_229),
.B1(n_233),
.B2(n_191),
.Y(n_274)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_140),
.A2(n_8),
.B1(n_10),
.B2(n_179),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_236),
.B1(n_173),
.B2(n_166),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_8),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_235),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_127),
.A2(n_161),
.B1(n_117),
.B2(n_155),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_119),
.B(n_123),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_140),
.A2(n_179),
.B1(n_146),
.B2(n_126),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_141),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_157),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_126),
.B1(n_146),
.B2(n_173),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_239),
.A2(n_260),
.B1(n_277),
.B2(n_282),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_141),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_244),
.B(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_250),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_170),
.B1(n_115),
.B2(n_129),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_188),
.B1(n_182),
.B2(n_201),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_133),
.B1(n_157),
.B2(n_117),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_254),
.A2(n_257),
.B(n_229),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_255),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_157),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_267),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_210),
.A2(n_128),
.B(n_209),
.C(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_128),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_219),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_273),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_199),
.A2(n_208),
.B1(n_223),
.B2(n_196),
.Y(n_272)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_194),
.B1(n_183),
.B2(n_235),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_202),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_234),
.B1(n_203),
.B2(n_186),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_221),
.A2(n_224),
.B1(n_211),
.B2(n_232),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_185),
.B(n_213),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_283),
.A2(n_293),
.B(n_304),
.Y(n_318)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_206),
.B1(n_228),
.B2(n_189),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_287),
.B1(n_294),
.B2(n_307),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_247),
.A2(n_218),
.B1(n_184),
.B2(n_187),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_244),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_258),
.B(n_227),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_290),
.B(n_299),
.Y(n_339)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_241),
.Y(n_292)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_266),
.A2(n_254),
.B1(n_240),
.B2(n_272),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_264),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_278),
.C(n_252),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_250),
.B1(n_253),
.B2(n_266),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_296),
.A2(n_279),
.B1(n_246),
.B2(n_243),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_303),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_238),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_275),
.B(n_259),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_256),
.A2(n_264),
.B(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_276),
.B1(n_262),
.B2(n_253),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_308),
.B(n_315),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_255),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_314),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_310),
.A2(n_312),
.B1(n_263),
.B2(n_268),
.Y(n_334)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_276),
.A2(n_238),
.B1(n_244),
.B2(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_281),
.B1(n_261),
.B2(n_242),
.Y(n_340)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_271),
.B(n_252),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_328),
.Y(n_358)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_244),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_333),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_344),
.B1(n_314),
.B2(n_283),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_338),
.C(n_309),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_265),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_335),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_292),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_265),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_274),
.B1(n_245),
.B2(n_251),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_343),
.B1(n_300),
.B2(n_301),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_286),
.C(n_306),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_300),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_308),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_341),
.Y(n_351)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_342),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_243),
.B1(n_261),
.B2(n_268),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_263),
.B1(n_282),
.B2(n_287),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_345),
.A2(n_315),
.B1(n_290),
.B2(n_303),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_335),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_346),
.B(n_326),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_322),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_306),
.B(n_293),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_331),
.B(n_330),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_318),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_354),
.C(n_356),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_328),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_331),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_341),
.B(n_299),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_353),
.B(n_325),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_286),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_311),
.C(n_306),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_361),
.C(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_364),
.B1(n_340),
.B2(n_324),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_311),
.C(n_306),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_307),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_336),
.B1(n_324),
.B2(n_326),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_322),
.A2(n_305),
.B1(n_301),
.B2(n_288),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_321),
.B1(n_333),
.B2(n_284),
.Y(n_384)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_359),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_358),
.B(n_319),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_374),
.A2(n_385),
.B1(n_351),
.B2(n_358),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_339),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_378),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_347),
.A2(n_325),
.B(n_337),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_377),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_351),
.A2(n_337),
.B(n_288),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_361),
.B(n_313),
.CI(n_339),
.CON(n_380),
.SN(n_380)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_382),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_384),
.Y(n_391)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_352),
.A2(n_342),
.B1(n_310),
.B2(n_332),
.Y(n_385)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_383),
.C(n_350),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_393),
.C(n_396),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_354),
.C(n_357),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_349),
.C(n_363),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_362),
.B1(n_360),
.B2(n_366),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_364),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_356),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_371),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_372),
.B1(n_398),
.B2(n_390),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_402),
.B(n_404),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_406),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_382),
.B1(n_373),
.B2(n_368),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_376),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_405),
.B(n_410),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_369),
.B1(n_370),
.B2(n_375),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_387),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_381),
.C(n_384),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_409),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_385),
.C(n_348),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_380),
.C(n_377),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_400),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_387),
.B(n_394),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_407),
.C(n_401),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_415),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_386),
.Y(n_415)
);

NOR3xp33_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_380),
.C(n_367),
.Y(n_418)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_418),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_367),
.C(n_355),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_401),
.B(n_411),
.Y(n_423)
);

AOI21xp33_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_414),
.B(n_355),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_421),
.A2(n_397),
.B1(n_406),
.B2(n_394),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_426),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_419),
.A2(n_417),
.B(n_420),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_424),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_415),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_428),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_422),
.B1(n_426),
.B2(n_342),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_432),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_433),
.A2(n_310),
.B(n_332),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_435),
.B(n_436),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_430),
.C(n_431),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_310),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_438),
.B(n_437),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_434),
.C(n_439),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_310),
.B(n_332),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_263),
.Y(n_443)
);


endmodule