module fake_jpeg_4320_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.Y(n_15)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_20),
.A3(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_19),
.B1(n_8),
.B2(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_2),
.CI(n_3),
.CON(n_20),
.SN(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_9),
.B(n_13),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_8),
.A3(n_11),
.B1(n_12),
.B2(n_9),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_15),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_30),
.B1(n_25),
.B2(n_3),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_20),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_25),
.B(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_18),
.B1(n_8),
.B2(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_41)
);

OAI31xp33_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_37),
.A3(n_41),
.B(n_2),
.Y(n_43)
);

AOI22x1_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_4),
.B1(n_42),
.B2(n_24),
.Y(n_44)
);


endmodule