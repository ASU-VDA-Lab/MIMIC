module fake_aes_5126_n_585 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_585);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_585;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_305;
wire n_100;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_70), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_30), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_38), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_72), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_68), .Y(n_89) );
INVx2_ASAP7_75t_SL g90 ( .A(n_36), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_50), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_77), .Y(n_92) );
INVxp33_ASAP7_75t_L g93 ( .A(n_34), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_10), .Y(n_96) );
BUFx10_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_18), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_25), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_69), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_80), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_12), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_10), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_81), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_63), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_74), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_59), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_58), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_64), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_5), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_43), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_41), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_99), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
NOR2xp33_ASAP7_75t_SL g128 ( .A(n_99), .B(n_29), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_106), .B(n_101), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_96), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_131) );
CKINVDCx8_ASAP7_75t_R g132 ( .A(n_112), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_106), .B(n_0), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_97), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_95), .B(n_1), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_109), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_98), .Y(n_146) );
INVx5_ASAP7_75t_L g147 ( .A(n_142), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_139), .B(n_97), .Y(n_148) );
OR2x6_ASAP7_75t_L g149 ( .A(n_139), .B(n_110), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_138), .B(n_90), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_138), .B(n_112), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_135), .A2(n_105), .B1(n_115), .B2(n_104), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_135), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_138), .B(n_89), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_138), .B(n_93), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_144), .B(n_90), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_144), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_144), .B(n_104), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_144), .Y(n_163) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_128), .B(n_94), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_123), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_124), .B(n_83), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_124), .B(n_105), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_146), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_133), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_143), .B(n_115), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_125), .B(n_94), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_143), .B(n_102), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_170), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_155), .B(n_132), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_161), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_156), .A2(n_134), .B(n_126), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_149), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_155), .B(n_132), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_168), .B(n_160), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g185 ( .A1(n_149), .A2(n_131), .B1(n_118), .B2(n_130), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_149), .B(n_130), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_156), .B(n_125), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_173), .B(n_102), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_148), .B(n_126), .Y(n_200) );
BUFx8_ASAP7_75t_L g201 ( .A(n_174), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_148), .B(n_127), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_173), .B(n_127), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_150), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_150), .B(n_131), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_166), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_150), .B(n_134), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
AND2x6_ASAP7_75t_L g211 ( .A(n_173), .B(n_116), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_174), .B1(n_172), .B2(n_164), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_184), .A2(n_159), .B(n_163), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_202), .A2(n_154), .B(n_172), .C(n_151), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_178), .A2(n_159), .B(n_163), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_210), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_210), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_206), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_186), .A2(n_164), .B1(n_152), .B2(n_157), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_178), .A2(n_164), .B(n_167), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_200), .B(n_174), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_192), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_205), .B1(n_185), .B2(n_211), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_181), .A2(n_118), .B1(n_141), .B2(n_140), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_181), .B(n_174), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_203), .A2(n_141), .B(n_140), .C(n_136), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_209), .B(n_174), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_209), .B(n_136), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_179), .A2(n_120), .B(n_116), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_205), .A2(n_137), .B1(n_145), .B2(n_117), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_200), .B(n_137), .Y(n_234) );
BUFx8_ASAP7_75t_SL g235 ( .A(n_175), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
OR2x6_ASAP7_75t_SL g238 ( .A(n_175), .B(n_117), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_196), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_198), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
AOI21xp33_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_114), .B(n_86), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_209), .B(n_145), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_195), .B(n_111), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_199), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_200), .B(n_205), .Y(n_247) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_179), .B(n_189), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_213), .A2(n_215), .B(n_246), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_218), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_212), .A2(n_224), .B1(n_246), .B2(n_225), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_223), .A2(n_187), .B(n_180), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_235), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_225), .A2(n_187), .B(n_189), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_247), .B(n_200), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_235), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_247), .B(n_187), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_228), .B(n_207), .C(n_204), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_239), .B(n_190), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_241), .A2(n_190), .B(n_199), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_220), .A2(n_211), .B1(n_198), .B2(n_207), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_219), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_233), .A2(n_204), .B(n_188), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_237), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_237), .B(n_201), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_226), .A2(n_85), .B(n_122), .Y(n_272) );
BUFx2_ASAP7_75t_R g273 ( .A(n_238), .Y(n_273) );
INVx8_ASAP7_75t_L g274 ( .A(n_227), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_214), .A2(n_231), .B(n_208), .C(n_233), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_232), .A2(n_198), .B1(n_211), .B2(n_234), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_230), .B(n_208), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_244), .B(n_87), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_258), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_265), .A2(n_222), .B(n_229), .C(n_233), .Y(n_280) );
AO31x2_ASAP7_75t_L g281 ( .A1(n_252), .A2(n_188), .A3(n_183), .B(n_191), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_251), .B(n_234), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_251), .B(n_227), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_249), .A2(n_245), .B(n_191), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_242), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_252), .A2(n_176), .B1(n_182), .B2(n_243), .C(n_238), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_261), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_261), .B(n_227), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_260), .B(n_197), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
AOI222xp33_ASAP7_75t_L g291 ( .A1(n_257), .A2(n_236), .B1(n_201), .B2(n_198), .C1(n_211), .C2(n_195), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_250), .A2(n_240), .B1(n_236), .B2(n_245), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_269), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_263), .A2(n_245), .B(n_197), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_260), .B(n_217), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_265), .A2(n_211), .B1(n_198), .B2(n_217), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_255), .Y(n_300) );
AO21x1_ASAP7_75t_SL g301 ( .A1(n_269), .A2(n_113), .B(n_103), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_260), .B(n_217), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_287), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_289), .B(n_267), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_267), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_296), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_278), .A2(n_248), .B(n_268), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_302), .B(n_267), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_293), .B(n_257), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_279), .B(n_257), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_297), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_290), .Y(n_318) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_286), .A2(n_273), .B(n_276), .C(n_271), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_290), .B(n_256), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_299), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_298), .A2(n_273), .B1(n_276), .B2(n_263), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_282), .B(n_285), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_320), .B(n_284), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_320), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_326), .A2(n_282), .B1(n_285), .B2(n_283), .C(n_288), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_306), .B(n_302), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_319), .B(n_254), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_311), .B(n_259), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_306), .B(n_302), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_311), .B(n_274), .Y(n_343) );
NAND2xp33_ASAP7_75t_R g344 ( .A(n_310), .B(n_2), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_307), .B(n_300), .Y(n_346) );
AOI211x1_ASAP7_75t_SL g347 ( .A1(n_325), .A2(n_271), .B(n_121), .C(n_275), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_321), .B(n_281), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_305), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_281), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_321), .B(n_281), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_328), .B(n_309), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_309), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_348), .B(n_309), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_352), .B(n_309), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_327), .A2(n_292), .B(n_294), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_332), .B(n_315), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_348), .B(n_281), .Y(n_365) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_331), .B(n_322), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_355), .B(n_315), .Y(n_367) );
NAND5xp2_ASAP7_75t_L g368 ( .A(n_336), .B(n_291), .C(n_316), .D(n_280), .E(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_356), .B(n_281), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_327), .B(n_317), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_330), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_333), .B(n_317), .Y(n_374) );
NAND4xp75_ASAP7_75t_SL g375 ( .A(n_344), .B(n_301), .C(n_291), .D(n_316), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_356), .B(n_281), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_349), .B(n_318), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_341), .B(n_3), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_334), .B(n_314), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_349), .B(n_318), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_338), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_323), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_323), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_338), .B(n_322), .Y(n_388) );
AND3x1_ASAP7_75t_L g389 ( .A(n_329), .B(n_301), .C(n_324), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_339), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_327), .B(n_323), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_340), .B(n_324), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_352), .B(n_278), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g397 ( .A(n_350), .B(n_278), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_351), .B(n_278), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_351), .B(n_310), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_335), .B(n_272), .Y(n_400) );
AO22x1_ASAP7_75t_L g401 ( .A1(n_337), .A2(n_300), .B1(n_302), .B2(n_270), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_353), .B(n_248), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_362), .B(n_354), .Y(n_404) );
NOR2x2_ASAP7_75t_L g405 ( .A(n_389), .B(n_121), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_361), .B(n_372), .Y(n_406) );
INVx5_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_361), .B(n_337), .Y(n_408) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_375), .B(n_354), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_346), .B1(n_343), .B2(n_342), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_372), .B(n_350), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_365), .B(n_350), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_372), .B(n_350), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_381), .B(n_368), .Y(n_414) );
NOR3xp33_ASAP7_75t_SL g415 ( .A(n_397), .B(n_108), .C(n_107), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_372), .B(n_284), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_399), .B(n_346), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_399), .B(n_346), .Y(n_418) );
NOR3xp33_ASAP7_75t_SL g419 ( .A(n_400), .B(n_100), .C(n_288), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_365), .B(n_347), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_369), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_370), .B(n_248), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_359), .B(n_119), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_359), .B(n_119), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_358), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_360), .B(n_391), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_373), .B(n_272), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_362), .B(n_295), .Y(n_430) );
OR2x6_ASAP7_75t_L g431 ( .A(n_366), .B(n_300), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_376), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_360), .B(n_119), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_382), .B(n_3), .Y(n_434) );
NAND2x1_ASAP7_75t_L g435 ( .A(n_378), .B(n_391), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_370), .B(n_272), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_379), .B(n_272), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_379), .B(n_119), .Y(n_438) );
OR2x6_ASAP7_75t_L g439 ( .A(n_366), .B(n_300), .Y(n_439) );
NOR2x1p5_ASAP7_75t_SL g440 ( .A(n_394), .B(n_268), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_378), .B(n_268), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_380), .B(n_4), .Y(n_442) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_358), .B(n_283), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_376), .B(n_142), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_358), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_377), .Y(n_446) );
AND2x4_ASAP7_75t_SL g447 ( .A(n_380), .B(n_270), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_377), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_383), .B(n_5), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_383), .B(n_6), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_390), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_392), .B(n_142), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
OAI21xp33_ASAP7_75t_SL g457 ( .A1(n_378), .A2(n_256), .B(n_264), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_392), .B(n_142), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_410), .A2(n_394), .B1(n_363), .B2(n_393), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_395), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_414), .A2(n_410), .B1(n_419), .B2(n_409), .Y(n_461) );
OAI21xp33_ASAP7_75t_SL g462 ( .A1(n_431), .A2(n_388), .B(n_374), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_415), .A2(n_396), .B(n_364), .C(n_367), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_427), .B(n_395), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_431), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_408), .B(n_386), .Y(n_470) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_438), .A2(n_396), .B(n_403), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_456), .B(n_387), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_445), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_411), .B(n_387), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_434), .A2(n_401), .B1(n_403), .B2(n_398), .Y(n_475) );
AOI32xp33_ASAP7_75t_L g476 ( .A1(n_442), .A2(n_398), .A3(n_402), .B1(n_371), .B2(n_384), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_438), .B(n_402), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_445), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_413), .B(n_384), .Y(n_480) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_431), .A2(n_384), .B1(n_371), .B2(n_401), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
OAI21xp33_ASAP7_75t_SL g483 ( .A1(n_439), .A2(n_371), .B(n_256), .Y(n_483) );
OAI322xp33_ASAP7_75t_L g484 ( .A1(n_436), .A2(n_142), .A3(n_9), .B1(n_11), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_SL g485 ( .A1(n_423), .A2(n_277), .B(n_9), .C(n_11), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_412), .B(n_7), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g487 ( .A1(n_457), .A2(n_255), .B(n_262), .C(n_253), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_451), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_439), .B(n_255), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_420), .A2(n_277), .B(n_262), .C(n_14), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_449), .B(n_7), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_450), .Y(n_494) );
AOI221x1_ASAP7_75t_SL g495 ( .A1(n_436), .A2(n_13), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_437), .A2(n_198), .B1(n_211), .B2(n_274), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_437), .A2(n_274), .B1(n_264), .B2(n_249), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_412), .B(n_16), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_420), .A2(n_274), .B1(n_264), .B2(n_249), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_439), .A2(n_274), .B1(n_217), .B2(n_216), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_440), .A2(n_169), .B(n_253), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_424), .B(n_433), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_435), .A2(n_274), .B(n_253), .C(n_19), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_417), .B(n_17), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_418), .B(n_18), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_422), .B(n_19), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_462), .A2(n_443), .B(n_422), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_466), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_469), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_483), .A2(n_416), .B(n_407), .Y(n_512) );
OAI22xp33_ASAP7_75t_SL g513 ( .A1(n_492), .A2(n_407), .B1(n_405), .B2(n_416), .Y(n_513) );
OA22x2_ASAP7_75t_L g514 ( .A1(n_461), .A2(n_426), .B1(n_454), .B2(n_453), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_478), .Y(n_516) );
XNOR2xp5_ASAP7_75t_L g517 ( .A(n_504), .B(n_430), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_494), .B(n_429), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_495), .A2(n_407), .B1(n_404), .B2(n_444), .C(n_455), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_482), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_488), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_493), .Y(n_523) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_506), .A2(n_458), .B1(n_455), .B2(n_444), .C(n_441), .Y(n_524) );
AOI21xp33_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_458), .B(n_441), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_480), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_407), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_473), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_476), .B(n_20), .Y(n_531) );
NAND4xp25_ASAP7_75t_SL g532 ( .A(n_475), .B(n_21), .C(n_22), .D(n_23), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_470), .B(n_468), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_485), .A2(n_26), .B(n_27), .C(n_32), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_479), .B(n_33), .Y(n_535) );
AOI322xp5_ASAP7_75t_L g536 ( .A1(n_491), .A2(n_217), .A3(n_216), .B1(n_169), .B2(n_40), .C1(n_44), .C2(n_45), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_459), .A2(n_216), .B1(n_169), .B2(n_147), .Y(n_538) );
AOI21xp33_ASAP7_75t_L g539 ( .A1(n_514), .A2(n_486), .B(n_498), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_514), .A2(n_503), .B(n_481), .Y(n_540) );
NAND2x2_ASAP7_75t_L g541 ( .A(n_531), .B(n_502), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_518), .B(n_471), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_534), .A2(n_464), .B(n_484), .C(n_505), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_518), .Y(n_544) );
AOI21xp33_ASAP7_75t_SL g545 ( .A1(n_513), .A2(n_500), .B(n_495), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_520), .Y(n_546) );
AOI211xp5_ASAP7_75t_L g547 ( .A1(n_525), .A2(n_484), .B(n_479), .C(n_487), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_517), .A2(n_489), .B1(n_497), .B2(n_499), .Y(n_548) );
AOI322xp5_ASAP7_75t_L g549 ( .A1(n_530), .A2(n_460), .A3(n_496), .B1(n_501), .B2(n_216), .C1(n_169), .C2(n_51), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_511), .B(n_35), .Y(n_550) );
AO221x1_ASAP7_75t_L g551 ( .A1(n_511), .A2(n_216), .B1(n_169), .B2(n_47), .C(n_49), .Y(n_551) );
NOR2xp33_ASAP7_75t_R g552 ( .A(n_532), .B(n_37), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_537), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_517), .B(n_39), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_535), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_508), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_544), .B(n_510), .Y(n_558) );
AOI221x1_ASAP7_75t_L g559 ( .A1(n_548), .A2(n_511), .B1(n_522), .B2(n_512), .C(n_507), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_554), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_539), .A2(n_519), .B1(n_523), .B2(n_515), .C(n_516), .Y(n_561) );
OAI211xp5_ASAP7_75t_L g562 ( .A1(n_545), .A2(n_538), .B(n_524), .C(n_536), .Y(n_562) );
AO22x2_ASAP7_75t_L g563 ( .A1(n_540), .A2(n_529), .B1(n_528), .B2(n_522), .Y(n_563) );
AOI211xp5_ASAP7_75t_L g564 ( .A1(n_543), .A2(n_522), .B(n_529), .C(n_528), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_547), .B(n_535), .C(n_527), .D(n_521), .Y(n_565) );
OAI221xp5_ASAP7_75t_SL g566 ( .A1(n_549), .A2(n_527), .B1(n_533), .B2(n_509), .C(n_526), .Y(n_566) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_555), .A2(n_533), .B(n_526), .C(n_169), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_541), .A2(n_147), .B1(n_53), .B2(n_54), .Y(n_568) );
AND3x4_ASAP7_75t_L g569 ( .A(n_559), .B(n_550), .C(n_552), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_564), .B(n_550), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_560), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_558), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_565), .B(n_542), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g575 ( .A1(n_574), .A2(n_566), .B1(n_568), .B2(n_563), .C1(n_556), .C2(n_561), .Y(n_575) );
AOI222xp33_ASAP7_75t_L g576 ( .A1(n_571), .A2(n_562), .B1(n_557), .B2(n_553), .C1(n_546), .C2(n_551), .Y(n_576) );
XOR2xp5_ASAP7_75t_L g577 ( .A(n_573), .B(n_567), .Y(n_577) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_576), .B(n_572), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_577), .A2(n_569), .B1(n_573), .B2(n_570), .Y(n_579) );
AOI22xp5_ASAP7_75t_SL g580 ( .A1(n_579), .A2(n_575), .B1(n_55), .B2(n_56), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_578), .Y(n_581) );
OAI311xp33_ASAP7_75t_L g582 ( .A1(n_581), .A2(n_52), .A3(n_57), .B1(n_61), .C1(n_65), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_582), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_580), .A3(n_67), .B1(n_71), .B2(n_76), .C1(n_78), .C2(n_66), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_584), .A2(n_147), .B(n_579), .C(n_581), .Y(n_585) );
endmodule