module real_jpeg_15441_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_413),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_0),
.B(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_2),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_2),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_3),
.Y(n_260)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_5),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_5),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_6),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_6),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_6),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_6),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

AND2x4_ASAP7_75t_SL g259 ( 
.A(n_6),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_9),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_23),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_42),
.Y(n_41)
);

NAND2x1p5_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_52),
.Y(n_51)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_10),
.B(n_92),
.Y(n_91)
);

AND2x4_ASAP7_75t_SL g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_10),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_11),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_37),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_12),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_12),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_13),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_97),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_58),
.B(n_96),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_17),
.B(n_58),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.C(n_39),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_19),
.A2(n_20),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_21),
.A2(n_33),
.B1(n_41),
.B2(n_89),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_41),
.B1(n_45),
.B2(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_22),
.B(n_138),
.C(n_142),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_22),
.A2(n_88),
.B(n_93),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_22),
.A2(n_45),
.B1(n_138),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_22),
.A2(n_45),
.B1(n_127),
.B2(n_164),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_25),
.A2(n_26),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_30),
.C(n_45),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_41),
.Y(n_93)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_30),
.A2(n_34),
.B1(n_51),
.B2(n_55),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_30),
.A2(n_34),
.B1(n_64),
.B2(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_30),
.B(n_177),
.C(n_185),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_30),
.B(n_144),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_30),
.B(n_64),
.C(n_131),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_30),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_30),
.B(n_142),
.C(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_30),
.A2(n_34),
.B1(n_185),
.B2(n_372),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_32),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_34),
.B(n_136),
.C(n_144),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.C(n_45),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_41),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_41),
.B(n_90),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_41),
.A2(n_259),
.B(n_275),
.C(n_277),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_41),
.B(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_41),
.A2(n_89),
.B1(n_259),
.B2(n_261),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_41),
.B(n_64),
.C(n_91),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_44),
.A2(n_110),
.B(n_117),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_44),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_45),
.B(n_127),
.C(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_55),
.B1(n_105),
.B2(n_114),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_110),
.C(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_51),
.A2(n_55),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_51),
.A2(n_55),
.B1(n_298),
.B2(n_302),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_51),
.B(n_113),
.C(n_298),
.Y(n_334)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_55),
.B(n_142),
.C(n_156),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.C(n_81),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_59),
.B(n_62),
.Y(n_225)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_72),
.C(n_77),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.C(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_64),
.A2(n_134),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_64),
.A2(n_134),
.B1(n_210),
.B2(n_211),
.Y(n_329)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_66),
.B(n_123),
.C(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_122),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_66),
.A2(n_90),
.B1(n_91),
.B2(n_122),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_66),
.A2(n_91),
.B(n_237),
.C(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_77),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_72),
.A2(n_86),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_72),
.B(n_90),
.C(n_106),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_72),
.A2(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_72),
.B(n_331),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_128),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_73),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_81),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.C(n_94),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_82),
.A2(n_83),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_87),
.B(n_94),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B(n_93),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_91),
.B1(n_106),
.B2(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_90),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_90),
.B(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_228),
.B(n_405),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_212),
.C(n_223),
.Y(n_99)
);

AND2x4_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_193),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_101),
.B(n_193),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_147),
.C(n_165),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_102),
.B(n_147),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_129),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_130),
.C(n_135),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.C(n_120),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_104),
.B(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_105),
.A2(n_114),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_113),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_110),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_106),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_106),
.A2(n_132),
.B1(n_182),
.B2(n_247),
.Y(n_313)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_117),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_110),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_110),
.A2(n_170),
.B1(n_244),
.B2(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_111),
.Y(n_332)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_113),
.B(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_114),
.A2(n_254),
.B(n_259),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_115),
.B(n_120),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_116),
.Y(n_323)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_117),
.A2(n_171),
.B1(n_255),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_117),
.A2(n_138),
.B1(n_171),
.B2(n_175),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_117),
.B(n_138),
.C(n_311),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_127),
.A2(n_164),
.B1(n_298),
.B2(n_302),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_132),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_136),
.A2(n_137),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_142),
.A2(n_155),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_144),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_178),
.C(n_182),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_152),
.C(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_163),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_164),
.B(n_302),
.C(n_343),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_165),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.C(n_189),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_166),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_173),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_172),
.Y(n_391)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_173),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_176),
.A2(n_189),
.B1(n_190),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_177),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_178),
.A2(n_182),
.B1(n_247),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_178),
.Y(n_353)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_182),
.Y(n_247)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_185),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_196),
.C(n_203),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

XNOR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_201),
.C(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_213),
.A2(n_408),
.B(n_409),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_214),
.B(n_222),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_223),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_224),
.B(n_226),
.Y(n_412)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI321xp33_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_359),
.A3(n_392),
.B1(n_398),
.B2(n_403),
.C(n_404),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_336),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_315),
.B(n_335),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_292),
.B(n_314),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_272),
.B(n_291),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_251),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_243),
.C(n_248),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_237),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_237),
.A2(n_241),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_248),
.B1(n_249),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_244),
.B(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_263),
.C(n_271),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_283),
.B(n_285),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_267),
.A2(n_311),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_281),
.B(n_290),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_278),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_287),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_286),
.B(n_289),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_294),
.Y(n_314)
);

XOR2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_303),
.C(n_304),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

OR2x6_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_309),
.C(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_317),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_320),
.C(n_327),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_324),
.C(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_334),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_330),
.C(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_333),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_338),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_349),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_339),
.B(n_350),
.C(n_358),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_347),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_345),
.C(n_347),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_358),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_356),
.C(n_357),
.Y(n_366)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_379),
.Y(n_359)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_377),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_377),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.C(n_373),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_374),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.C(n_368),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_369),
.B1(n_370),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI31xp67_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_393),
.A3(n_399),
.B(n_402),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_382),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.C(n_388),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_383),
.A2(n_384),
.B1(n_388),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_388),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_394),
.B(n_397),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_410),
.B(n_411),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);


endmodule