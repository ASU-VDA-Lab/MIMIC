module fake_jpeg_28115_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_24),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_15),
.B1(n_37),
.B2(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_44),
.B1(n_49),
.B2(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_15),
.B1(n_22),
.B2(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B1(n_16),
.B2(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_58),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_48),
.C(n_45),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_65),
.C(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_68),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_14),
.B1(n_19),
.B2(n_22),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_30),
.C(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_72),
.B1(n_16),
.B2(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_38),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_81),
.B(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_25),
.B1(n_23),
.B2(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.C(n_10),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_5),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_16),
.C(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_25),
.B(n_16),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_97),
.B(n_71),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_1),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_103),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_8),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_11),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_11),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_65),
.B1(n_77),
.B2(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_112),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_62),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_116),
.B(n_100),
.C(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_67),
.B(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_12),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_102),
.C(n_95),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_133),
.C(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_105),
.Y(n_143)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_117),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_102),
.C(n_87),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_112),
.B(n_110),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_93),
.C(n_97),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_134),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_139),
.B(n_145),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_108),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_106),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_113),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_146),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_114),
.B1(n_109),
.B2(n_89),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_106),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_134),
.C(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_134),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_140),
.B1(n_146),
.B2(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_157),
.B1(n_148),
.B2(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_111),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_148),
.B1(n_152),
.B2(n_130),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_126),
.B(n_92),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_166),
.B(n_118),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_162),
.B(n_165),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_63),
.B1(n_92),
.B2(n_12),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_169),
.B1(n_104),
.B2(n_126),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_171),
.B(n_13),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_171),
.Y(n_173)
);


endmodule