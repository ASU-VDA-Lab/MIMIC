module fake_jpeg_7806_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_20),
.Y(n_81)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_35),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_32),
.B1(n_26),
.B2(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_67),
.B(n_73),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_40),
.C(n_37),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_18),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_38),
.B1(n_22),
.B2(n_26),
.Y(n_100)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_59),
.B1(n_57),
.B2(n_53),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_39),
.Y(n_86)
);

XNOR2x1_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_92),
.B1(n_22),
.B2(n_40),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_38),
.B1(n_45),
.B2(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_93),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_95),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_151)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_108),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_21),
.C(n_27),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_76),
.B(n_33),
.Y(n_128)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_117),
.B1(n_31),
.B2(n_79),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_37),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_27),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_18),
.B1(n_33),
.B2(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_14),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_72),
.B1(n_86),
.B2(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_135),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_103),
.B1(n_116),
.B2(n_106),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_72),
.B1(n_70),
.B2(n_93),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_70),
.B(n_95),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_101),
.B(n_108),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_74),
.B1(n_75),
.B2(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_84),
.B1(n_75),
.B2(n_88),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_24),
.B(n_80),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_147),
.B(n_23),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_105),
.B1(n_100),
.B2(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_80),
.B(n_71),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_101),
.B(n_21),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_12),
.B(n_14),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_24),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_126),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_122),
.C(n_121),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_84),
.B1(n_91),
.B2(n_29),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_91),
.B1(n_29),
.B2(n_30),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_171),
.C(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_174),
.Y(n_200)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_172),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_166),
.B(n_169),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_138),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_115),
.B(n_118),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_178),
.B(n_185),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_123),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_181),
.B(n_191),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_25),
.C(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_188),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_25),
.C(n_28),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_149),
.C(n_21),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_134),
.B(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_196),
.A2(n_212),
.B(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_210),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_202),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_132),
.B1(n_134),
.B2(n_148),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_176),
.B1(n_161),
.B2(n_162),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_132),
.B1(n_152),
.B2(n_141),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_185),
.B1(n_174),
.B2(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_132),
.B1(n_144),
.B2(n_145),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_216),
.C(n_186),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_144),
.B(n_11),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_25),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_219),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_242),
.B1(n_221),
.B2(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_166),
.B1(n_188),
.B2(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_230),
.C(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_243),
.B1(n_221),
.B2(n_220),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_167),
.C(n_170),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_176),
.B1(n_169),
.B2(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_192),
.C(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_165),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_163),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_23),
.Y(n_240)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_29),
.B1(n_30),
.B2(n_19),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_21),
.C(n_28),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_245),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_193),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_27),
.C(n_19),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_226),
.C(n_244),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_206),
.CI(n_212),
.CON(n_252),
.SN(n_252)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_258),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_202),
.B1(n_193),
.B2(n_217),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_259),
.B1(n_265),
.B2(n_267),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_197),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_223),
.A2(n_194),
.B1(n_211),
.B2(n_198),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_198),
.B(n_222),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_0),
.B(n_1),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_195),
.B1(n_214),
.B2(n_30),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_214),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_227),
.A3(n_236),
.B1(n_232),
.B2(n_230),
.C1(n_229),
.C2(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_274),
.C(n_277),
.Y(n_299)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_272),
.B(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_27),
.C(n_19),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_6),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_6),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_5),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_256),
.B(n_8),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_282),
.B1(n_254),
.B2(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_286),
.B(n_291),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_266),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_292),
.C(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_257),
.B1(n_262),
.B2(n_259),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_253),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_256),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_264),
.B1(n_249),
.B2(n_9),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_283),
.B1(n_270),
.B2(n_280),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_14),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_5),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_2),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_3),
.B1(n_4),
.B2(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_11),
.C(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_309),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_1),
.C(n_2),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_4),
.C(n_303),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_2),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_3),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_3),
.C(n_4),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_4),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_290),
.B(n_289),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_317),
.B(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_318),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_290),
.B1(n_296),
.B2(n_3),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_310),
.B(n_316),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_320),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_308),
.C(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_314),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_321),
.B(n_323),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_328),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_313),
.C(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_313),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_325),
.Y(n_335)
);


endmodule