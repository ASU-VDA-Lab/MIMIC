module fake_jpeg_20945_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_20),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_12),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_11),
.C(n_8),
.Y(n_35)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_24),
.B1(n_23),
.B2(n_13),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_11),
.B1(n_10),
.B2(n_27),
.Y(n_39)
);

XOR2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_7),
.C(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_17),
.C(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_15),
.C(n_22),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_29),
.B1(n_7),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_36),
.B1(n_38),
.B2(n_29),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_50),
.B1(n_47),
.B2(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_25),
.C(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.C(n_48),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_52),
.C(n_3),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.A3(n_0),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_36),
.Y(n_58)
);

XNOR2x1_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_4),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVxp33_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_2),
.Y(n_61)
);


endmodule