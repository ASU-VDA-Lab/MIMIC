module fake_jpeg_751_n_696 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_696);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_696;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_59),
.Y(n_181)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_61),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_62),
.Y(n_190)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_81),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_69),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_71),
.B(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_73),
.Y(n_234)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_9),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_85),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_88),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_51),
.B(n_9),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_100),
.B(n_104),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_103),
.B(n_124),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_10),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_120),
.Y(n_192)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_37),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_45),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_26),
.Y(n_131)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_56),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_135),
.B(n_147),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_82),
.A2(n_45),
.B(n_48),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_150),
.B(n_211),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_62),
.A2(n_33),
.B1(n_26),
.B2(n_35),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_159),
.A2(n_165),
.B1(n_183),
.B2(n_200),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_61),
.B(n_43),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_162),
.B(n_90),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_62),
.A2(n_33),
.B1(n_26),
.B2(n_35),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_65),
.A2(n_47),
.B1(n_35),
.B2(n_54),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_166),
.A2(n_85),
.B1(n_80),
.B2(n_75),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_64),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_167),
.B(n_187),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_89),
.A2(n_23),
.B1(n_32),
.B2(n_43),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_168),
.A2(n_199),
.B1(n_214),
.B2(n_217),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_47),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_171),
.B(n_178),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_32),
.B(n_23),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_172),
.A2(n_86),
.B(n_1),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_83),
.B(n_47),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_69),
.A2(n_33),
.B1(n_21),
.B2(n_54),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_111),
.B(n_28),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_58),
.A2(n_54),
.B1(n_21),
.B2(n_38),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_69),
.A2(n_21),
.B1(n_32),
.B2(n_23),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_94),
.B(n_40),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_96),
.Y(n_207)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_94),
.B(n_47),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_107),
.B(n_40),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_40),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_216),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_88),
.A2(n_38),
.B1(n_24),
.B2(n_20),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_91),
.B(n_38),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_109),
.A2(n_24),
.B1(n_20),
.B2(n_52),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_70),
.B(n_24),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_225),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_77),
.B(n_20),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_136),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_84),
.B(n_121),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_128),
.B(n_52),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_105),
.B(n_52),
.Y(n_227)
);

AOI22x1_ASAP7_75t_L g229 ( 
.A1(n_124),
.A2(n_42),
.B1(n_10),
.B2(n_11),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_229),
.A2(n_236),
.B1(n_0),
.B2(n_1),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_117),
.B(n_42),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_66),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_131),
.A2(n_42),
.B1(n_11),
.B2(n_12),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_231),
.A2(n_181),
.B1(n_182),
.B2(n_220),
.Y(n_296)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

HAxp5_ASAP7_75t_SL g236 ( 
.A(n_90),
.B(n_8),
.CON(n_236),
.SN(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_192),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_239),
.B(n_260),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_240),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_168),
.A2(n_211),
.B1(n_130),
.B2(n_110),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_241),
.A2(n_262),
.B1(n_272),
.B2(n_299),
.Y(n_387)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_249),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_250),
.B(n_275),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_200),
.A2(n_125),
.B1(n_122),
.B2(n_113),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_251),
.A2(n_179),
.B1(n_153),
.B2(n_148),
.Y(n_392)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_252),
.Y(n_360)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx4_ASAP7_75t_SL g384 ( 
.A(n_254),
.Y(n_384)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_156),
.Y(n_255)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_197),
.B(n_73),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_259),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_172),
.A2(n_101),
.B1(n_112),
.B2(n_72),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_261),
.A2(n_292),
.B1(n_295),
.B2(n_308),
.Y(n_328)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_264),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_204),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_265),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_266),
.B(n_279),
.Y(n_336)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_269),
.Y(n_386)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_271),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_185),
.A2(n_67),
.B1(n_196),
.B2(n_214),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_171),
.B(n_0),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_274),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_157),
.B(n_12),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_149),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_278),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_193),
.B(n_12),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_146),
.B(n_143),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_280),
.B(n_284),
.Y(n_382)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_234),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_289),
.Y(n_348)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_285),
.Y(n_376)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_173),
.Y(n_286)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_287),
.B(n_298),
.Y(n_359)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_137),
.Y(n_288)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_201),
.B(n_12),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_290),
.Y(n_380)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_137),
.Y(n_291)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_229),
.A2(n_86),
.B1(n_7),
.B2(n_13),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_178),
.B(n_0),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_293),
.Y(n_379)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_202),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_294),
.B(n_297),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_206),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_296),
.A2(n_310),
.B1(n_313),
.B2(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_169),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_184),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_180),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_300),
.Y(n_346)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_184),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_303),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_218),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_302),
.Y(n_385)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_174),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_175),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_307),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_177),
.Y(n_306)
);

INVx11_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_141),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_139),
.A2(n_164),
.B1(n_161),
.B2(n_158),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_138),
.B(n_16),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_322),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_181),
.A2(n_150),
.B1(n_189),
.B2(n_163),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_142),
.Y(n_312)
);

INVx11_ASAP7_75t_L g372 ( 
.A(n_312),
.Y(n_372)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_159),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_154),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_314),
.B(n_319),
.Y(n_378)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_218),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_323),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_142),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_139),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_141),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_140),
.B(n_2),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_321),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_160),
.B(n_2),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_210),
.B(n_16),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_144),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_236),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_215),
.B(n_19),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_148),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_170),
.B1(n_223),
.B2(n_144),
.Y(n_351)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_221),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_300),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_339),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_271),
.A2(n_217),
.B(n_165),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_343),
.A2(n_356),
.B(n_290),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_256),
.A2(n_203),
.B(n_231),
.C(n_152),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_347),
.A2(n_369),
.B(n_254),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_305),
.A2(n_313),
.B1(n_258),
.B2(n_253),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_350),
.A2(n_351),
.B1(n_388),
.B2(n_392),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_262),
.A2(n_170),
.B1(n_223),
.B2(n_209),
.Y(n_353)
);

AOI22x1_ASAP7_75t_L g405 ( 
.A1(n_353),
.A2(n_323),
.B1(n_318),
.B2(n_293),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_256),
.A2(n_188),
.B(n_220),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_248),
.B(n_209),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_381),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_268),
.A2(n_182),
.B(n_152),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_245),
.B(n_152),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_259),
.C(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_243),
.B(n_213),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_311),
.A2(n_284),
.B(n_299),
.C(n_241),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_383),
.A2(n_133),
.B(n_265),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_257),
.A2(n_213),
.B1(n_186),
.B2(n_179),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_320),
.B(n_186),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_321),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_387),
.A2(n_256),
.B1(n_311),
.B2(n_272),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_393),
.A2(n_404),
.B1(n_407),
.B2(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_335),
.Y(n_394)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_396),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_398),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_259),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_387),
.A2(n_311),
.B1(n_295),
.B2(n_308),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_400),
.A2(n_426),
.B1(n_346),
.B2(n_385),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_333),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_403),
.B(n_424),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_363),
.A2(n_383),
.B1(n_357),
.B2(n_381),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_405),
.A2(n_378),
.B1(n_434),
.B2(n_433),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_321),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_413),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_383),
.A2(n_311),
.B1(n_274),
.B2(n_293),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_238),
.C(n_244),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_439),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_330),
.B(n_240),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_409),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_303),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_410),
.Y(n_464)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_274),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

NOR2x1p5_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_267),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_425),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_332),
.A2(n_153),
.B1(n_291),
.B2(n_288),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_419),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_334),
.B(n_316),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_420),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_331),
.B(n_237),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_421),
.B(n_422),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_242),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_343),
.A2(n_270),
.B(n_269),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_423),
.A2(n_430),
.B(n_436),
.Y(n_457)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_329),
.B(n_247),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_382),
.A2(n_307),
.B1(n_255),
.B2(n_249),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_336),
.B(n_301),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_427),
.B(n_429),
.Y(n_476)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_435),
.B1(n_384),
.B2(n_252),
.Y(n_448)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_432),
.Y(n_461)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_433),
.B(n_437),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_328),
.A2(n_317),
.B1(n_312),
.B2(n_263),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_438),
.B1(n_442),
.B2(n_384),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_328),
.A2(n_246),
.B1(n_298),
.B2(n_273),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_375),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_368),
.A2(n_133),
.B1(n_281),
.B2(n_134),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_379),
.B(n_228),
.C(n_134),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_369),
.B(n_228),
.C(n_302),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_356),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_334),
.B(n_306),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_384),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_447),
.A2(n_466),
.B1(n_469),
.B2(n_454),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_448),
.A2(n_418),
.B(n_360),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_439),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_359),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_450),
.B(n_452),
.C(n_483),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_397),
.B(n_359),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g501 ( 
.A1(n_454),
.A2(n_480),
.B1(n_428),
.B2(n_394),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_455),
.B(n_456),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_329),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_353),
.B1(n_351),
.B2(n_378),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_458),
.A2(n_459),
.B1(n_465),
.B2(n_478),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_407),
.A2(n_378),
.B1(n_359),
.B2(n_391),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_404),
.A2(n_382),
.B1(n_389),
.B2(n_339),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_442),
.A2(n_342),
.B1(n_389),
.B2(n_362),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_395),
.B(n_390),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_477),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_395),
.B(n_371),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_431),
.A2(n_380),
.B1(n_362),
.B2(n_371),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_415),
.A2(n_371),
.B1(n_346),
.B2(n_344),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_481),
.A2(n_405),
.B1(n_423),
.B2(n_421),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_399),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_484),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_344),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_385),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_413),
.B(n_355),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_376),
.C(n_373),
.Y(n_515)
);

OAI32xp33_ASAP7_75t_L g487 ( 
.A1(n_463),
.A2(n_415),
.A3(n_440),
.B1(n_403),
.B2(n_430),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_488),
.A2(n_444),
.B1(n_470),
.B2(n_461),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_490),
.B(n_473),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_452),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_492),
.B(n_518),
.C(n_377),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_457),
.A2(n_416),
.B(n_405),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_493),
.A2(n_494),
.B(n_505),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_429),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_451),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_501),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_445),
.A2(n_422),
.B1(n_396),
.B2(n_412),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_496),
.A2(n_510),
.B1(n_472),
.B2(n_486),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_498),
.A2(n_500),
.B1(n_511),
.B2(n_512),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_445),
.A2(n_401),
.B1(n_424),
.B2(n_419),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_408),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_502),
.B(n_517),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_451),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_503),
.B(n_513),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_402),
.Y(n_504)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_463),
.A2(n_417),
.B(n_414),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_506),
.A2(n_521),
.B(n_523),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_466),
.A2(n_467),
.B1(n_482),
.B2(n_464),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_507),
.Y(n_543)
);

XOR2x2_ASAP7_75t_L g509 ( 
.A(n_450),
.B(n_411),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_509),
.B(n_473),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_458),
.A2(n_465),
.B1(n_447),
.B2(n_459),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_476),
.A2(n_386),
.B1(n_341),
.B2(n_370),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_484),
.A2(n_386),
.B1(n_337),
.B2(n_341),
.Y(n_512)
);

OAI32xp33_ASAP7_75t_L g513 ( 
.A1(n_477),
.A2(n_355),
.A3(n_358),
.B1(n_377),
.B2(n_366),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_470),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_474),
.A2(n_481),
.B1(n_478),
.B2(n_449),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_516),
.A2(n_520),
.B1(n_526),
.B2(n_361),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_479),
.A2(n_360),
.B(n_370),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_460),
.B(n_366),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_474),
.A2(n_361),
.B1(n_365),
.B2(n_333),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_453),
.A2(n_375),
.B(n_345),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_485),
.B(n_333),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_522),
.B(n_528),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_443),
.A2(n_468),
.B(n_475),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_443),
.A2(n_376),
.B(n_373),
.C(n_358),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_524),
.B(n_5),
.Y(n_567)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_444),
.A2(n_461),
.B1(n_483),
.B2(n_475),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_468),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_532),
.A2(n_503),
.B1(n_495),
.B2(n_489),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_560),
.Y(n_569)
);

MAJx2_ASAP7_75t_L g571 ( 
.A(n_537),
.B(n_538),
.C(n_548),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_499),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_539),
.B(n_555),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_514),
.B(n_365),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_541),
.B(n_519),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_494),
.A2(n_472),
.B(n_486),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_542),
.A2(n_562),
.B(n_566),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_545),
.A2(n_547),
.B1(n_552),
.B2(n_556),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_349),
.C(n_276),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_559),
.C(n_518),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_498),
.A2(n_349),
.B1(n_372),
.B2(n_315),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_188),
.Y(n_553)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_553),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_17),
.Y(n_554)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_554),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_499),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_510),
.A2(n_507),
.B1(n_516),
.B2(n_500),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_497),
.B(n_17),
.Y(n_557)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_557),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_19),
.Y(n_558)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_490),
.B(n_345),
.C(n_372),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_508),
.B(n_19),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_506),
.A2(n_2),
.B(n_3),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_508),
.B(n_5),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_487),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_505),
.B(n_3),
.Y(n_564)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_564),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_523),
.Y(n_565)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_565),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_517),
.A2(n_494),
.B(n_488),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_564),
.B(n_565),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_568),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_573),
.B(n_578),
.Y(n_607)
);

CKINVDCx14_ASAP7_75t_R g624 ( 
.A(n_575),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_548),
.B(n_509),
.C(n_526),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_577),
.C(n_594),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_509),
.C(n_522),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_491),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_580),
.B(n_583),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_532),
.B(n_491),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_537),
.B(n_494),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_584),
.B(n_586),
.Y(n_625)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_535),
.Y(n_585)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_585),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_545),
.A2(n_489),
.B1(n_496),
.B2(n_494),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_587),
.A2(n_588),
.B1(n_590),
.B2(n_544),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_556),
.A2(n_493),
.B1(n_524),
.B2(n_501),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_547),
.A2(n_501),
.B1(n_527),
.B2(n_525),
.Y(n_590)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_593),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_549),
.B(n_501),
.C(n_528),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_539),
.A2(n_511),
.B1(n_520),
.B2(n_512),
.Y(n_595)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_595),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_538),
.B(n_513),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_SL g616 ( 
.A(n_596),
.B(n_551),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_521),
.C(n_4),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_597),
.B(n_560),
.C(n_564),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_555),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_598)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_598),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_561),
.B(n_3),
.Y(n_599)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_592),
.A2(n_566),
.B(n_561),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_622),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_533),
.Y(n_603)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_603),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_606),
.A2(n_621),
.B1(n_595),
.B2(n_531),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_616),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_573),
.B(n_540),
.C(n_543),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_617),
.C(n_623),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_591),
.A2(n_544),
.B(n_529),
.C(n_542),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_612),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_591),
.A2(n_530),
.B(n_529),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_615),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_589),
.A2(n_530),
.B(n_543),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_580),
.B(n_576),
.C(n_577),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_571),
.B(n_533),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_618),
.B(n_626),
.C(n_584),
.Y(n_638)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_598),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_570),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_571),
.B(n_551),
.C(n_546),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_588),
.A2(n_546),
.B(n_542),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_583),
.C(n_594),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_628),
.B(n_632),
.Y(n_656)
);

BUFx24_ASAP7_75t_SL g630 ( 
.A(n_624),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_630),
.B(n_646),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_604),
.B(n_596),
.C(n_586),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_617),
.B(n_569),
.C(n_578),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_633),
.B(n_637),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_623),
.B(n_581),
.Y(n_636)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_636),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_619),
.A2(n_581),
.B1(n_590),
.B2(n_587),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_638),
.B(n_639),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_569),
.C(n_542),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_642),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_607),
.B(n_531),
.C(n_552),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_644),
.C(n_645),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_607),
.B(n_568),
.C(n_534),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_534),
.C(n_550),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_609),
.A2(n_574),
.B1(n_572),
.B2(n_579),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_609),
.A2(n_579),
.B1(n_567),
.B2(n_582),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_614),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_620),
.B(n_550),
.C(n_597),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_648),
.B(n_625),
.C(n_615),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_651),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_640),
.A2(n_641),
.B1(n_635),
.B2(n_629),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_L g652 ( 
.A(n_634),
.B(n_618),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_652),
.A2(n_659),
.B(n_658),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_628),
.B(n_625),
.C(n_601),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_660),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_627),
.B(n_616),
.C(n_600),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_606),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_662),
.B(n_665),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_636),
.A2(n_603),
.B1(n_613),
.B2(n_611),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_663),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_602),
.Y(n_664)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_605),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_632),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_627),
.C(n_633),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_668),
.B(n_670),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_660),
.A2(n_642),
.B(n_631),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_669),
.A2(n_671),
.B(n_673),
.Y(n_683)
);

BUFx24_ASAP7_75t_SL g670 ( 
.A(n_653),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_657),
.A2(n_631),
.B(n_626),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_SL g672 ( 
.A(n_661),
.B(n_643),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_672),
.B(n_650),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_656),
.A2(n_612),
.B(n_645),
.Y(n_673)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_674),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_677),
.A2(n_654),
.B(n_663),
.Y(n_684)
);

XOR2xp5_ASAP7_75t_L g678 ( 
.A(n_675),
.B(n_649),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_678),
.B(n_685),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_666),
.B(n_649),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_679),
.B(n_681),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_667),
.B(n_662),
.C(n_661),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_666),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_688),
.B(n_681),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_680),
.A2(n_667),
.B(n_676),
.Y(n_689)
);

A2O1A1O1Ixp25_ASAP7_75t_L g691 ( 
.A1(n_689),
.A2(n_679),
.B(n_682),
.C(n_683),
.D(n_678),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_690),
.B(n_691),
.Y(n_692)
);

MAJx2_ASAP7_75t_L g693 ( 
.A(n_692),
.B(n_687),
.C(n_686),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_693),
.B(n_611),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_621),
.C(n_608),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_562),
.Y(n_696)
);


endmodule