module real_jpeg_3885_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_0),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_0),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_0),
.B(n_137),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_0),
.B(n_184),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_0),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_0),
.B(n_312),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_1),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_2),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_2),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_4),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_4),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_189),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_4),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_4),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_4),
.B(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_4),
.B(n_146),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_56),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_5),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_5),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_215),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_6),
.Y(n_148)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_8),
.Y(n_191)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_8),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_8),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_8),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_9),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_9),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_9),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_62),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_9),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_9),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_9),
.B(n_421),
.Y(n_420)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_11),
.B(n_48),
.Y(n_171)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_11),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_11),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_11),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_11),
.B(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_12),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_12),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_12),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_13),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_13),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_13),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_13),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_13),
.B(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_15),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_15),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_15),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_15),
.B(n_215),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_15),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_15),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_16),
.B(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_16),
.B(n_71),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_16),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_16),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_16),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_16),
.B(n_361),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_17),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_17),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_17),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_17),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_17),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_17),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_18),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_18),
.B(n_69),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_18),
.B(n_200),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_18),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_18),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_18),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_18),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_18),
.B(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_538),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_23),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_44),
.B(n_80),
.C(n_537),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_51),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_27),
.B(n_51),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.C(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_29),
.A2(n_33),
.B1(n_43),
.B2(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_33),
.B(n_55),
.C(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_36),
.Y(n_195)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_37),
.Y(n_202)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_37),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_50),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_76),
.C(n_78),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.C(n_66),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_60),
.B1(n_72),
.B2(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_56),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_57),
.Y(n_359)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_58),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_58),
.Y(n_394)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_58),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_67),
.C(n_72),
.Y(n_66)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_66),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_68),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_72),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_507)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_75),
.Y(n_339)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_75),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_122),
.B(n_536),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_119),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_82),
.B(n_119),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_116),
.C(n_117),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_83),
.A2(n_84),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_100),
.C(n_112),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_85),
.A2(n_86),
.B1(n_511),
.B2(n_513),
.Y(n_510)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_98),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_92),
.B(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_501)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_100),
.A2(n_112),
.B1(n_113),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_100),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_111),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_101),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_103),
.Y(n_265)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_106),
.A2(n_107),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_107),
.B(n_199),
.C(n_204),
.Y(n_508)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_110),
.Y(n_290)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_116),
.B(n_117),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_530),
.B(n_535),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_494),
.B(n_527),
.Y(n_123)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_295),
.B(n_493),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_244),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_126),
.B(n_244),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_196),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_127),
.B(n_197),
.C(n_226),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_169),
.C(n_178),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_128),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_143),
.C(n_158),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_129),
.B(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_136),
.C(n_140),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_134),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_143),
.A2(n_144),
.B1(n_158),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_154),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_145),
.B(n_154),
.Y(n_469)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_148),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_149),
.B(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_158),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_159),
.B(n_161),
.C(n_166),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_163),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_164),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_204),
.C(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_165),
.A2(n_166),
.B1(n_204),
.B2(n_207),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_178),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_175),
.C(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_172),
.A2(n_176),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_174),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_176),
.B(n_231),
.C(n_237),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_190),
.C(n_192),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_179),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_187),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_180),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_183),
.B(n_187),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_190),
.B(n_192),
.Y(n_273)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_195),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_226),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_198),
.B(n_209),
.C(n_225),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_217),
.B1(n_224),
.B2(n_225),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_214),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_218),
.B(n_220),
.C(n_223),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_228),
.B(n_230),
.C(n_238),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_246),
.B(n_249),
.Y(n_489)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_251),
.B(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_271),
.C(n_274),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_253),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_262),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_254),
.A2(n_255),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_257),
.A2(n_258),
.B(n_261),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_257),
.B(n_262),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_437)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_268),
.B(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_269),
.B(n_372),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_274),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_286),
.C(n_291),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_276),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.C(n_283),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_277),
.B(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_279),
.A2(n_283),
.B1(n_284),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_279),
.Y(n_450)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_286),
.B(n_291),
.Y(n_471)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_487),
.B(n_492),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_474),
.B(n_486),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_456),
.B(n_473),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_430),
.B(n_455),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_398),
.B(n_429),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_364),
.B(n_397),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_341),
.B(n_363),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_319),
.B(n_340),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_316),
.B(n_318),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_314),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_314),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_311),
.Y(n_320)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_321),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_329),
.B2(n_330),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_332),
.C(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_327),
.Y(n_352)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_336),
.B2(n_337),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_362),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_362),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_353),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_352),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_352),
.C(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_349),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_383),
.C(n_384),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_360),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_367),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_381),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_382),
.C(n_385),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_371),
.C(n_374),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_377),
.B1(n_378),
.B2(n_380),
.Y(n_374)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_375),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_392),
.C(n_395),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_392),
.B1(n_395),
.B2(n_396),
.Y(n_388)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_389),
.Y(n_395)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_392),
.Y(n_396)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_428),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_428),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_409),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_408),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_408),
.C(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_407),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_444),
.C(n_445),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_419),
.C(n_426),
.Y(n_433)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_410),
.Y(n_543)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.CI(n_414),
.CON(n_410),
.SN(n_410)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_413),
.C(n_414),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_426),
.B2(n_427),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_425),
.Y(n_440)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_453),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_453),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_442),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_434),
.C(n_442),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_465),
.C(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_440),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_447),
.C(n_452),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_452),
.Y(n_446)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_448),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_472),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_472),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_463),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_462),
.C(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_468),
.C(n_470),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_484),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_484),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_481),
.C(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_490),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_522),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_515),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_515),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_498),
.B1(n_504),
.B2(n_514),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_505),
.C(n_510),
.Y(n_534)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.C(n_502),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_499),
.B(n_518),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_500),
.A2(n_502),
.B1(n_503),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_504),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_510),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.C(n_509),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_506),
.B(n_508),
.CI(n_509),
.CON(n_520),
.SN(n_520)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_520),
.C(n_521),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_517),
.B1(n_520),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_520),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_520),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_524),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_526),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);


endmodule