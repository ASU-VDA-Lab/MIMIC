module fake_jpeg_2014_n_554 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_554);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_554;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_0),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_0),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_64),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_1),
.C(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_37),
.C(n_47),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_101),
.Y(n_112)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_30),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_89),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_5),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_95),
.Y(n_157)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_20),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_96),
.B(n_100),
.Y(n_163)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_5),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_37),
.B(n_17),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_52),
.B1(n_39),
.B2(n_51),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_20),
.B1(n_41),
.B2(n_43),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_147),
.B1(n_154),
.B2(n_158),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_24),
.B1(n_35),
.B2(n_23),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_118),
.B(n_79),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_55),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_78),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_63),
.A2(n_24),
.B1(n_35),
.B2(n_23),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_56),
.A2(n_46),
.B1(n_43),
.B2(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_165),
.B1(n_47),
.B2(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_52),
.B1(n_28),
.B2(n_51),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_63),
.A2(n_24),
.B1(n_35),
.B2(n_53),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_43),
.B1(n_46),
.B2(n_53),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_53),
.B1(n_44),
.B2(n_46),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_102),
.A2(n_69),
.B1(n_75),
.B2(n_73),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_57),
.C(n_71),
.Y(n_200)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_54),
.B1(n_21),
.B2(n_25),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_62),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_169),
.B(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_87),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_80),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_181),
.Y(n_243)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_173),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_112),
.A2(n_37),
.B(n_104),
.C(n_39),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_27),
.Y(n_241)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_177),
.A2(n_136),
.B1(n_111),
.B2(n_142),
.Y(n_249)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_21),
.B(n_25),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_180),
.B(n_210),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_81),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_182),
.B(n_184),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_81),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_77),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_192),
.B(n_133),
.Y(n_257)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_67),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_204),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_79),
.B(n_97),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_223),
.C(n_132),
.Y(n_236)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_84),
.B1(n_92),
.B2(n_68),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_202),
.A2(n_117),
.B1(n_144),
.B2(n_129),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_26),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

BUFx4f_ASAP7_75t_SL g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_120),
.B(n_165),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_222),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_272)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_137),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_218),
.A2(n_221),
.B1(n_146),
.B2(n_148),
.Y(n_265)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_115),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_115),
.B(n_111),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_159),
.B(n_31),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_151),
.B(n_113),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_226),
.A2(n_233),
.B1(n_235),
.B2(n_247),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_93),
.B1(n_26),
.B2(n_31),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_231),
.A2(n_249),
.B1(n_220),
.B2(n_209),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_160),
.B1(n_166),
.B2(n_137),
.Y(n_233)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_212),
.B1(n_202),
.B2(n_179),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_236),
.B(n_257),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_184),
.C(n_182),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_238),
.C(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_182),
.C(n_180),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g286 ( 
.A(n_241),
.B(n_223),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_167),
.B1(n_156),
.B2(n_136),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_132),
.C(n_142),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_179),
.A2(n_156),
.B1(n_133),
.B2(n_113),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_251),
.A2(n_224),
.B1(n_216),
.B2(n_213),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_175),
.B(n_153),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_266),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_197),
.A2(n_146),
.B1(n_91),
.B2(n_148),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_218),
.B1(n_199),
.B2(n_198),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_5),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_174),
.B(n_138),
.C(n_60),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_176),
.C(n_188),
.Y(n_295)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_273),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_192),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_284),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_278),
.A2(n_227),
.B1(n_266),
.B2(n_252),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_185),
.B1(n_211),
.B2(n_203),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_226),
.B1(n_247),
.B2(n_256),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_203),
.B1(n_211),
.B2(n_183),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_280),
.A2(n_291),
.B1(n_300),
.B2(n_260),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_281),
.B(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_177),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_286),
.A2(n_294),
.B(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_223),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_311),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_205),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_301),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_293),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_256),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_263),
.A2(n_173),
.B(n_193),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_241),
.A2(n_209),
.B(n_195),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_238),
.B(n_138),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_263),
.A2(n_201),
.B(n_191),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_260),
.B(n_253),
.Y(n_350)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_138),
.C(n_60),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_308),
.Y(n_351)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_168),
.C(n_186),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_208),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_225),
.B(n_189),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_313),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_225),
.B(n_178),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_228),
.B(n_6),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_301),
.C(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_354),
.C(n_327),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_332),
.B1(n_336),
.B2(n_346),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_282),
.A2(n_235),
.B1(n_249),
.B2(n_243),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_331),
.B1(n_341),
.B2(n_347),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_326),
.A2(n_330),
.B(n_353),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_276),
.A2(n_233),
.B1(n_251),
.B2(n_258),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_282),
.A2(n_242),
.B1(n_257),
.B2(n_265),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_242),
.B1(n_271),
.B2(n_248),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_274),
.A2(n_271),
.B1(n_245),
.B2(n_254),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_277),
.B(n_257),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_277),
.B(n_244),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_274),
.A2(n_244),
.B1(n_230),
.B2(n_245),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_254),
.B1(n_230),
.B2(n_239),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_310),
.A2(n_311),
.B1(n_276),
.B2(n_275),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_350),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_269),
.B(n_253),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_250),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_289),
.A2(n_239),
.B1(n_240),
.B2(n_270),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_292),
.B1(n_293),
.B2(n_288),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_261),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_310),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_355),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_322),
.A2(n_310),
.B1(n_291),
.B2(n_315),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_331),
.B1(n_332),
.B2(n_337),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_329),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_380),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_294),
.B(n_303),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_366),
.A2(n_374),
.B(n_334),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_308),
.B1(n_300),
.B2(n_287),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_367),
.A2(n_372),
.B1(n_346),
.B2(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_322),
.B1(n_335),
.B2(n_338),
.Y(n_369)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_373),
.C(n_382),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_352),
.B(n_296),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_371),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_283),
.B1(n_298),
.B2(n_306),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_295),
.C(n_307),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_302),
.B(n_299),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_381),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_297),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_273),
.C(n_270),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_351),
.C(n_353),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_316),
.B(n_240),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_391),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_6),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_386),
.Y(n_405)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_6),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_390),
.Y(n_415)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_336),
.B(n_6),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_406),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_394),
.A2(n_420),
.B1(n_367),
.B2(n_366),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_343),
.B(n_350),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_396),
.A2(n_404),
.B(n_419),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_361),
.B(n_351),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_398),
.B(n_409),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_7),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_333),
.B(n_342),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_339),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_339),
.C(n_333),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_408),
.C(n_418),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_342),
.C(n_344),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_365),
.B(n_344),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_378),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_376),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_417),
.B(n_387),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_372),
.C(n_365),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_358),
.A2(n_334),
.B1(n_345),
.B2(n_99),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_364),
.B(n_345),
.C(n_88),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_398),
.C(n_409),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_426),
.A2(n_427),
.B1(n_437),
.B2(n_395),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_399),
.A2(n_358),
.B1(n_363),
.B2(n_423),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_414),
.B(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_430),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_419),
.B(n_364),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_432),
.C(n_435),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_362),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_374),
.C(n_357),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_439),
.C(n_440),
.Y(n_465)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_436),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_399),
.A2(n_358),
.B1(n_389),
.B2(n_388),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_380),
.C(n_386),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_390),
.C(n_381),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_415),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_444),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_443),
.B(n_447),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_400),
.B(n_377),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_379),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_448),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_404),
.A2(n_359),
.B(n_27),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_446),
.A2(n_424),
.B(n_411),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_38),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_38),
.C(n_48),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_451),
.C(n_452),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_38),
.C(n_48),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_394),
.B(n_38),
.C(n_27),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_412),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_449),
.A2(n_422),
.B1(n_401),
.B2(n_402),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_458),
.Y(n_483)
);

BUFx12f_ASAP7_75t_SL g455 ( 
.A(n_441),
.Y(n_455)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_474),
.C(n_430),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_401),
.B1(n_396),
.B2(n_420),
.Y(n_456)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_429),
.A2(n_446),
.B1(n_445),
.B2(n_441),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_466),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_460),
.B(n_472),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_433),
.A2(n_412),
.B1(n_405),
.B2(n_410),
.Y(n_466)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_469),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_451),
.A2(n_413),
.B1(n_424),
.B2(n_411),
.Y(n_470)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_470),
.Y(n_482)
);

AO221x1_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_416),
.B1(n_405),
.B2(n_421),
.C(n_27),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_438),
.B(n_416),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_473),
.B(n_438),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_8),
.B(n_9),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_452),
.A2(n_38),
.B1(n_10),
.B2(n_12),
.Y(n_475)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_439),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_477),
.B(n_484),
.Y(n_506)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_465),
.B(n_425),
.Y(n_479)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_479),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_457),
.B(n_462),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_425),
.C(n_431),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_487),
.C(n_491),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_431),
.C(n_435),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_462),
.B(n_464),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_474),
.Y(n_508)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_450),
.C(n_447),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_492),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_38),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_480),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_499),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_454),
.B1(n_461),
.B2(n_463),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_495),
.A2(n_459),
.B(n_455),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_501),
.A2(n_491),
.B(n_478),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_466),
.C(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_502),
.B(n_511),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_495),
.A2(n_461),
.B1(n_481),
.B2(n_486),
.Y(n_505)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_505),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_483),
.A2(n_460),
.B1(n_471),
.B2(n_476),
.Y(n_507)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_493),
.C(n_494),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_510),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_481),
.A2(n_472),
.B1(n_468),
.B2(n_476),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_515),
.A2(n_512),
.B(n_504),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_487),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_516),
.B(n_520),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_519),
.A2(n_526),
.B(n_509),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_9),
.C(n_10),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_9),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_523),
.B(n_524),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_497),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_10),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_525),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_501),
.A2(n_10),
.B(n_12),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_12),
.C(n_13),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_504),
.B(n_503),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_530),
.Y(n_542)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_529),
.A2(n_535),
.B(n_536),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_513),
.B(n_502),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_514),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_531),
.B(n_533),
.Y(n_544)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_532),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_503),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_522),
.A2(n_511),
.B(n_500),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_525),
.C(n_527),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_541),
.A2(n_13),
.B(n_15),
.Y(n_548)
);

AOI211xp5_ASAP7_75t_L g543 ( 
.A1(n_537),
.A2(n_500),
.B(n_515),
.C(n_526),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_543),
.A2(n_545),
.B(n_537),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_535),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_546),
.A2(n_547),
.B(n_549),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_545),
.A2(n_520),
.B(n_538),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_548),
.A2(n_544),
.B(n_16),
.Y(n_551)
);

AOI321xp33_ASAP7_75t_L g549 ( 
.A1(n_540),
.A2(n_13),
.A3(n_16),
.B1(n_17),
.B2(n_539),
.C(n_542),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_550),
.C(n_13),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_17),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_17),
.Y(n_554)
);


endmodule