module real_jpeg_4099_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_2),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_159),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_2),
.A2(n_111),
.B1(n_112),
.B2(n_159),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_2),
.A2(n_159),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_3),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_4),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_4),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_5),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_203),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_5),
.A2(n_68),
.B1(n_203),
.B2(n_308),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_5),
.A2(n_155),
.B1(n_203),
.B2(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_80),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_80),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_36),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_10),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_11),
.A2(n_243),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_11),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_11),
.A2(n_37),
.B1(n_267),
.B2(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_11),
.A2(n_267),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_11),
.A2(n_93),
.B1(n_267),
.B2(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_13),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_13),
.A2(n_91),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_13),
.A2(n_91),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_13),
.A2(n_91),
.B1(n_188),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_14),
.A2(n_48),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_14),
.A2(n_48),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_15),
.A2(n_49),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_15),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_15),
.B(n_71),
.C(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_15),
.B(n_146),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_85),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_15),
.B(n_222),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_16),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_16),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_16),
.A2(n_69),
.B1(n_108),
.B2(n_243),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_16),
.A2(n_28),
.B1(n_108),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_16),
.A2(n_108),
.B1(n_318),
.B2(n_320),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_229),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_227),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_206),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_20),
.B(n_206),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_125),
.C(n_173),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_21),
.A2(n_22),
.B1(n_125),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_86),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_23),
.A2(n_24),
.B(n_88),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_24),
.A2(n_87),
.B1(n_88),
.B2(n_124),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_24),
.A2(n_46),
.B1(n_124),
.B2(n_428),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_25),
.A2(n_35),
.B1(n_176),
.B2(n_182),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_25),
.A2(n_252),
.B(n_257),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_25),
.A2(n_240),
.B(n_257),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_25),
.A2(n_392),
.B1(n_393),
.B2(n_396),
.Y(n_391)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_26),
.B(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_26),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_26),
.A2(n_326),
.B1(n_363),
.B2(n_368),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_26),
.A2(n_33),
.B1(n_397),
.B2(n_434),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_27),
.Y(n_296)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_39),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_46),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_79),
.B2(n_85),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_47),
.A2(n_56),
.B1(n_85),
.B2(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_51),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_52),
.Y(n_170)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_52),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_53),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_53),
.Y(n_339)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_56),
.A2(n_79),
.B1(n_85),
.B2(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_56),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_56),
.B(n_242),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_70),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_64),
.B2(n_68),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_70),
.A2(n_265),
.B(n_268),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_75),
.Y(n_400)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_76),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_76),
.Y(n_401)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_84),
.Y(n_309)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_85),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_85),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_92),
.Y(n_380)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_95),
.B(n_107),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_95),
.Y(n_212)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_96),
.B(n_240),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_96),
.A2(n_199),
.B1(n_200),
.B2(n_437),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_104),
.Y(n_96)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_97),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_99),
.Y(n_319)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_99),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_100),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_101),
.A2(n_378),
.A3(n_381),
.B1(n_383),
.B2(n_389),
.Y(n_377)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_102),
.Y(n_224)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_105),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_106),
.A2(n_212),
.B(n_437),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_SL g408 ( 
.A1(n_112),
.A2(n_240),
.B(n_389),
.Y(n_408)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_114),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_114),
.A2(n_408),
.B(n_409),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_125),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_165),
.B(n_172),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_146),
.B1(n_153),
.B2(n_160),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_128),
.A2(n_312),
.B(n_316),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_128),
.B(n_359),
.Y(n_358)
);

AOI22x1_ASAP7_75t_L g440 ( 
.A1(n_128),
.A2(n_146),
.B1(n_359),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_128),
.A2(n_316),
.B(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_129),
.A2(n_154),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_129),
.A2(n_197),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_129),
.A2(n_197),
.B1(n_353),
.B2(n_412),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_146),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_133),
.Y(n_336)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_135),
.Y(n_342)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_138),
.Y(n_416)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_145),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_145),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_145),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_146),
.Y(n_197)
);

AO22x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_157),
.Y(n_354)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_171),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_207),
.CI(n_208),
.CON(n_206),
.SN(n_206)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_173),
.B(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_192),
.C(n_198),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_174),
.B(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_186),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_175),
.B(n_186),
.Y(n_451)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_176),
.Y(n_434)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_179),
.Y(n_283)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_179),
.Y(n_365)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_185),
.Y(n_286)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_185),
.Y(n_395)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_187),
.Y(n_432)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_192),
.B(n_198),
.Y(n_426)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_193),
.Y(n_441)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_197),
.B(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_197),
.A2(n_353),
.B(n_358),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B(n_205),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_202),
.B(n_240),
.Y(n_389)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_205),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_206),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_226),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_225),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_238),
.B(n_241),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_216),
.A2(n_217),
.B1(n_265),
.B2(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_216),
.A2(n_241),
.B(n_307),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_216),
.A2(n_217),
.B1(n_418),
.B2(n_432),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_217),
.A2(n_268),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI311xp33_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_422),
.A3(n_459),
.B1(n_477),
.C1(n_478),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_371),
.B(n_421),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_344),
.B(n_370),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_301),
.B(n_343),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_271),
.B(n_300),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_250),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_236),
.B(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_245),
.B1(n_246),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_240),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g334 ( 
.A(n_243),
.Y(n_334)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_263),
.C(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_290),
.B(n_299),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B(n_289),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_288),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_284),
.B(n_287),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_325),
.B(n_331),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_303),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_323),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_310),
.B2(n_311),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_310),
.C(n_323),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_333),
.A3(n_334),
.B1(n_335),
.B2(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_332),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_332),
.Y(n_350)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_345),
.B(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_351),
.B2(n_369),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_350),
.C(n_369),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_360),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_361),
.C(n_362),
.Y(n_402)
);

INVx4_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_372),
.B(n_373),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_405),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_374)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_390),
.B2(n_391),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_402),
.B(n_403),
.C(n_405),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_410),
.B2(n_420),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_406),
.B(n_411),
.C(n_417),
.Y(n_468)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_412),
.Y(n_457)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_445),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_423),
.A2(n_445),
.B(n_479),
.C(n_482),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_442),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_442),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.C(n_429),
.Y(n_424)
);

FAx1_ASAP7_75t_SL g458 ( 
.A(n_425),
.B(n_427),
.CI(n_429),
.CON(n_458),
.SN(n_458)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_435),
.C(n_440),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_433),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_435),
.A2(n_436),
.B1(n_440),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_440),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_458),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_456),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_453),
.A2(n_454),
.B1(n_456),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_458),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.C(n_468),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_467),
.B1(n_468),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_474),
.Y(n_480)
);


endmodule