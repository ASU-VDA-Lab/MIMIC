module fake_jpeg_1086_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_48),
.Y(n_49)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_33),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_26),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_42),
.C(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_32),
.B(n_3),
.C(n_4),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_32),
.C(n_31),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_62),
.C(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_44),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_2),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_31),
.C(n_14),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_31),
.C(n_13),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_44),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_44),
.B(n_4),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_8),
.B(n_10),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_77),
.B(n_7),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_82),
.B1(n_72),
.B2(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_84),
.B1(n_81),
.B2(n_73),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_11),
.C(n_12),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_20),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_21),
.Y(n_91)
);


endmodule