module fake_aes_7574_n_1339 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1339);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1339;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_167), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_253), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_60), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_76), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_181), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_95), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_52), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_105), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_189), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_180), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_256), .Y(n_300) );
INVxp33_ASAP7_75t_SL g301 ( .A(n_96), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_80), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_91), .Y(n_303) );
BUFx2_ASAP7_75t_SL g304 ( .A(n_103), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_249), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_44), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_146), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_20), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_134), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_11), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_279), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_260), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_88), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_1), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_204), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_110), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_136), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_28), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_233), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_235), .Y(n_321) );
INVxp33_ASAP7_75t_L g322 ( .A(n_29), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_264), .Y(n_323) );
INVxp33_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_196), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_153), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_221), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_207), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_218), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_286), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_165), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_115), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_30), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_127), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_144), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_231), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_129), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_158), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_38), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_220), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_65), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_148), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_52), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_66), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_124), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_228), .B(n_267), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_150), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_15), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_1), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_89), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_117), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_282), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_47), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_174), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_35), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_226), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_99), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_141), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_168), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_285), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_169), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_208), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_61), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_247), .Y(n_365) );
INVxp33_ASAP7_75t_L g366 ( .A(n_92), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_45), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_212), .Y(n_368) );
INVxp33_ASAP7_75t_SL g369 ( .A(n_51), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_26), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_164), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_140), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_131), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_8), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_224), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_186), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_125), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_31), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_10), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_142), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_145), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_83), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_38), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_32), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_216), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_194), .Y(n_386) );
INVxp33_ASAP7_75t_SL g387 ( .A(n_161), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_163), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_2), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_100), .B(n_243), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_114), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_184), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_70), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_65), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_44), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_245), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_37), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_270), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_60), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_205), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_18), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_61), .Y(n_402) );
INVxp33_ASAP7_75t_L g403 ( .A(n_262), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_17), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_23), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_133), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_213), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_21), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_261), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_69), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_273), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_147), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_254), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_274), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_8), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_237), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_97), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_112), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_265), .Y(n_419) );
INVxp33_ASAP7_75t_L g420 ( .A(n_50), .Y(n_420) );
INVxp33_ASAP7_75t_L g421 ( .A(n_239), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_93), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_206), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_241), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_122), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_284), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_201), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_55), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_94), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_188), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_130), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_120), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_25), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_305), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_369), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_322), .B(n_0), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_305), .Y(n_437) );
BUFx8_ASAP7_75t_L g438 ( .A(n_380), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_325), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_355), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_305), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_314), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_294), .Y(n_443) );
NAND2xp33_ASAP7_75t_L g444 ( .A(n_321), .B(n_75), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_314), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_297), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_343), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_427), .B(n_3), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_343), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_350), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_350), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_297), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_291), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_338), .B(n_416), .Y(n_454) );
INVxp33_ASAP7_75t_L g455 ( .A(n_322), .Y(n_455) );
INVx6_ASAP7_75t_L g456 ( .A(n_297), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_4), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_293), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_297), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_315), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_321), .B(n_4), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_294), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_306), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_338), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_306), .B(n_5), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_295), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_292), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_452), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_436), .A2(n_420), .B1(n_333), .B2(n_341), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_437), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_438), .B(n_324), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_441), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_455), .B(n_324), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_454), .B(n_313), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_455), .A2(n_349), .B1(n_354), .B2(n_318), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_454), .B(n_366), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_467), .B(n_374), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_454), .B(n_385), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_436), .A2(n_339), .B1(n_370), .B2(n_356), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_441), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_434), .B(n_454), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_434), .B(n_416), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_436), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_454), .B(n_378), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_457), .B(n_308), .C(n_393), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_464), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
NOR3xp33_ASAP7_75t_SL g496 ( .A(n_439), .B(n_349), .C(n_318), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_464), .B(n_366), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_438), .B(n_403), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_467), .B(n_403), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_456), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_438), .B(n_421), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_443), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_457), .B(n_421), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_453), .B(n_365), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_453), .B(n_298), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_354), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_452), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_458), .B(n_373), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_504), .B(n_510), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_481), .B(n_440), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_510), .B(n_438), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_478), .B(n_448), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_492), .A2(n_461), .B1(n_448), .B2(n_369), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_478), .B(n_461), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_470), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_470), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_478), .B(n_458), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_504), .B(n_462), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_478), .B(n_466), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
NOR3xp33_ASAP7_75t_SL g529 ( .A(n_490), .B(n_401), .C(n_395), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_482), .B(n_466), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_487), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_481), .B(n_465), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_502), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_492), .A2(n_328), .B1(n_444), .B2(n_401), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_472), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_502), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_482), .B(n_289), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_482), .B(n_301), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_490), .A2(n_328), .B1(n_410), .B2(n_395), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_482), .A2(n_433), .B1(n_410), .B2(n_435), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_480), .B(n_289), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_487), .B(n_435), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_491), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_513), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_493), .B(n_299), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_508), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_513), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_472), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_491), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_494), .B(n_300), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_474), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_496), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_491), .B(n_442), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_501), .B(n_303), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_474), .Y(n_562) );
BUFx4f_ASAP7_75t_L g563 ( .A(n_494), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_476), .B(n_303), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_475), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_475), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_486), .Y(n_567) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_484), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_473), .B(n_301), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_484), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_503), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_511), .B(n_311), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_489), .Y(n_574) );
INVx5_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_515), .A2(n_387), .B1(n_433), .B2(n_312), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_495), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_507), .A2(n_296), .B1(n_364), .B2(n_387), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_512), .Y(n_581) );
INVxp67_ASAP7_75t_SL g582 ( .A(n_479), .Y(n_582) );
NOR2x2_ASAP7_75t_L g583 ( .A(n_496), .B(n_463), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_483), .B(n_302), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_469), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_497), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_471), .A2(n_445), .B1(n_447), .B2(n_442), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_497), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_505), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_498), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_505), .B(n_445), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_477), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_509), .B(n_311), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_509), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_509), .B(n_312), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_514), .B(n_447), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_514), .A2(n_404), .B1(n_383), .B2(n_384), .Y(n_600) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_514), .B(n_347), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_477), .B(n_307), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_477), .B(n_323), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_469), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_499), .B(n_465), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_499), .B(n_449), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_499), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_500), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_500), .B(n_345), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_521), .A2(n_368), .B(n_290), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
BUFx2_ASAP7_75t_SL g612 ( .A(n_532), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_532), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_578), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_519), .B(n_323), .Y(n_615) );
BUFx12f_ASAP7_75t_L g616 ( .A(n_553), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_542), .A2(n_348), .B(n_335), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_547), .B(n_304), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_581), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_519), .B(n_335), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_550), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_584), .A2(n_389), .B(n_394), .C(n_379), .Y(n_623) );
O2A1O1Ixp5_ASAP7_75t_SL g624 ( .A1(n_584), .A2(n_450), .B(n_451), .C(n_449), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_519), .B(n_348), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_547), .A2(n_516), .B1(n_582), .B2(n_549), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_554), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_567), .B(n_358), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_568), .A2(n_345), .B1(n_367), .B2(n_361), .Y(n_629) );
OAI21x1_ASAP7_75t_L g630 ( .A1(n_601), .A2(n_500), .B(n_309), .Y(n_630) );
INVx5_ASAP7_75t_L g631 ( .A(n_565), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_567), .B(n_358), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_565), .Y(n_633) );
OR2x6_ASAP7_75t_L g634 ( .A(n_547), .B(n_397), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_565), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_568), .A2(n_367), .B1(n_361), .B2(n_363), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_525), .A2(n_377), .B(n_317), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_565), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_536), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_572), .Y(n_640) );
CKINVDCx6p67_ASAP7_75t_R g641 ( .A(n_526), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_520), .A2(n_406), .B1(n_424), .B2(n_363), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_576), .B(n_406), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_560), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_542), .A2(n_424), .B1(n_402), .B2(n_405), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_530), .A2(n_320), .B(n_316), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_544), .A2(n_408), .B1(n_415), .B2(n_399), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_553), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_537), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_527), .B(n_428), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_450), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_518), .A2(n_451), .B(n_413), .C(n_327), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_609), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_537), .Y(n_655) );
AO22x1_ASAP7_75t_L g656 ( .A1(n_559), .A2(n_330), .B1(n_326), .B2(n_329), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_527), .A2(n_310), .B1(n_336), .B2(n_332), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_529), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_548), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_560), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_517), .B(n_337), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_549), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_556), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_556), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_531), .B(n_310), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_539), .B(n_310), .Y(n_666) );
INVx4_ASAP7_75t_L g667 ( .A(n_563), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_546), .A2(n_344), .B(n_346), .C(n_340), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_605), .B(n_351), .Y(n_669) );
OR2x6_ASAP7_75t_L g670 ( .A(n_533), .B(n_310), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_535), .B(n_352), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_557), .A2(n_357), .B(n_353), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_541), .B(n_359), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_538), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_577), .B(n_360), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_569), .B(n_362), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_538), .Y(n_677) );
O2A1O1Ixp5_ASAP7_75t_L g678 ( .A1(n_557), .A2(n_309), .B(n_331), .C(n_298), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_569), .A2(n_372), .B1(n_375), .B2(n_371), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_570), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_522), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_570), .A2(n_386), .B1(n_388), .B2(n_376), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_563), .B(n_392), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_564), .B(n_396), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_573), .B(n_5), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_574), .Y(n_687) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_534), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_588), .A2(n_414), .B1(n_432), .B2(n_425), .C1(n_423), .C2(n_422), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_529), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_580), .A2(n_411), .B1(n_412), .B2(n_398), .Y(n_691) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_534), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_555), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_561), .B(n_417), .Y(n_694) );
O2A1O1Ixp5_ASAP7_75t_SL g695 ( .A1(n_602), .A2(n_418), .B(n_426), .C(n_419), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_552), .A2(n_431), .B(n_429), .Y(n_696) );
BUFx3_ASAP7_75t_L g697 ( .A(n_593), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_522), .B(n_390), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_579), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_579), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g701 ( .A(n_559), .B(n_583), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_588), .B(n_6), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_600), .B(n_6), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_603), .A2(n_334), .B(n_331), .Y(n_704) );
INVx5_ASAP7_75t_L g705 ( .A(n_540), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_593), .Y(n_706) );
AND2x6_ASAP7_75t_L g707 ( .A(n_540), .B(n_334), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_558), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_562), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_L g710 ( .A1(n_566), .A2(n_342), .B(n_391), .C(n_400), .Y(n_710) );
AND2x6_ASAP7_75t_L g711 ( .A(n_545), .B(n_342), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_571), .A2(n_391), .B(n_400), .C(n_407), .Y(n_712) );
BUFx12f_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_523), .A2(n_409), .B(n_407), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_524), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_596), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_545), .Y(n_717) );
INVx4_ASAP7_75t_L g718 ( .A(n_575), .Y(n_718) );
INVx4_ASAP7_75t_L g719 ( .A(n_575), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_528), .A2(n_430), .B(n_409), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_590), .B(n_7), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_575), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_586), .A2(n_430), .B1(n_460), .B2(n_459), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_575), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_587), .B(n_7), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_606), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_606), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_589), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_599), .A2(n_459), .B(n_460), .C(n_315), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_551), .A2(n_460), .B(n_459), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_606), .Y(n_731) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_585), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_585), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_592), .B(n_9), .Y(n_734) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_598), .A2(n_9), .B(n_10), .C(n_11), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_599), .A2(n_382), .B(n_381), .C(n_319), .Y(n_736) );
INVx8_ASAP7_75t_L g737 ( .A(n_583), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g738 ( .A1(n_595), .A2(n_382), .B(n_381), .C(n_319), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_591), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_597), .B(n_12), .Y(n_740) );
OAI222xp33_ASAP7_75t_SL g741 ( .A1(n_608), .A2(n_12), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_608), .B(n_315), .Y(n_742) );
OR2x6_ASAP7_75t_SL g743 ( .A(n_594), .B(n_13), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_594), .B(n_14), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_607), .B(n_16), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_607), .A2(n_488), .B(n_469), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g747 ( .A1(n_626), .A2(n_315), .B1(n_319), .B2(n_381), .C1(n_382), .C2(n_456), .Y(n_747) );
OAI21x1_ASAP7_75t_SL g748 ( .A1(n_611), .A2(n_17), .B(n_18), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_704), .A2(n_604), .B(n_585), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_616), .Y(n_750) );
OAI21x1_ASAP7_75t_SL g751 ( .A1(n_611), .A2(n_19), .B(n_20), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_680), .B(n_585), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_621), .Y(n_753) );
OAI21x1_ASAP7_75t_SL g754 ( .A1(n_655), .A2(n_19), .B(n_21), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_614), .A2(n_382), .B1(n_381), .B2(n_319), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_619), .A2(n_456), .B1(n_604), .B2(n_24), .Y(n_756) );
OAI21x1_ASAP7_75t_L g757 ( .A1(n_624), .A2(n_604), .B(n_506), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_612), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_613), .B(n_22), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_655), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_627), .A2(n_629), .B1(n_634), .B2(n_636), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_680), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_634), .B(n_22), .Y(n_763) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_630), .A2(n_506), .B(n_488), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_746), .A2(n_506), .B(n_488), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_645), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_732), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_680), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_641), .B(n_23), .Y(n_769) );
BUFx2_ASAP7_75t_L g770 ( .A(n_713), .Y(n_770) );
OAI21x1_ASAP7_75t_L g771 ( .A1(n_695), .A2(n_506), .B(n_78), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_649), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_652), .B(n_618), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_622), .B(n_24), .Y(n_774) );
AND2x2_ASAP7_75t_SL g775 ( .A(n_721), .B(n_25), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_685), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_644), .B(n_26), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_685), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_725), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_678), .A2(n_79), .B(n_77), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_685), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_665), .A2(n_82), .B(n_81), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_618), .A2(n_456), .B1(n_28), .B2(n_29), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_670), .B(n_27), .Y(n_784) );
AO21x2_ASAP7_75t_L g785 ( .A1(n_736), .A2(n_85), .B(n_84), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_639), .A2(n_677), .B(n_650), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_702), .A2(n_27), .B1(n_30), .B2(n_31), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_693), .Y(n_788) );
OAI21xp5_ASAP7_75t_SL g789 ( .A1(n_642), .A2(n_32), .B(n_33), .Y(n_789) );
INVx3_ASAP7_75t_L g790 ( .A(n_645), .Y(n_790) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_732), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_735), .A2(n_33), .B(n_34), .C(n_35), .Y(n_792) );
INVx4_ASAP7_75t_L g793 ( .A(n_631), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_654), .A2(n_34), .B1(n_36), .B2(n_37), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_714), .A2(n_87), .B(n_86), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_L g796 ( .A1(n_668), .A2(n_36), .B(n_39), .C(n_40), .Y(n_796) );
BUFx4_ASAP7_75t_R g797 ( .A(n_697), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_666), .A2(n_98), .B(n_90), .Y(n_798) );
OAI21x1_ASAP7_75t_SL g799 ( .A1(n_709), .A2(n_39), .B(n_40), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_744), .A2(n_102), .B(n_101), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_670), .B(n_41), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g802 ( .A1(n_648), .A2(n_41), .B1(n_42), .B2(n_43), .C(n_45), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_671), .B(n_42), .Y(n_803) );
BUFx2_ASAP7_75t_L g804 ( .A(n_743), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_631), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_669), .B(n_43), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_728), .Y(n_807) );
AOI21x1_ASAP7_75t_L g808 ( .A1(n_720), .A2(n_175), .B(n_287), .Y(n_808) );
OR2x6_ASAP7_75t_L g809 ( .A(n_737), .B(n_46), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_737), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_707), .Y(n_811) );
OA21x2_ASAP7_75t_L g812 ( .A1(n_738), .A2(n_172), .B(n_283), .Y(n_812) );
OA21x2_ASAP7_75t_L g813 ( .A1(n_729), .A2(n_171), .B(n_281), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_721), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_674), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_633), .A2(n_176), .B(n_280), .Y(n_816) );
AO31x2_ASAP7_75t_L g817 ( .A1(n_709), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_699), .Y(n_818) );
OA21x2_ASAP7_75t_L g819 ( .A1(n_696), .A2(n_177), .B(n_278), .Y(n_819) );
A2O1A1Ixp33_ASAP7_75t_L g820 ( .A1(n_623), .A2(n_49), .B(n_51), .C(n_53), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_734), .A2(n_178), .B(n_277), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_700), .A2(n_170), .B(n_276), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_645), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_708), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_669), .B(n_53), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_617), .B(n_54), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_739), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_638), .A2(n_166), .B(n_275), .Y(n_828) );
OAI21x1_ASAP7_75t_L g829 ( .A1(n_742), .A2(n_162), .B(n_269), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_660), .B(n_54), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_687), .A2(n_179), .B(n_268), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_715), .A2(n_160), .B(n_266), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_646), .B(n_55), .Y(n_833) );
OAI21x1_ASAP7_75t_L g834 ( .A1(n_722), .A2(n_159), .B(n_263), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g835 ( .A1(n_610), .A2(n_157), .B(n_259), .Y(n_835) );
O2A1O1Ixp33_ASAP7_75t_L g836 ( .A1(n_676), .A2(n_56), .B(n_57), .C(n_58), .Y(n_836) );
OA21x2_ASAP7_75t_L g837 ( .A1(n_730), .A2(n_156), .B(n_258), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_631), .Y(n_838) );
OR2x2_ASAP7_75t_L g839 ( .A(n_703), .B(n_56), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_706), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_689), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_716), .B(n_59), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_710), .A2(n_183), .B(n_257), .Y(n_843) );
OA21x2_ASAP7_75t_L g844 ( .A1(n_694), .A2(n_182), .B(n_255), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_647), .A2(n_155), .B(n_252), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_667), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_727), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_686), .Y(n_848) );
INVx5_ASAP7_75t_L g849 ( .A(n_635), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_635), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_684), .A2(n_154), .B(n_251), .Y(n_851) );
AO31x2_ASAP7_75t_L g852 ( .A1(n_723), .A2(n_62), .A3(n_63), .B(n_64), .Y(n_852) );
OAI21x1_ASAP7_75t_L g853 ( .A1(n_722), .A2(n_187), .B(n_250), .Y(n_853) );
BUFx8_ASAP7_75t_L g854 ( .A(n_707), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_667), .B(n_66), .Y(n_855) );
INVx1_ASAP7_75t_SL g856 ( .A(n_707), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_707), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_635), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_726), .Y(n_859) );
NAND2x1_ASAP7_75t_L g860 ( .A(n_711), .B(n_104), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_726), .A2(n_731), .B1(n_651), .B2(n_673), .Y(n_861) );
INVx4_ASAP7_75t_L g862 ( .A(n_659), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_724), .A2(n_190), .B(n_248), .Y(n_863) );
OA21x2_ASAP7_75t_L g864 ( .A1(n_672), .A2(n_185), .B(n_246), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_745), .A2(n_152), .B(n_244), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_731), .Y(n_866) );
INVx1_ASAP7_75t_SL g867 ( .A(n_711), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_664), .Y(n_868) );
OAI21x1_ASAP7_75t_L g869 ( .A1(n_724), .A2(n_151), .B(n_242), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_659), .B(n_67), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_732), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_615), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_733), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_733), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_640), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_679), .B(n_68), .Y(n_876) );
OAI21x1_ASAP7_75t_SL g877 ( .A1(n_712), .A2(n_70), .B(n_71), .Y(n_877) );
INVx5_ASAP7_75t_L g878 ( .A(n_659), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_733), .Y(n_879) );
BUFx2_ASAP7_75t_L g880 ( .A(n_711), .Y(n_880) );
AO21x2_ASAP7_75t_L g881 ( .A1(n_675), .A2(n_192), .B(n_240), .Y(n_881) );
INVxp33_ASAP7_75t_L g882 ( .A(n_628), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_698), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_662), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_691), .A2(n_71), .B1(n_72), .B2(n_73), .C(n_74), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_637), .A2(n_620), .B(n_625), .Y(n_886) );
AOI21x1_ASAP7_75t_L g887 ( .A1(n_698), .A2(n_191), .B(n_238), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_653), .A2(n_149), .B(n_236), .Y(n_888) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_643), .A2(n_143), .B(n_234), .Y(n_889) );
OAI21x1_ASAP7_75t_L g890 ( .A1(n_682), .A2(n_139), .B(n_232), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_681), .B(n_72), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_632), .A2(n_195), .B(n_230), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_775), .A2(n_690), .B1(n_658), .B2(n_701), .Y(n_893) );
AO21x1_ASAP7_75t_L g894 ( .A1(n_870), .A2(n_661), .B(n_740), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_753), .Y(n_895) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_789), .A2(n_657), .B1(n_683), .B2(n_663), .C(n_688), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_807), .B(n_681), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_827), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_761), .A2(n_662), .B1(n_719), .B2(n_718), .C(n_741), .Y(n_899) );
INVx3_ASAP7_75t_L g900 ( .A(n_793), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_775), .A2(n_711), .B1(n_662), .B2(n_718), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_753), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_804), .A2(n_705), .B1(n_717), .B2(n_692), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_773), .B(n_719), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_752), .A2(n_705), .B(n_717), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_752), .A2(n_705), .B(n_717), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_861), .A2(n_692), .B1(n_656), .B2(n_73), .C(n_74), .Y(n_907) );
INVx3_ASAP7_75t_L g908 ( .A(n_793), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_833), .A2(n_692), .B1(n_107), .B2(n_108), .Y(n_909) );
AOI221x1_ASAP7_75t_SL g910 ( .A1(n_794), .A2(n_106), .B1(n_109), .B2(n_111), .C(n_113), .Y(n_910) );
NOR2x1_ASAP7_75t_SL g911 ( .A(n_809), .B(n_116), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_758), .A2(n_854), .B1(n_801), .B2(n_809), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_848), .A2(n_118), .B1(n_119), .B2(n_121), .C(n_123), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_758), .A2(n_854), .B1(n_809), .B2(n_855), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_760), .A2(n_126), .B1(n_128), .B2(n_132), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_886), .A2(n_135), .B(n_137), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_760), .A2(n_138), .B1(n_197), .B2(n_198), .Y(n_917) );
AOI21xp33_ASAP7_75t_SL g918 ( .A1(n_750), .A2(n_288), .B(n_200), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_861), .B(n_199), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_774), .A2(n_202), .B1(n_203), .B2(n_209), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_764), .A2(n_210), .B(n_211), .Y(n_921) );
BUFx3_ASAP7_75t_L g922 ( .A(n_772), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_788), .Y(n_923) );
OAI21xp5_ASAP7_75t_L g924 ( .A1(n_786), .A2(n_214), .B(n_215), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_833), .A2(n_217), .B1(n_219), .B2(n_222), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_779), .B(n_223), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_763), .A2(n_225), .B1(n_227), .B2(n_229), .Y(n_927) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_767), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_826), .A2(n_806), .B1(n_882), .B2(n_777), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_818), .Y(n_930) );
NAND2x1_ASAP7_75t_L g931 ( .A(n_818), .B(n_862), .Y(n_931) );
OAI21xp33_ASAP7_75t_L g932 ( .A1(n_792), .A2(n_826), .B(n_882), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_824), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_774), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_840), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_764), .A2(n_757), .B(n_765), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_868), .B(n_803), .Y(n_937) );
AND2x4_ASAP7_75t_L g938 ( .A(n_878), .B(n_811), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_870), .Y(n_939) );
INVxp67_ASAP7_75t_L g940 ( .A(n_842), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_774), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_878), .B(n_857), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_839), .A2(n_784), .B1(n_814), .B2(n_783), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_777), .A2(n_876), .B1(n_841), .B2(n_825), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_777), .A2(n_841), .B1(n_855), .B2(n_891), .Y(n_945) );
OA21x2_ASAP7_75t_L g946 ( .A1(n_757), .A2(n_771), .B(n_821), .Y(n_946) );
AND3x1_ASAP7_75t_L g947 ( .A(n_769), .B(n_885), .C(n_787), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_770), .B(n_759), .Y(n_948) );
OAI21xp33_ASAP7_75t_L g949 ( .A1(n_792), .A2(n_747), .B(n_820), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_859), .B(n_866), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_855), .A2(n_891), .B1(n_883), .B2(n_854), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_891), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_799), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_846), .B(n_805), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_888), .A2(n_768), .B(n_871), .Y(n_955) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_797), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_766), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_830), .B(n_762), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_820), .B(n_836), .C(n_796), .Y(n_959) );
AND2x4_ASAP7_75t_L g960 ( .A(n_878), .B(n_880), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_787), .A2(n_856), .B1(n_867), .B2(n_847), .Y(n_961) );
OAI21x1_ASAP7_75t_L g962 ( .A1(n_800), .A2(n_816), .B(n_828), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_802), .A2(n_872), .B1(n_877), .B2(n_875), .C(n_815), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_748), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_846), .B(n_805), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g966 ( .A1(n_772), .A2(n_751), .B1(n_754), .B2(n_797), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_838), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_847), .A2(n_756), .B1(n_810), .B2(n_750), .C(n_835), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_817), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_810), .A2(n_845), .B1(n_838), .B2(n_822), .C(n_755), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_878), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_852), .B(n_817), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_768), .A2(n_871), .B(n_879), .Y(n_973) );
AOI21xp5_ASAP7_75t_L g974 ( .A1(n_873), .A2(n_879), .B(n_874), .Y(n_974) );
AOI222xp33_ASAP7_75t_L g975 ( .A1(n_862), .A2(n_790), .B1(n_766), .B2(n_823), .C1(n_884), .C2(n_890), .Y(n_975) );
CKINVDCx6p67_ASAP7_75t_R g976 ( .A(n_849), .Y(n_976) );
OA21x2_ASAP7_75t_L g977 ( .A1(n_843), .A2(n_780), .B(n_795), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_817), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_852), .B(n_817), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_852), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_860), .A2(n_819), .B1(n_849), .B2(n_844), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_790), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_852), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_823), .A2(n_884), .B1(n_865), .B2(n_776), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_890), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_834), .Y(n_986) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_873), .A2(n_874), .B(n_767), .Y(n_987) );
OAI21x1_ASAP7_75t_L g988 ( .A1(n_782), .A2(n_798), .B(n_831), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_849), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_889), .A2(n_851), .B1(n_892), .B2(n_865), .C(n_778), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_853), .Y(n_991) );
OAI211xp5_ASAP7_75t_L g992 ( .A1(n_887), .A2(n_819), .B(n_844), .C(n_808), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_762), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_776), .A2(n_778), .B1(n_781), .B2(n_819), .Y(n_994) );
AND2x4_ASAP7_75t_L g995 ( .A(n_849), .B(n_781), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_844), .A2(n_767), .B1(n_791), .B2(n_850), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_863), .Y(n_997) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_881), .A2(n_785), .B1(n_850), .B2(n_858), .C(n_791), .Y(n_998) );
INVx2_ASAP7_75t_SL g999 ( .A(n_767), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_869), .Y(n_1000) );
AO21x2_ASAP7_75t_L g1001 ( .A1(n_843), .A2(n_881), .B(n_780), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_858), .A2(n_785), .B1(n_813), .B2(n_864), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_795), .B(n_813), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_791), .B(n_864), .Y(n_1004) );
INVx3_ASAP7_75t_L g1005 ( .A(n_791), .Y(n_1005) );
OA21x2_ASAP7_75t_L g1006 ( .A1(n_832), .A2(n_829), .B(n_837), .Y(n_1006) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_864), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_L g1008 ( .A1(n_813), .A2(n_886), .B(n_826), .C(n_796), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_812), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_812), .Y(n_1010) );
OAI21xp33_ASAP7_75t_L g1011 ( .A1(n_837), .A2(n_661), .B(n_526), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_837), .A2(n_775), .B1(n_760), .B2(n_774), .Y(n_1012) );
AND2x4_ASAP7_75t_SL g1013 ( .A(n_812), .B(n_772), .Y(n_1013) );
NOR2x1_ASAP7_75t_SL g1014 ( .A(n_809), .B(n_612), .Y(n_1014) );
OR2x6_ASAP7_75t_L g1015 ( .A(n_797), .B(n_612), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_848), .A2(n_492), .B1(n_516), .B2(n_669), .C(n_582), .Y(n_1016) );
OA21x2_ASAP7_75t_L g1017 ( .A1(n_757), .A2(n_749), .B(n_771), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_775), .A2(n_463), .B1(n_462), .B2(n_443), .Y(n_1018) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_761), .A2(n_443), .B1(n_462), .B2(n_634), .Y(n_1019) );
OAI221xp5_ASAP7_75t_L g1020 ( .A1(n_789), .A2(n_626), .B1(n_761), .B2(n_861), .C(n_544), .Y(n_1020) );
NAND2x1_ASAP7_75t_L g1021 ( .A(n_1012), .B(n_928), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_922), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1016), .B(n_1019), .Y(n_1023) );
AO21x2_ASAP7_75t_L g1024 ( .A1(n_936), .A2(n_992), .B(n_1009), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_929), .B(n_898), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_930), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_923), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_895), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_943), .B(n_937), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_933), .Y(n_1030) );
OAI21xp5_ASAP7_75t_L g1031 ( .A1(n_959), .A2(n_1008), .B(n_896), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_902), .B(n_980), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_945), .B(n_935), .Y(n_1033) );
INVx8_ASAP7_75t_L g1034 ( .A(n_1015), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_993), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_897), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_972), .B(n_979), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1004), .Y(n_1038) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_981), .A2(n_1011), .B(n_970), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_928), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_983), .B(n_967), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_897), .Y(n_1042) );
INVx3_ASAP7_75t_L g1043 ( .A(n_976), .Y(n_1043) );
OAI221xp5_ASAP7_75t_SL g1044 ( .A1(n_1020), .A2(n_1018), .B1(n_932), .B2(n_947), .C(n_914), .Y(n_1044) );
INVx4_ASAP7_75t_L g1045 ( .A(n_1015), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_952), .B(n_937), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_950), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_1015), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_940), .B(n_965), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_951), .B(n_934), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_912), .B(n_1020), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_941), .B(n_969), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_950), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_948), .B(n_904), .Y(n_1054) );
INVxp67_ASAP7_75t_L g1055 ( .A(n_954), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_928), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_978), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_985), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_926), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_926), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_1012), .Y(n_1061) );
NAND4xp25_ASAP7_75t_L g1062 ( .A(n_893), .B(n_910), .C(n_963), .D(n_968), .Y(n_1062) );
NAND2x1p5_ASAP7_75t_L g1063 ( .A(n_995), .B(n_931), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_971), .B(n_944), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_956), .B(n_900), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_900), .B(n_908), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1014), .B(n_901), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_986), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_903), .B(n_966), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_908), .B(n_953), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_989), .B(n_964), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_949), .B(n_896), .Y(n_1072) );
BUFx2_ASAP7_75t_L g1073 ( .A(n_939), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_938), .Y(n_1074) );
AND2x2_ASAP7_75t_SL g1075 ( .A(n_1013), .B(n_1010), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_958), .B(n_938), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_991), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_911), .B(n_995), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_957), .B(n_982), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_899), .Y(n_1080) );
INVxp67_ASAP7_75t_L g1081 ( .A(n_907), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_899), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_942), .B(n_960), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_942), .B(n_960), .Y(n_1084) );
INVx1_ASAP7_75t_SL g1085 ( .A(n_1005), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_907), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_920), .B(n_958), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_920), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_910), .B(n_961), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1005), .B(n_999), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_915), .B(n_917), .Y(n_1091) );
AOI21xp5_ASAP7_75t_L g1092 ( .A1(n_970), .A2(n_955), .B(n_996), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1000), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_915), .Y(n_1094) );
INVxp67_ASAP7_75t_L g1095 ( .A(n_919), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_917), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_961), .B(n_919), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_924), .B(n_984), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_894), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_975), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_909), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_997), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_924), .B(n_975), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1003), .B(n_925), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g1105 ( .A1(n_996), .A2(n_1007), .B1(n_977), .B2(n_916), .Y(n_1105) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_1017), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_905), .B(n_906), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_927), .B(n_974), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1017), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_918), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_973), .B(n_987), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_913), .B(n_990), .Y(n_1112) );
AO21x2_ASAP7_75t_L g1113 ( .A1(n_1001), .A2(n_962), .B(n_988), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1001), .B(n_946), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_946), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_994), .B(n_1002), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_977), .B(n_1006), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_998), .A2(n_1016), .B1(n_618), .B2(n_761), .C(n_804), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1006), .B(n_921), .Y(n_1119) );
OAI221xp5_ASAP7_75t_L g1120 ( .A1(n_1044), .A2(n_1118), .B1(n_1023), .B2(n_1051), .C(n_1029), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1121 ( .A(n_1028), .Y(n_1121) );
OAI31xp33_ASAP7_75t_L g1122 ( .A1(n_1062), .A2(n_1080), .A3(n_1082), .B(n_1072), .Y(n_1122) );
AO21x2_ASAP7_75t_L g1123 ( .A1(n_1092), .A2(n_1039), .B(n_1031), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1037), .B(n_1032), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1037), .B(n_1052), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1047), .B(n_1053), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1052), .B(n_1033), .Y(n_1127) );
OAI321xp33_ASAP7_75t_L g1128 ( .A1(n_1089), .A2(n_1091), .A3(n_1081), .B1(n_1069), .B2(n_1099), .C(n_1100), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1076), .Y(n_1129) );
A2O1A1Ixp33_ASAP7_75t_L g1130 ( .A1(n_1091), .A2(n_1034), .B(n_1088), .C(n_1094), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_1025), .A2(n_1086), .B1(n_1055), .B2(n_1054), .C(n_1033), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1038), .B(n_1057), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1038), .B(n_1087), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1058), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1135 ( .A1(n_1027), .A2(n_1030), .B1(n_1042), .B2(n_1036), .C(n_1050), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_1034), .A2(n_1050), .B1(n_1045), .B2(n_1096), .Y(n_1136) );
BUFx2_ASAP7_75t_L g1137 ( .A(n_1075), .Y(n_1137) );
NOR2x1_ASAP7_75t_L g1138 ( .A(n_1045), .B(n_1070), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1032), .B(n_1041), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1068), .Y(n_1140) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_1111), .B(n_1107), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1041), .B(n_1076), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1087), .B(n_1046), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1068), .Y(n_1144) );
BUFx6f_ASAP7_75t_L g1145 ( .A(n_1107), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1026), .B(n_1035), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1077), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1071), .B(n_1097), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1077), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1026), .B(n_1035), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1151 ( .A1(n_1064), .A2(n_1034), .B1(n_1059), .B2(n_1060), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1093), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1061), .B(n_1064), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1093), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1103), .B(n_1098), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1115), .Y(n_1156) );
BUFx6f_ASAP7_75t_L g1157 ( .A(n_1107), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1103), .B(n_1098), .Y(n_1158) );
AO22x1_ASAP7_75t_L g1159 ( .A1(n_1045), .A2(n_1048), .B1(n_1078), .B2(n_1043), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1097), .B(n_1073), .Y(n_1160) );
OR2x6_ASAP7_75t_L g1161 ( .A(n_1034), .B(n_1021), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1073), .B(n_1079), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1102), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1164 ( .A1(n_1049), .A2(n_1071), .A3(n_1070), .B1(n_1110), .B2(n_1067), .B3(n_1065), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1083), .B(n_1084), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1102), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1117), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1116), .B(n_1065), .Y(n_1168) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1109), .Y(n_1169) );
NAND4xp25_ASAP7_75t_SL g1170 ( .A(n_1022), .B(n_1083), .C(n_1084), .D(n_1078), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1117), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1106), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1079), .B(n_1116), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1111), .B(n_1104), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1106), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1104), .B(n_1095), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1114), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1178 ( .A(n_1066), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1066), .B(n_1090), .Y(n_1179) );
INVx4_ASAP7_75t_L g1180 ( .A(n_1043), .Y(n_1180) );
AND2x4_ASAP7_75t_SL g1181 ( .A(n_1043), .B(n_1022), .Y(n_1181) );
INVx1_ASAP7_75t_SL g1182 ( .A(n_1074), .Y(n_1182) );
AND2x4_ASAP7_75t_L g1183 ( .A(n_1040), .B(n_1056), .Y(n_1183) );
BUFx6f_ASAP7_75t_L g1184 ( .A(n_1113), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1185 ( .A1(n_1112), .A2(n_1101), .B(n_1108), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1063), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1114), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1021), .B(n_1085), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1090), .B(n_1119), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1101), .B(n_1063), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1063), .B(n_1024), .Y(n_1191) );
INVx3_ASAP7_75t_SL g1192 ( .A(n_1181), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1125), .B(n_1127), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1125), .B(n_1119), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1169), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1169), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1140), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1124), .B(n_1155), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_1120), .A2(n_1024), .B1(n_1105), .B2(n_1155), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1124), .B(n_1139), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1127), .B(n_1189), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1144), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1144), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1204 ( .A(n_1138), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1205 ( .A(n_1181), .B(n_1165), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1147), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1189), .B(n_1174), .Y(n_1207) );
OAI31xp33_ASAP7_75t_L g1208 ( .A1(n_1137), .A2(n_1170), .A3(n_1122), .B(n_1130), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1147), .Y(n_1209) );
NAND2xp5_ASAP7_75t_SL g1210 ( .A(n_1180), .B(n_1128), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1174), .B(n_1143), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1143), .B(n_1133), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1133), .B(n_1158), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1149), .Y(n_1214) );
CKINVDCx16_ASAP7_75t_R g1215 ( .A(n_1180), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1173), .B(n_1153), .Y(n_1216) );
INVxp67_ASAP7_75t_L g1217 ( .A(n_1121), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1149), .Y(n_1218) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1180), .B(n_1126), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1173), .B(n_1153), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1139), .B(n_1148), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1152), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1167), .B(n_1160), .Y(n_1223) );
NAND5xp2_ASAP7_75t_L g1224 ( .A(n_1131), .B(n_1136), .C(n_1151), .D(n_1185), .E(n_1135), .Y(n_1224) );
AND2x4_ASAP7_75t_L g1225 ( .A(n_1141), .B(n_1157), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1167), .B(n_1160), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1177), .B(n_1187), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1154), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1129), .B(n_1142), .Y(n_1229) );
NOR3xp33_ASAP7_75t_SL g1230 ( .A(n_1164), .B(n_1190), .C(n_1163), .Y(n_1230) );
AND2x2_ASAP7_75t_SL g1231 ( .A(n_1148), .B(n_1191), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1132), .B(n_1176), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1134), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1168), .B(n_1171), .Y(n_1234) );
AND2x4_ASAP7_75t_SL g1235 ( .A(n_1161), .B(n_1186), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1141), .B(n_1171), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1141), .B(n_1179), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1193), .B(n_1162), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1221), .Y(n_1239) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1195), .Y(n_1240) );
INVxp67_ASAP7_75t_L g1241 ( .A(n_1219), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1195), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1213), .B(n_1168), .Y(n_1243) );
AOI211x1_ASAP7_75t_L g1244 ( .A1(n_1210), .A2(n_1159), .B(n_1179), .C(n_1166), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1200), .B(n_1178), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1212), .B(n_1163), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1229), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1212), .B(n_1166), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1213), .B(n_1150), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1223), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1211), .B(n_1175), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1196), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1211), .B(n_1175), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1224), .B(n_1182), .Y(n_1254) );
AOI211xp5_ASAP7_75t_L g1255 ( .A1(n_1208), .A2(n_1159), .B(n_1157), .C(n_1145), .Y(n_1255) );
NAND4xp25_ASAP7_75t_L g1256 ( .A(n_1208), .B(n_1191), .C(n_1188), .D(n_1172), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1207), .B(n_1172), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1207), .B(n_1123), .Y(n_1258) );
AND2x4_ASAP7_75t_L g1259 ( .A(n_1225), .B(n_1157), .Y(n_1259) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1217), .B(n_1123), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1226), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1201), .B(n_1157), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1236), .B(n_1145), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1198), .B(n_1145), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1216), .B(n_1146), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1216), .B(n_1183), .Y(n_1266) );
INVx3_ASAP7_75t_L g1267 ( .A(n_1215), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1226), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1232), .B(n_1156), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1246), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1248), .Y(n_1271) );
AOI222xp33_ASAP7_75t_L g1272 ( .A1(n_1254), .A2(n_1231), .B1(n_1220), .B2(n_1199), .C1(n_1192), .C2(n_1194), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_1255), .A2(n_1192), .B1(n_1231), .B2(n_1205), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1269), .Y(n_1274) );
AOI22xp5_ASAP7_75t_L g1275 ( .A1(n_1254), .A2(n_1231), .B1(n_1192), .B2(n_1230), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1241), .B(n_1232), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1258), .B(n_1220), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1247), .B(n_1237), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1245), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1240), .Y(n_1280) );
HB1xp67_ASAP7_75t_L g1281 ( .A(n_1251), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1258), .Y(n_1282) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1240), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1239), .Y(n_1284) );
O2A1O1Ixp33_ASAP7_75t_L g1285 ( .A1(n_1256), .A2(n_1204), .B(n_1222), .C(n_1197), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1250), .Y(n_1286) );
OAI21xp33_ASAP7_75t_L g1287 ( .A1(n_1260), .A2(n_1227), .B(n_1234), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1262), .B(n_1225), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1261), .B(n_1234), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1242), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1268), .B(n_1218), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1290), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1290), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1282), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1282), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1281), .B(n_1262), .Y(n_1296) );
NAND2xp5_ASAP7_75t_SL g1297 ( .A(n_1273), .B(n_1244), .Y(n_1297) );
AOI21xp5_ASAP7_75t_L g1298 ( .A1(n_1285), .A2(n_1267), .B(n_1235), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1274), .Y(n_1299) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1280), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1291), .Y(n_1301) );
NAND2xp5_ASAP7_75t_SL g1302 ( .A(n_1272), .B(n_1253), .Y(n_1302) );
NAND2xp5_ASAP7_75t_SL g1303 ( .A(n_1275), .B(n_1253), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1288), .B(n_1257), .Y(n_1304) );
OAI221xp5_ASAP7_75t_SL g1305 ( .A1(n_1287), .A2(n_1243), .B1(n_1238), .B2(n_1266), .C(n_1264), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1299), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_1297), .A2(n_1276), .B1(n_1278), .B2(n_1279), .C(n_1284), .Y(n_1307) );
INVxp67_ASAP7_75t_L g1308 ( .A(n_1303), .Y(n_1308) );
INVx3_ASAP7_75t_L g1309 ( .A(n_1300), .Y(n_1309) );
AOI222xp33_ASAP7_75t_L g1310 ( .A1(n_1302), .A2(n_1278), .B1(n_1286), .B2(n_1270), .C1(n_1271), .C2(n_1277), .Y(n_1310) );
AOI21xp33_ASAP7_75t_L g1311 ( .A1(n_1301), .A2(n_1264), .B(n_1145), .Y(n_1311) );
AOI221x1_ASAP7_75t_L g1312 ( .A1(n_1298), .A2(n_1289), .B1(n_1288), .B2(n_1283), .C(n_1280), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1296), .B(n_1263), .Y(n_1313) );
O2A1O1Ixp33_ASAP7_75t_L g1314 ( .A1(n_1305), .A2(n_1283), .B(n_1249), .C(n_1265), .Y(n_1314) );
NOR2x1_ASAP7_75t_L g1315 ( .A(n_1296), .B(n_1209), .Y(n_1315) );
AOI222xp33_ASAP7_75t_L g1316 ( .A1(n_1307), .A2(n_1295), .B1(n_1294), .B2(n_1293), .C1(n_1292), .C2(n_1304), .Y(n_1316) );
OAI21xp5_ASAP7_75t_L g1317 ( .A1(n_1308), .A2(n_1295), .B(n_1294), .Y(n_1317) );
O2A1O1Ixp33_ASAP7_75t_L g1318 ( .A1(n_1310), .A2(n_1293), .B(n_1292), .C(n_1300), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g1319 ( .A(n_1315), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1314), .B(n_1214), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1321 ( .A(n_1306), .Y(n_1321) );
AOI221x1_ASAP7_75t_L g1322 ( .A1(n_1311), .A2(n_1214), .B1(n_1209), .B2(n_1206), .C(n_1233), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1321), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1320), .B(n_1309), .Y(n_1324) );
OAI22x1_ASAP7_75t_L g1325 ( .A1(n_1319), .A2(n_1312), .B1(n_1313), .B2(n_1259), .Y(n_1325) );
OAI211xp5_ASAP7_75t_SL g1326 ( .A1(n_1318), .A2(n_1228), .B(n_1203), .C(n_1202), .Y(n_1326) );
HB1xp67_ASAP7_75t_L g1327 ( .A(n_1323), .Y(n_1327) );
NOR3xp33_ASAP7_75t_L g1328 ( .A(n_1326), .B(n_1317), .C(n_1316), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1324), .B(n_1322), .Y(n_1329) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1327), .Y(n_1330) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_1329), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1328), .B(n_1325), .Y(n_1332) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_1330), .Y(n_1333) );
INVx3_ASAP7_75t_L g1334 ( .A(n_1332), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1331), .Y(n_1335) );
INVxp67_ASAP7_75t_SL g1336 ( .A(n_1335), .Y(n_1336) );
OAI21xp5_ASAP7_75t_L g1337 ( .A1(n_1336), .A2(n_1334), .B(n_1333), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1337), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_1338), .A2(n_1184), .B1(n_1252), .B2(n_1242), .Y(n_1339) );
endmodule