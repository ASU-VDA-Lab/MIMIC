module fake_jpeg_31038_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_15),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_0),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_66),
.B1(n_68),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_87),
.B1(n_90),
.B2(n_96),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_66),
.B1(n_63),
.B2(n_61),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_92),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_67),
.B1(n_72),
.B2(n_63),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_61),
.B1(n_71),
.B2(n_60),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_72),
.B(n_67),
.C(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_2),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_60),
.B1(n_73),
.B2(n_52),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_107),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_54),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_62),
.B1(n_59),
.B2(n_51),
.Y(n_106)
);

XNOR2x2_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_56),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_73),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_11),
.C(n_12),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_65),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_84),
.Y(n_122)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_20),
.B1(n_45),
.B2(n_43),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_117),
.B1(n_22),
.B2(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_12),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_19),
.B1(n_41),
.B2(n_39),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_84),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AO221x1_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_126),
.B1(n_135),
.B2(n_16),
.C(n_17),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_24),
.C(n_37),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_115),
.C(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_27),
.A3(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_11),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_38),
.B1(n_32),
.B2(n_31),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_134),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_105),
.B(n_98),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_149),
.B(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_109),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_148),
.C(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_117),
.C(n_30),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_13),
.B(n_15),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_149),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_121),
.B1(n_131),
.B2(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_152),
.B(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_144),
.C(n_143),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_154),
.B(n_157),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_164),
.A3(n_163),
.B1(n_140),
.B2(n_142),
.C1(n_150),
.C2(n_156),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_142),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_165),
.A3(n_148),
.B1(n_120),
.B2(n_128),
.C1(n_29),
.C2(n_18),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_17),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_18),
.Y(n_171)
);


endmodule