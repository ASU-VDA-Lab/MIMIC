module real_jpeg_8323_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_45),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_45),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_1),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_1),
.B(n_90),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_26),
.B(n_30),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_1),
.A2(n_24),
.B1(n_32),
.B2(n_129),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_8),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_8),
.A2(n_43),
.B1(n_45),
.B2(n_113),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_113),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_8),
.A2(n_24),
.B1(n_32),
.B2(n_113),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_9),
.A2(n_43),
.B1(n_45),
.B2(n_108),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_108),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_24),
.B1(n_32),
.B2(n_108),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_10),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_10),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_43),
.B1(n_45),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_11),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_120),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_11),
.A2(n_24),
.B1(n_32),
.B2(n_120),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_12),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_12),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_12),
.A2(n_33),
.B1(n_43),
.B2(n_45),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_14),
.A2(n_24),
.B1(n_32),
.B2(n_47),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_24),
.B1(n_32),
.B2(n_53),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_15),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_15),
.A2(n_43),
.B1(n_45),
.B2(n_53),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_72),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_20),
.A2(n_21),
.B1(n_68),
.B2(n_317),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_36),
.B1(n_37),
.B2(n_67),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_23),
.A2(n_28),
.B1(n_224),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_23),
.A2(n_28),
.B1(n_233),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_23),
.A2(n_252),
.B(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_23),
.A2(n_89),
.B(n_298),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_24),
.A2(n_25),
.B(n_129),
.C(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_31),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_40),
.B(n_41),
.C(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_41),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_30),
.B(n_129),
.CON(n_158),
.SN(n_158)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_39),
.A2(n_75),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_40),
.A2(n_49),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_40),
.A2(n_49),
.B1(n_77),
.B2(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_41),
.B(n_45),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_43),
.A2(n_50),
.B1(n_158),
.B2(n_164),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_56),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_46),
.A2(n_49),
.B(n_79),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_48),
.A2(n_80),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_65),
.C(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_54),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_58),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_58),
.B1(n_119),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_55),
.A2(n_58),
.B1(n_146),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_55),
.A2(n_156),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_55),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_55),
.A2(n_58),
.B1(n_239),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_55),
.A2(n_258),
.B(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_58),
.B(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_58),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_58),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_59),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_59),
.B(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_59),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_60),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_64),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_64),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_68),
.C(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_68),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_68),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_71),
.A2(n_90),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_72),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_78),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_75),
.A2(n_80),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_75),
.A2(n_80),
.B1(n_178),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_90),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_314),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_332),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_266),
.A3(n_290),
.B1(n_307),
.B2(n_313),
.C(n_333),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_226),
.C(n_262),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_197),
.B(n_225),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_171),
.B(n_196),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_151),
.B(n_170),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_140),
.B(n_150),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_126),
.B(n_139),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_109),
.B(n_168),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_132),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_125),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_134),
.B(n_138),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_133),
.B1(n_182),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_132),
.A2(n_167),
.B(n_207),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_132),
.A2(n_133),
.B(n_166),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_142),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_152),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.CI(n_147),
.CON(n_143),
.SN(n_143)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_148),
.B(n_183),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_162),
.B2(n_169),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_161),
.C(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_173),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_188),
.B2(n_189),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_191),
.C(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B1(n_180),
.B2(n_187),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_192),
.B(n_240),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_199),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_210),
.C(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_218),
.C(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_216),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_227),
.B(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.C(n_243),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_231),
.C(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_237),
.B1(n_243),
.B2(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_255),
.C(n_259),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_267),
.A2(n_308),
.B(n_312),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_268),
.B(n_269),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_289),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_282),
.B2(n_283),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_283),
.C(n_289),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_275),
.C(n_281),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_281),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_280),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_285),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_297),
.B(n_300),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_286),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_291),
.B(n_292),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_292),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_301),
.CI(n_306),
.CON(n_292),
.SN(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_299),
.B2(n_300),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_304),
.B(n_305),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_304),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_305),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_305),
.A2(n_316),
.B1(n_320),
.B2(n_328),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B(n_311),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_322),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.C(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);


endmodule