module fake_jpeg_3613_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_12),
.B(n_7),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_43),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_71),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_66),
.B1(n_64),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_88),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_64),
.B1(n_59),
.B2(n_51),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_56),
.B1(n_55),
.B2(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_66),
.B1(n_61),
.B2(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_74),
.B1(n_65),
.B2(n_57),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_76),
.B1(n_4),
.B2(n_5),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_49),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_50),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_52),
.B(n_70),
.C(n_2),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_1),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_105),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_76),
.B1(n_80),
.B2(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_121),
.B1(n_110),
.B2(n_123),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_16),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_42),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_40),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_99),
.B(n_94),
.C(n_105),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_143),
.B(n_145),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_19),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.C(n_21),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_135),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_5),
.B(n_6),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_145),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_6),
.B(n_7),
.Y(n_139)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_10),
.C(n_11),
.D(n_13),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_8),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_9),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_9),
.B(n_10),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_153),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_129),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_107),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_129),
.B1(n_125),
.B2(n_143),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_154)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_15),
.B1(n_29),
.B2(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_161),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_149),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_141),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_155),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_156),
.B(n_161),
.Y(n_177)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_148),
.A3(n_163),
.B1(n_159),
.B2(n_164),
.C(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.C(n_158),
.Y(n_178)
);

CKINVDCx11_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_130),
.C(n_171),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_172),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_151),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_R g185 ( 
.A(n_184),
.B(n_160),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_158),
.Y(n_186)
);


endmodule