module fake_netlist_5_517_n_4802 (n_137, n_924, n_676, n_294, n_431, n_318, n_380, n_419, n_977, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_1060, n_82, n_194, n_316, n_785, n_389, n_843, n_855, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_865, n_61, n_913, n_678, n_664, n_376, n_697, n_503, n_967, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_928, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_1055, n_916, n_452, n_885, n_397, n_493, n_111, n_525, n_880, n_703, n_698, n_980, n_483, n_544, n_683, n_1007, n_155, n_780, n_649, n_552, n_1057, n_1051, n_547, n_43, n_721, n_998, n_116, n_841, n_1050, n_956, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_983, n_139, n_38, n_105, n_280, n_744, n_1021, n_590, n_629, n_672, n_4, n_873, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_898, n_254, n_690, n_33, n_1013, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_1022, n_526, n_915, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_859, n_864, n_951, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_909, n_625, n_854, n_949, n_621, n_753, n_997, n_100, n_455, n_674, n_1008, n_932, n_417, n_946, n_1048, n_612, n_1001, n_212, n_385, n_498, n_516, n_933, n_788, n_507, n_119, n_497, n_689, n_738, n_912, n_606, n_559, n_275, n_640, n_968, n_252, n_624, n_825, n_26, n_295, n_133, n_1010, n_330, n_877, n_508, n_739, n_506, n_2, n_737, n_610, n_972, n_692, n_986, n_755, n_6, n_509, n_568, n_936, n_39, n_147, n_373, n_820, n_757, n_947, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_1024, n_556, n_106, n_209, n_259, n_448, n_758, n_999, n_668, n_733, n_991, n_375, n_301, n_828, n_779, n_576, n_941, n_929, n_981, n_1032, n_68, n_804, n_93, n_867, n_186, n_537, n_134, n_902, n_191, n_587, n_945, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_878, n_524, n_943, n_399, n_341, n_204, n_394, n_250, n_579, n_992, n_1049, n_938, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_984, n_320, n_694, n_518, n_505, n_286, n_883, n_122, n_282, n_752, n_331, n_10, n_905, n_906, n_24, n_406, n_519, n_470, n_908, n_782, n_919, n_325, n_449, n_132, n_862, n_90, n_900, n_724, n_856, n_546, n_1016, n_101, n_760, n_658, n_281, n_918, n_240, n_942, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_959, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_940, n_896, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_920, n_894, n_1046, n_271, n_934, n_1017, n_94, n_831, n_826, n_335, n_123, n_886, n_978, n_964, n_1054, n_654, n_370, n_167, n_976, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_1045, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_1033, n_988, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_1009, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_961, n_995, n_955, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_882, n_183, n_185, n_243, n_398, n_396, n_1036, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_897, n_215, n_350, n_196, n_798, n_662, n_459, n_1020, n_646, n_1062, n_211, n_218, n_400, n_930, n_181, n_436, n_962, n_3, n_290, n_580, n_221, n_178, n_622, n_1040, n_723, n_1035, n_386, n_578, n_994, n_926, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_1030, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_1043, n_496, n_355, n_958, n_849, n_1034, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_922, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_974, n_395, n_164, n_432, n_553, n_727, n_839, n_901, n_311, n_813, n_957, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_888, n_296, n_613, n_871, n_241, n_637, n_357, n_875, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_858, n_114, n_96, n_923, n_772, n_691, n_881, n_717, n_165, n_468, n_499, n_939, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_866, n_969, n_236, n_388, n_761, n_1012, n_1, n_1019, n_249, n_903, n_1006, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_889, n_80, n_973, n_35, n_73, n_277, n_1061, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_990, n_84, n_462, n_975, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_907, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_1031, n_263, n_471, n_609, n_852, n_989, n_1041, n_1039, n_44, n_224, n_40, n_34, n_228, n_283, n_1028, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_892, n_893, n_1015, n_1000, n_891, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_979, n_1002, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_874, n_465, n_838, n_76, n_358, n_1058, n_362, n_876, n_170, n_332, n_27, n_1053, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_953, n_601, n_279, n_917, n_1014, n_966, n_70, n_987, n_253, n_261, n_174, n_289, n_745, n_963, n_1052, n_954, n_627, n_767, n_172, n_206, n_217, n_993, n_440, n_726, n_478, n_793, n_545, n_982, n_441, n_860, n_450, n_648, n_312, n_476, n_818, n_429, n_861, n_534, n_948, n_884, n_899, n_345, n_210, n_944, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_1059, n_176, n_970, n_911, n_557, n_182, n_143, n_83, n_1005, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_857, n_560, n_656, n_340, n_207, n_561, n_1044, n_37, n_346, n_937, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_879, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_863, n_910, n_971, n_490, n_805, n_1027, n_117, n_326, n_794, n_768, n_921, n_996, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_1042, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_895, n_1037, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_1038, n_1025, n_887, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_870, n_931, n_159, n_334, n_599, n_766, n_811, n_952, n_541, n_807, n_391, n_701, n_434, n_1023, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_868, n_238, n_639, n_799, n_914, n_99, n_687, n_715, n_411, n_414, n_1026, n_319, n_364, n_965, n_927, n_20, n_536, n_531, n_935, n_1004, n_121, n_242, n_817, n_872, n_360, n_36, n_594, n_764, n_200, n_890, n_1056, n_162, n_960, n_64, n_759, n_1018, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_1011, n_904, n_985, n_1047, n_869, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_1029, n_166, n_626, n_11, n_925, n_424, n_1003, n_7, n_706, n_746, n_256, n_305, n_533, n_950, n_747, n_52, n_278, n_784, n_110, n_4802);

input n_137;
input n_924;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_977;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_1060;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_855;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_865;
input n_61;
input n_913;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_967;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_928;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_1055;
input n_916;
input n_452;
input n_885;
input n_397;
input n_493;
input n_111;
input n_525;
input n_880;
input n_703;
input n_698;
input n_980;
input n_483;
input n_544;
input n_683;
input n_1007;
input n_155;
input n_780;
input n_649;
input n_552;
input n_1057;
input n_1051;
input n_547;
input n_43;
input n_721;
input n_998;
input n_116;
input n_841;
input n_1050;
input n_956;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_983;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_1021;
input n_590;
input n_629;
input n_672;
input n_4;
input n_873;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_898;
input n_254;
input n_690;
input n_33;
input n_1013;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_1022;
input n_526;
input n_915;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_859;
input n_864;
input n_951;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_909;
input n_625;
input n_854;
input n_949;
input n_621;
input n_753;
input n_997;
input n_100;
input n_455;
input n_674;
input n_1008;
input n_932;
input n_417;
input n_946;
input n_1048;
input n_612;
input n_1001;
input n_212;
input n_385;
input n_498;
input n_516;
input n_933;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_912;
input n_606;
input n_559;
input n_275;
input n_640;
input n_968;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_1010;
input n_330;
input n_877;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_972;
input n_692;
input n_986;
input n_755;
input n_6;
input n_509;
input n_568;
input n_936;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_947;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_1024;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_999;
input n_668;
input n_733;
input n_991;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_941;
input n_929;
input n_981;
input n_1032;
input n_68;
input n_804;
input n_93;
input n_867;
input n_186;
input n_537;
input n_134;
input n_902;
input n_191;
input n_587;
input n_945;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_878;
input n_524;
input n_943;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_992;
input n_1049;
input n_938;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_984;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_883;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_905;
input n_906;
input n_24;
input n_406;
input n_519;
input n_470;
input n_908;
input n_782;
input n_919;
input n_325;
input n_449;
input n_132;
input n_862;
input n_90;
input n_900;
input n_724;
input n_856;
input n_546;
input n_1016;
input n_101;
input n_760;
input n_658;
input n_281;
input n_918;
input n_240;
input n_942;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_959;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_940;
input n_896;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_920;
input n_894;
input n_1046;
input n_271;
input n_934;
input n_1017;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_886;
input n_978;
input n_964;
input n_1054;
input n_654;
input n_370;
input n_167;
input n_976;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_1045;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_1033;
input n_988;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_1009;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_961;
input n_995;
input n_955;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_882;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_1036;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_1020;
input n_646;
input n_1062;
input n_211;
input n_218;
input n_400;
input n_930;
input n_181;
input n_436;
input n_962;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_1040;
input n_723;
input n_1035;
input n_386;
input n_578;
input n_994;
input n_926;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_1030;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_1043;
input n_496;
input n_355;
input n_958;
input n_849;
input n_1034;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_922;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_974;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_901;
input n_311;
input n_813;
input n_957;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_888;
input n_296;
input n_613;
input n_871;
input n_241;
input n_637;
input n_357;
input n_875;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_772;
input n_691;
input n_881;
input n_717;
input n_165;
input n_468;
input n_499;
input n_939;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_866;
input n_969;
input n_236;
input n_388;
input n_761;
input n_1012;
input n_1;
input n_1019;
input n_249;
input n_903;
input n_1006;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_889;
input n_80;
input n_973;
input n_35;
input n_73;
input n_277;
input n_1061;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_990;
input n_84;
input n_462;
input n_975;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_907;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_1031;
input n_263;
input n_471;
input n_609;
input n_852;
input n_989;
input n_1041;
input n_1039;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_1028;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_892;
input n_893;
input n_1015;
input n_1000;
input n_891;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_979;
input n_1002;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_874;
input n_465;
input n_838;
input n_76;
input n_358;
input n_1058;
input n_362;
input n_876;
input n_170;
input n_332;
input n_27;
input n_1053;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_953;
input n_601;
input n_279;
input n_917;
input n_1014;
input n_966;
input n_70;
input n_987;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_993;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_982;
input n_441;
input n_860;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_861;
input n_534;
input n_948;
input n_884;
input n_899;
input n_345;
input n_210;
input n_944;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_1059;
input n_176;
input n_970;
input n_911;
input n_557;
input n_182;
input n_143;
input n_83;
input n_1005;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_857;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_1044;
input n_37;
input n_346;
input n_937;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_879;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_863;
input n_910;
input n_971;
input n_490;
input n_805;
input n_1027;
input n_117;
input n_326;
input n_794;
input n_768;
input n_921;
input n_996;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_1042;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_895;
input n_1037;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_1038;
input n_1025;
input n_887;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_870;
input n_931;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_952;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_1023;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_868;
input n_238;
input n_639;
input n_799;
input n_914;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_1026;
input n_319;
input n_364;
input n_965;
input n_927;
input n_20;
input n_536;
input n_531;
input n_935;
input n_1004;
input n_121;
input n_242;
input n_817;
input n_872;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_890;
input n_1056;
input n_162;
input n_960;
input n_64;
input n_759;
input n_1018;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_1011;
input n_904;
input n_985;
input n_1047;
input n_869;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_1029;
input n_166;
input n_626;
input n_11;
input n_925;
input n_424;
input n_1003;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_950;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_4802;

wire n_1263;
wire n_3304;
wire n_1378;
wire n_2417;
wire n_2253;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_4706;
wire n_2739;
wire n_2380;
wire n_1166;
wire n_1751;
wire n_2771;
wire n_3241;
wire n_1508;
wire n_4129;
wire n_4604;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_4798;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_4419;
wire n_2746;
wire n_1677;
wire n_4477;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_3256;
wire n_3732;
wire n_1780;
wire n_1488;
wire n_4250;
wire n_2899;
wire n_2955;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4699;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_1370;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_4577;
wire n_4240;
wire n_4508;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_4639;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_2487;
wire n_1695;
wire n_3766;
wire n_1353;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_3813;
wire n_1535;
wire n_1789;
wire n_3350;
wire n_1666;
wire n_2389;
wire n_4165;
wire n_4238;
wire n_1451;
wire n_4038;
wire n_4109;
wire n_2302;
wire n_2374;
wire n_1545;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_4412;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_1462;
wire n_2069;
wire n_2396;
wire n_1799;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_4013;
wire n_2011;
wire n_2096;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_4780;
wire n_3163;
wire n_4425;
wire n_1118;
wire n_1686;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_2543;
wire n_1860;
wire n_4155;
wire n_1359;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_3695;
wire n_2482;
wire n_3891;
wire n_1728;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4131;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_4561;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_4548;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_4501;
wire n_3937;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_4525;
wire n_4622;
wire n_1243;
wire n_4315;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_3277;
wire n_1280;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_4499;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_2091;
wire n_2652;
wire n_2466;
wire n_2635;
wire n_1517;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_4691;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_1449;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_4483;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1484;
wire n_1328;
wire n_1374;
wire n_4715;
wire n_4793;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_3049;
wire n_1598;
wire n_4394;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_2384;
wire n_4485;
wire n_4626;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_4468;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1070;
wire n_1547;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_3985;
wire n_1801;
wire n_1391;
wire n_4615;
wire n_4760;
wire n_4652;
wire n_3361;
wire n_2908;
wire n_2970;
wire n_1513;
wire n_1600;
wire n_4624;
wire n_4758;
wire n_3744;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_2551;
wire n_1796;
wire n_3291;
wire n_4255;
wire n_4716;
wire n_1587;
wire n_2682;
wire n_1473;
wire n_3755;
wire n_4484;
wire n_2432;
wire n_3668;
wire n_4258;
wire n_1521;
wire n_4498;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_4745;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_4569;
wire n_2506;
wire n_2699;
wire n_4064;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_3550;
wire n_1626;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_2118;
wire n_2985;
wire n_1151;
wire n_2944;
wire n_4770;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_4629;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_4741;
wire n_1322;
wire n_2101;
wire n_1986;
wire n_1471;
wire n_2863;
wire n_4752;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_4552;
wire n_3252;
wire n_4421;
wire n_2275;
wire n_2855;
wire n_4503;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4464;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_3096;
wire n_2251;
wire n_1447;
wire n_1377;
wire n_3915;
wire n_4414;
wire n_2370;
wire n_3496;
wire n_4469;
wire n_3954;
wire n_4114;
wire n_2544;
wire n_4532;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3735;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_4067;
wire n_4674;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_4385;
wire n_3320;
wire n_4556;
wire n_3007;
wire n_2688;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_2622;
wire n_1278;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_1667;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_4504;
wire n_2241;
wire n_4717;
wire n_4788;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_3781;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_4531;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_4609;
wire n_2987;
wire n_2042;
wire n_1527;
wire n_4567;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_3328;
wire n_4130;
wire n_4234;
wire n_1754;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4471;
wire n_4161;
wire n_4472;
wire n_4462;
wire n_3433;
wire n_4024;
wire n_3392;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_2305;
wire n_3430;
wire n_3975;
wire n_4444;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_3331;
wire n_1319;
wire n_2379;
wire n_3447;
wire n_3992;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4148;
wire n_4151;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_4415;
wire n_1387;
wire n_4466;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4702;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_4457;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_4786;
wire n_1156;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_4160;
wire n_2945;
wire n_2331;
wire n_2798;
wire n_2293;
wire n_3989;
wire n_4475;
wire n_2837;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_2319;
wire n_1393;
wire n_3296;
wire n_2979;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2808;
wire n_3009;
wire n_1276;
wire n_2548;
wire n_1412;
wire n_2676;
wire n_2679;
wire n_1709;
wire n_3981;
wire n_4683;
wire n_2108;
wire n_3640;
wire n_4491;
wire n_4388;
wire n_1162;
wire n_2930;
wire n_1538;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_2434;
wire n_1884;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_2967;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_4647;
wire n_3923;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_4696;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_2454;
wire n_4371;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_2801;
wire n_3120;
wire n_1293;
wire n_4473;
wire n_1876;
wire n_4007;
wire n_1743;
wire n_4620;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_1175;
wire n_2763;
wire n_4613;
wire n_1479;
wire n_1810;
wire n_4480;
wire n_4649;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_3643;
wire n_2009;
wire n_1888;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_4438;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_3218;
wire n_3748;
wire n_1766;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_4795;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4623;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_4553;
wire n_3819;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_2491;
wire n_1788;
wire n_3747;
wire n_1537;
wire n_3833;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_4262;
wire n_2671;
wire n_4184;
wire n_4618;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2022;
wire n_1798;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_4585;
wire n_2876;
wire n_4720;
wire n_2629;
wire n_1415;
wire n_4099;
wire n_2592;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2838;
wire n_2181;
wire n_2479;
wire n_1647;
wire n_4340;
wire n_1829;
wire n_3513;
wire n_3133;
wire n_1464;
wire n_4295;
wire n_4685;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_4645;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_4490;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_4511;
wire n_2928;
wire n_3128;
wire n_4694;
wire n_1734;
wire n_4533;
wire n_3038;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_3068;
wire n_2871;
wire n_2178;
wire n_1308;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_4757;
wire n_4603;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_4648;
wire n_2469;
wire n_1333;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_4391;
wire n_4641;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_3855;
wire n_1539;
wire n_2736;
wire n_4283;
wire n_4157;
wire n_4681;
wire n_2054;
wire n_1503;
wire n_3765;
wire n_1468;
wire n_4638;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_3816;
wire n_2623;
wire n_1617;
wire n_1744;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_1279;
wire n_3108;
wire n_1406;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_3760;
wire n_2577;
wire n_1837;
wire n_4108;
wire n_4486;
wire n_4557;
wire n_4707;
wire n_4078;
wire n_4451;
wire n_1760;
wire n_2875;
wire n_2960;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_4527;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_4627;
wire n_1851;
wire n_4156;
wire n_3205;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_4787;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_4541;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_2580;
wire n_1871;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_3271;
wire n_4771;
wire n_2039;
wire n_1207;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_2084;
wire n_1781;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_4432;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_2459;
wire n_3031;
wire n_4692;
wire n_4154;
wire n_4619;
wire n_4673;
wire n_3396;
wire n_3701;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_4420;
wire n_3243;
wire n_1773;
wire n_1169;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1596;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_4299;
wire n_2314;
wire n_2116;
wire n_1434;
wire n_4801;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2320;
wire n_2339;
wire n_2473;
wire n_1208;
wire n_2038;
wire n_3287;
wire n_4637;
wire n_2137;
wire n_3378;
wire n_4640;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_3767;
wire n_4279;
wire n_4769;
wire n_4785;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_3820;
wire n_4367;
wire n_4589;
wire n_3741;
wire n_3410;
wire n_4578;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_4413;
wire n_3502;
wire n_2523;
wire n_3098;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_4387;
wire n_2312;
wire n_3990;
wire n_4493;
wire n_4790;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4453;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_2536;
wire n_1592;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_2338;
wire n_1758;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_2725;
wire n_1548;
wire n_1421;
wire n_4510;
wire n_4610;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_4489;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_4570;
wire n_4542;
wire n_1119;
wire n_2261;
wire n_2156;
wire n_2729;
wire n_1240;
wire n_3268;
wire n_1820;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_4281;
wire n_2519;
wire n_3354;
wire n_4661;
wire n_2724;
wire n_4447;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_2897;
wire n_2077;
wire n_3614;
wire n_1416;
wire n_4198;
wire n_2909;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_1724;
wire n_4285;
wire n_4651;
wire n_3466;
wire n_4534;
wire n_4500;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_4514;
wire n_1366;
wire n_4606;
wire n_4800;
wire n_1300;
wire n_3960;
wire n_4774;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_4597;
wire n_3905;
wire n_4329;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_3200;
wire n_1664;
wire n_4271;
wire n_1486;
wire n_3586;
wire n_4672;
wire n_1332;
wire n_3519;
wire n_4433;
wire n_2231;
wire n_1390;
wire n_4682;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_4766;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_4460;
wire n_2400;
wire n_4633;
wire n_3645;
wire n_4614;
wire n_3838;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3929;
wire n_3077;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_4732;
wire n_2272;
wire n_3984;
wire n_1140;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_4665;
wire n_1913;
wire n_2878;
wire n_4693;
wire n_1823;
wire n_4434;
wire n_4662;
wire n_3679;
wire n_3779;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4744;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_4545;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_2490;
wire n_1903;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_3154;
wire n_1551;
wire n_3229;
wire n_4213;
wire n_4463;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_3692;
wire n_1816;
wire n_4687;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_4595;
wire n_1849;
wire n_3788;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_2410;
wire n_1131;
wire n_4313;
wire n_1084;
wire n_1961;
wire n_4037;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_2240;
wire n_2696;
wire n_1351;
wire n_4063;
wire n_4428;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_4650;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3995;
wire n_4669;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_4339;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4583;
wire n_4060;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_4763;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_4594;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_4666;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_2555;
wire n_1381;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_4015;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_4494;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_4714;
wire n_3465;
wire n_1316;
wire n_2419;
wire n_3215;
wire n_1708;
wire n_4796;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_3961;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_1630;
wire n_4540;
wire n_4102;
wire n_4776;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_4799;
wire n_1437;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_1092;
wire n_2694;
wire n_3559;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_4775;
wire n_3993;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_3462;
wire n_3588;
wire n_1424;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_4590;
wire n_2910;
wire n_1893;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_4455;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_4664;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_2969;
wire n_2191;
wire n_2864;
wire n_1311;
wire n_3941;
wire n_4754;
wire n_3195;
wire n_3190;
wire n_1519;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_4443;
wire n_3847;
wire n_2664;
wire n_4507;
wire n_4554;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_4575;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_4663;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3569;
wire n_3548;
wire n_4348;
wire n_4452;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_3953;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_3110;
wire n_1632;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_4572;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_4608;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_4104;
wire n_4512;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_4784;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4791;
wire n_4384;
wire n_4536;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_4521;
wire n_4488;
wire n_2086;
wire n_3537;
wire n_4423;
wire n_4773;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_4497;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_4611;
wire n_1763;
wire n_4755;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_4588;
wire n_2475;
wire n_2733;
wire n_2993;
wire n_1719;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_4598;
wire n_4478;
wire n_2785;
wire n_4658;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2415;
wire n_2309;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_4519;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_4470;
wire n_2816;
wire n_1228;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_4422;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_2903;
wire n_3482;
wire n_3417;
wire n_3866;
wire n_1967;
wire n_3921;
wire n_1143;
wire n_2233;
wire n_1579;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_4555;
wire n_2827;
wire n_3052;
wire n_1688;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_3326;
wire n_4689;
wire n_3956;
wire n_3572;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4721;
wire n_4047;
wire n_3734;
wire n_3237;
wire n_2082;
wire n_4778;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_4550;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_4441;
wire n_4496;
wire n_4761;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1557;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_3196;
wire n_1422;
wire n_4095;
wire n_3078;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_4727;
wire n_3952;
wire n_4568;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_4599;
wire n_3633;
wire n_3363;
wire n_4479;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_1735;
wire n_1697;
wire n_2020;
wire n_4628;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_4495;
wire n_4762;
wire n_1881;
wire n_4416;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2751;
wire n_2793;
wire n_2707;
wire n_3372;
wire n_3451;
wire n_4539;
wire n_2971;
wire n_4657;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_4458;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_2285;
wire n_1446;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_2471;
wire n_2298;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_4476;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_3342;
wire n_4748;
wire n_2303;
wire n_1824;
wire n_2295;
wire n_1917;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_4667;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_4690;
wire n_1814;
wire n_2822;
wire n_4437;
wire n_4710;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_4607;
wire n_2126;
wire n_4547;
wire n_4117;
wire n_2893;
wire n_4573;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_4668;
wire n_2600;
wire n_4487;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_2795;
wire n_4091;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3460;
wire n_3409;
wire n_2352;
wire n_4759;
wire n_3538;
wire n_1413;
wire n_4040;
wire n_2207;
wire n_4467;
wire n_2080;
wire n_2619;
wire n_2377;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_1110;
wire n_4474;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_3123;
wire n_1895;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_4728;
wire n_4316;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_4247;
wire n_2638;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4617;
wire n_4062;
wire n_4524;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1998;
wire n_1105;
wire n_4686;
wire n_4518;
wire n_3759;
wire n_1338;
wire n_4409;
wire n_4411;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_2034;
wire n_1637;
wire n_1687;
wire n_2711;
wire n_1419;
wire n_4631;
wire n_4336;
wire n_3933;
wire n_2270;
wire n_1653;
wire n_1506;
wire n_3206;
wire n_4777;
wire n_4792;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_2794;
wire n_2259;
wire n_1256;
wire n_1702;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_1122;
wire n_4068;
wire n_4290;
wire n_4253;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_4709;
wire n_2995;
wire n_2494;
wire n_1375;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_4398;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1929;
wire n_1392;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_1834;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_3324;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_4625;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_4431;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_3736;
wire n_4656;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_4729;
wire n_1116;
wire n_2000;
wire n_3402;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4679;
wire n_4115;
wire n_3174;
wire n_4701;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_2217;
wire n_1453;
wire n_3746;
wire n_1731;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_2722;
wire n_1658;
wire n_2201;
wire n_1737;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_3835;
wire n_3432;
wire n_2493;
wire n_2205;
wire n_1628;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_4537;
wire n_3090;
wire n_2067;
wire n_2437;
wire n_1168;
wire n_2219;
wire n_3762;
wire n_2885;
wire n_3902;
wire n_4730;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_3654;
wire n_3839;
wire n_3035;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_4659;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_3972;
wire n_4616;
wire n_4579;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_3358;
wire n_2605;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_4747;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1991;
wire n_2224;
wire n_1543;
wire n_1979;
wire n_3368;
wire n_1533;
wire n_1399;
wire n_2924;
wire n_4772;
wire n_3467;
wire n_2484;
wire n_4111;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_4587;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_4743;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_4538;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_3928;
wire n_4653;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_4654;
wire n_2264;
wire n_4677;
wire n_2754;
wire n_3534;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_4632;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_3438;
wire n_4098;
wire n_2012;
wire n_3792;
wire n_4733;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_2245;
wire n_3561;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_4789;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_2806;
wire n_1485;
wire n_4269;
wire n_2184;
wire n_1184;
wire n_4695;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_2965;
wire n_3661;
wire n_1855;
wire n_4150;
wire n_3635;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_2926;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_2213;
wire n_2023;
wire n_1170;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_4442;
wire n_3968;
wire n_4698;
wire n_4634;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_4704;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_2697;
wire n_1461;
wire n_4551;
wire n_3074;
wire n_3204;
wire n_4779;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_2861;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_4781;
wire n_2977;
wire n_3606;
wire n_4738;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_4424;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_4700;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_4426;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2284;
wire n_2187;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_4436;
wire n_3878;
wire n_1762;
wire n_4450;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_4601;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_4746;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_1890;
wire n_4220;
wire n_4251;
wire n_1817;
wire n_1944;
wire n_1683;
wire n_1497;
wire n_1530;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_3431;
wire n_4621;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_4737;
wire n_3070;
wire n_3284;
wire n_1326;
wire n_4066;
wire n_3647;
wire n_4459;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_4515;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_4559;
wire n_4403;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_4368;
wire n_1663;
wire n_1718;
wire n_4050;
wire n_4509;
wire n_3700;
wire n_4740;
wire n_3609;
wire n_4136;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_4642;
wire n_4393;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_4535;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_2326;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_4522;
wire n_2188;
wire n_4794;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_4724;
wire n_4644;
wire n_4456;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_4520;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_1861;
wire n_4546;
wire n_3584;
wire n_1425;
wire n_4592;
wire n_3858;
wire n_4675;
wire n_1901;
wire n_3069;
wire n_4502;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1727;
wire n_1554;
wire n_4382;
wire n_4435;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_4571;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_2447;
wire n_3761;
wire n_1813;
wire n_4764;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4723;
wire n_2382;
wire n_4719;
wire n_1707;
wire n_4178;
wire n_4655;
wire n_3062;
wire n_3161;
wire n_4581;
wire n_2317;
wire n_3289;
wire n_4558;
wire n_2799;
wire n_4454;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_1083;
wire n_1142;
wire n_4739;
wire n_2376;
wire n_2488;
wire n_4722;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_4768;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_2250;
wire n_2678;
wire n_2778;
wire n_1756;
wire n_4782;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_2451;
wire n_1520;
wire n_2887;
wire n_4363;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_1550;
wire n_4465;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_4605;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_3842;
wire n_3050;
wire n_3265;
wire n_1536;
wire n_1857;
wire n_4056;
wire n_4482;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_2957;
wire n_3551;
wire n_3903;
wire n_1769;
wire n_4783;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_3314;
wire n_4158;
wire n_4530;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_2173;
wire n_1250;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_1585;
wire n_3245;
wire n_4417;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_3527;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_2030;
wire n_1348;
wire n_2453;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_1525;
wire n_1752;
wire n_4287;
wire n_4749;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_4516;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_4270;
wire n_4505;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_4574;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_3497;
wire n_4602;
wire n_1487;
wire n_4449;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_4750;
wire n_1495;
wire n_1337;
wire n_4445;
wire n_4566;
wire n_4231;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3322;
wire n_3232;
wire n_4576;
wire n_3652;
wire n_1245;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1975;
wire n_1321;
wire n_4061;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_4083;
wire n_2112;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3125;
wire n_2594;
wire n_3114;
wire n_3234;
wire n_2394;
wire n_1914;
wire n_3612;
wire n_4461;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_4430;
wire n_2381;
wire n_4767;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_4407;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4676;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_4544;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_4429;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_4591;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_4646;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4446;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_4797;
wire n_2366;
wire n_4563;
wire n_4725;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_1275;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_2820;
wire n_1402;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4320;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_4596;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_4492;
wire n_2708;
wire n_3809;
wire n_1621;
wire n_2113;
wire n_3694;
wire n_2586;
wire n_1448;
wire n_4288;
wire n_4245;
wire n_4364;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_4378;
wire n_4726;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_1879;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_4751;
wire n_1181;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_4636;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_1558;
wire n_4584;
wire n_4241;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_4711;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_4309;
wire n_2256;
wire n_3152;
wire n_1704;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_4680;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_1186;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_4560;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_4671;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_3693;
wire n_1542;
wire n_1251;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_4705;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;
wire n_4580;

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_983),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_942),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_954),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_37),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_13),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_945),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_0),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_498),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_959),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_427),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_510),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_823),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_725),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_545),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_85),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_358),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_946),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_464),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_979),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_350),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_700),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_101),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_980),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_444),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_943),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_231),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_641),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_991),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_97),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_56),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_169),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_956),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_851),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_860),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_875),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_334),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_660),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_330),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_40),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_621),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_128),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_160),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_376),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_39),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_704),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_952),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_360),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_689),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_93),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_554),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_927),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_990),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_802),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_447),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_380),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_520),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_221),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_700),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_788),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_123),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_486),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_862),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_368),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1058),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_907),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_119),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_143),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_670),
.Y(n_1130)
);

CKINVDCx16_ASAP7_75t_R g1131 ( 
.A(n_947),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_394),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_940),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_869),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_266),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_358),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1015),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_348),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_972),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_262),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_216),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_123),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_489),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_993),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_918),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_269),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_182),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_924),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_832),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_862),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_992),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_276),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_929),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_220),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_828),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_279),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_170),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1017),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_462),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_21),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_39),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_92),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_645),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_994),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_855),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_71),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_135),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_268),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_922),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_469),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_53),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1006),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_165),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_4),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_247),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_521),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_968),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_971),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_553),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_88),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_587),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_158),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_613),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_96),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1057),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_130),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_647),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_767),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_883),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_439),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_386),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_430),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_384),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_488),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_580),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_793),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_739),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_321),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_964),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_866),
.Y(n_1200)
);

CKINVDCx12_ASAP7_75t_R g1201 ( 
.A(n_15),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_136),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_129),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_140),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_302),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_625),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_185),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_773),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_663),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_595),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_143),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_984),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_814),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_788),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_434),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_164),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_417),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_544),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_884),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_97),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_352),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_492),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_594),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_58),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_894),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_768),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_472),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_353),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_993),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_73),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_977),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_540),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_549),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_607),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_487),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_119),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_848),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_718),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_995),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_176),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_885),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_726),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_79),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_229),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_477),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_663),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_450),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_963),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_944),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_880),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_205),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_381),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_19),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_331),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_369),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_189),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_523),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_556),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_530),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_850),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_116),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_268),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_947),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_941),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_867),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_916),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_238),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_966),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_410),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_199),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_898),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_602),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_363),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_935),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_233),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_571),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_709),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_231),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_343),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_77),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_479),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_925),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_798),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_683),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_419),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_999),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_647),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_837),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_807),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_156),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_244),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_773),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_14),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_82),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_486),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_5),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_438),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_46),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1010),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_29),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_378),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_775),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_921),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_900),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_754),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_811),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_892),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_658),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_691),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_485),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_887),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_821),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_140),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1047),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_798),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_908),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_360),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_437),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_350),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_60),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_795),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_954),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1003),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_449),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_193),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_213),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_505),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_817),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_79),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_952),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_262),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_955),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_380),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_90),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_299),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_909),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_990),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_523),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_215),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_688),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_864),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_14),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_434),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_845),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_745),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_168),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_62),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_978),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_939),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_372),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_771),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_258),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_728),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_806),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_321),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_166),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1005),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_560),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_981),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_820),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_65),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_483),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_242),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_363),
.Y(n_1365)
);

BUFx10_ASAP7_75t_L g1366 ( 
.A(n_261),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_508),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1041),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_677),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_236),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_543),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_836),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1060),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_594),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_422),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_969),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_866),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_420),
.Y(n_1378)
);

CKINVDCx14_ASAP7_75t_R g1379 ( 
.A(n_898),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_357),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1001),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_929),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_840),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_392),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_730),
.Y(n_1385)
);

CKINVDCx16_ASAP7_75t_R g1386 ( 
.A(n_846),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_893),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_712),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_248),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_521),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_692),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_438),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_894),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_401),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_529),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_138),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_901),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_25),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_849),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_451),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_391),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_469),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_874),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_988),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_235),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_695),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_914),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_178),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_853),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_926),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_790),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_619),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_37),
.Y(n_1413)
);

BUFx5_ASAP7_75t_L g1414 ( 
.A(n_578),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1010),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_937),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_25),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_302),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1000),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_42),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_320),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_960),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_355),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_456),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_986),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_753),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_882),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_216),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_602),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_219),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_601),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_592),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_290),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_743),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_948),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_14),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_889),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_846),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_979),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_887),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_291),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_910),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_856),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_392),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_550),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_597),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_835),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_156),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1036),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1017),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_685),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_914),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_895),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_951),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_542),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_201),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_933),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_28),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_987),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_876),
.Y(n_1461)
);

CKINVDCx16_ASAP7_75t_R g1462 ( 
.A(n_813),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_675),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1046),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1062),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_28),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_941),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_985),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_149),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_897),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_389),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_774),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_366),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_472),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_868),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_185),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_855),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1056),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_271),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_343),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_718),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_930),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_902),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_890),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_80),
.Y(n_1485)
);

BUFx5_ASAP7_75t_L g1486 ( 
.A(n_531),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_720),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_705),
.Y(n_1488)
);

CKINVDCx14_ASAP7_75t_R g1489 ( 
.A(n_349),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_915),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_545),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_917),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_720),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_985),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_353),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_580),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_907),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_495),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_32),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_800),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_170),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_776),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_316),
.Y(n_1503)
);

BUFx10_ASAP7_75t_L g1504 ( 
.A(n_1030),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_957),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_646),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_11),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_842),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_870),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_121),
.Y(n_1510)
);

BUFx10_ASAP7_75t_L g1511 ( 
.A(n_355),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_879),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_316),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_751),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_899),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_557),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_398),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_672),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_346),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_689),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_141),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_42),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_43),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_198),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_429),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_260),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_419),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_325),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_383),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_888),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1046),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_716),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_36),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_630),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_286),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_137),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1054),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1029),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_982),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_628),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_923),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_853),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_374),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_909),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_47),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_856),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_655),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_950),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_137),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_286),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_590),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_181),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_844),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_332),
.Y(n_1554)
);

BUFx8_ASAP7_75t_SL g1555 ( 
.A(n_157),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_944),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_341),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_886),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_31),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_125),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_55),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_891),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_742),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_98),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_198),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_873),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_408),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_895),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_807),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_163),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_197),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_764),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_515),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_739),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_656),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_740),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_13),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_588),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_624),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_843),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_859),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_512),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_698),
.Y(n_1583)
);

INVx4_ASAP7_75t_R g1584 ( 
.A(n_841),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_683),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_975),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_479),
.Y(n_1587)
);

CKINVDCx14_ASAP7_75t_R g1588 ( 
.A(n_975),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_557),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_871),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_977),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_440),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_481),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_994),
.Y(n_1594)
);

CKINVDCx16_ASAP7_75t_R g1595 ( 
.A(n_719),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_640),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_627),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1058),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_847),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_881),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_649),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_620),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_681),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_17),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_299),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_378),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_219),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_676),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_931),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_447),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_385),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_473),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_369),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_120),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_109),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_202),
.Y(n_1616)
);

BUFx5_ASAP7_75t_L g1617 ( 
.A(n_974),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_637),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_183),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_695),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_217),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_938),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_305),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_404),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_583),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_401),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1029),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_430),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_865),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_487),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_90),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_461),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_964),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_159),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_674),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_613),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_920),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_595),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_608),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_252),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_997),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_901),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_631),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_676),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_93),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_806),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_931),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_240),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_714),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_324),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_494),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_300),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_490),
.Y(n_1653)
);

BUFx10_ASAP7_75t_L g1654 ( 
.A(n_921),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_617),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_741),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_351),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_970),
.Y(n_1658)
);

BUFx10_ASAP7_75t_L g1659 ( 
.A(n_18),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_858),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_519),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_276),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_796),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1049),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_854),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_181),
.Y(n_1666)
);

BUFx10_ASAP7_75t_L g1667 ( 
.A(n_869),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_872),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_478),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1038),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_120),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_387),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_936),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_320),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_607),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_312),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1040),
.Y(n_1677)
);

BUFx10_ASAP7_75t_L g1678 ( 
.A(n_1035),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1000),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1008),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_145),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_511),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_168),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_517),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_224),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_265),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_193),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_519),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_657),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_383),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_912),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_159),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_732),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_692),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_893),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_127),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_367),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_511),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_905),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_803),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_374),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_381),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_483),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_514),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_906),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_879),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_845),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_969),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_601),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_520),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_217),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_556),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_395),
.Y(n_1713)
);

CKINVDCx20_ASAP7_75t_R g1714 ( 
.A(n_951),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_904),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_421),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_517),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_989),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_885),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_138),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_750),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_976),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_292),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_971),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_970),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_813),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_50),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_912),
.Y(n_1728)
);

CKINVDCx20_ASAP7_75t_R g1729 ( 
.A(n_45),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_183),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_584),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_781),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_105),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_263),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_616),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_228),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_624),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_932),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_214),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_311),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_868),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_70),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_965),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_102),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_23),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_347),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_690),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_643),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_923),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1049),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_878),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_339),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_284),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_340),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_934),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_395),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_182),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_510),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_956),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_31),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_292),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_668),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_861),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_76),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_945),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_289),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1043),
.Y(n_1767)
);

BUFx8_ASAP7_75t_SL g1768 ( 
.A(n_1050),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_420),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_645),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_377),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_527),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_592),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_49),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_118),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_611),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_777),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_410),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_934),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_967),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_505),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_573),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_911),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_439),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_107),
.Y(n_1785)
);

BUFx10_ASAP7_75t_L g1786 ( 
.A(n_641),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_961),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_878),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_778),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1003),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_408),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_394),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_753),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_303),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_953),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_863),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_41),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_352),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_118),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_273),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_704),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_2),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_266),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_368),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_567),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_999),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_539),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_877),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_717),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_86),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_759),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_73),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_175),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_145),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_284),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_802),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_62),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_508),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_770),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_808),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_882),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_614),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_59),
.Y(n_1823)
);

CKINVDCx20_ASAP7_75t_R g1824 ( 
.A(n_13),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_903),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_155),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_354),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_128),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1055),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_356),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_393),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_264),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_27),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_494),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1026),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_913),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_617),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_89),
.Y(n_1838)
);

BUFx2_ASAP7_75t_SL g1839 ( 
.A(n_200),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_658),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_83),
.Y(n_1841)
);

CKINVDCx12_ASAP7_75t_R g1842 ( 
.A(n_949),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_697),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_633),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_896),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_375),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_370),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_682),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_867),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_160),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_748),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_206),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_728),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_715),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_857),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_537),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_397),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_110),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_165),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_226),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_962),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_484),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_297),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_225),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_34),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_190),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_192),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_329),
.Y(n_1868)
);

INVxp33_ASAP7_75t_SL g1869 ( 
.A(n_732),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_768),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_957),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_634),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_698),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_777),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_324),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_967),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_852),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_800),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_474),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_15),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_797),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1033),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_480),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_767),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_341),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_577),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_414),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_919),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_714),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_375),
.Y(n_1890)
);

CKINVDCx20_ASAP7_75t_R g1891 ( 
.A(n_631),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_628),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_880),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_196),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_973),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1024),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_482),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_124),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_699),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_148),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_544),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_958),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_716),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_187),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_245),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_991),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_471),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_179),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_87),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_618),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_45),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_463),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_502),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_4),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_75),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_928),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_465),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1414),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1379),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1414),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1414),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1414),
.Y(n_1922)
);

INVxp33_ASAP7_75t_L g1923 ( 
.A(n_1306),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1414),
.Y(n_1924)
);

INVxp33_ASAP7_75t_SL g1925 ( 
.A(n_1066),
.Y(n_1925)
);

INVxp33_ASAP7_75t_SL g1926 ( 
.A(n_1066),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1378),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1414),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1489),
.Y(n_1929)
);

INVxp33_ASAP7_75t_SL g1930 ( 
.A(n_1160),
.Y(n_1930)
);

INVxp33_ASAP7_75t_SL g1931 ( 
.A(n_1160),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1414),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1486),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1486),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1486),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1486),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1127),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1555),
.Y(n_1938)
);

INVxp33_ASAP7_75t_SL g1939 ( 
.A(n_1161),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1486),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1486),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1588),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1486),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1100),
.Y(n_1944)
);

CKINVDCx16_ASAP7_75t_R g1945 ( 
.A(n_1522),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1617),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1131),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1617),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1617),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1768),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1617),
.Y(n_1951)
);

INVxp67_ASAP7_75t_SL g1952 ( 
.A(n_1174),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1675),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1617),
.Y(n_1954)
);

INVx4_ASAP7_75t_R g1955 ( 
.A(n_1185),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1444),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1617),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1617),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1248),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1132),
.Y(n_1960)
);

CKINVDCx20_ASAP7_75t_R g1961 ( 
.A(n_1386),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1257),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1174),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1659),
.Y(n_1964)
);

INVxp67_ASAP7_75t_SL g1965 ( 
.A(n_1174),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1174),
.Y(n_1966)
);

CKINVDCx20_ASAP7_75t_R g1967 ( 
.A(n_1456),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1436),
.Y(n_1968)
);

NOR2xp67_ASAP7_75t_L g1969 ( 
.A(n_1315),
.B(n_0),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1436),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1297),
.Y(n_1971)
);

INVxp33_ASAP7_75t_SL g1972 ( 
.A(n_1161),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1436),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1436),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1315),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1301),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1315),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1398),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1420),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1459),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1499),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1523),
.Y(n_1982)
);

CKINVDCx14_ASAP7_75t_R g1983 ( 
.A(n_1659),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1533),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1745),
.Y(n_1985)
);

INVx1_ASAP7_75t_SL g1986 ( 
.A(n_1483),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1462),
.Y(n_1987)
);

INVxp67_ASAP7_75t_SL g1988 ( 
.A(n_1791),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1301),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1760),
.Y(n_1990)
);

INVxp33_ASAP7_75t_L g1991 ( 
.A(n_1858),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1201),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1595),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1132),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1302),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1302),
.Y(n_1996)
);

INVxp33_ASAP7_75t_SL g1997 ( 
.A(n_1880),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1842),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1494),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1880),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1559),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1914),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1494),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1559),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1779),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1544),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1544),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1132),
.Y(n_2008)
);

INVxp33_ASAP7_75t_L g2009 ( 
.A(n_1889),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1570),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1570),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1634),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1634),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1711),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1132),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1711),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1723),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1723),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1870),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1638),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1870),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1162),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1162),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1162),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1162),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1226),
.Y(n_2026)
);

CKINVDCx20_ASAP7_75t_R g2027 ( 
.A(n_1064),
.Y(n_2027)
);

CKINVDCx20_ASAP7_75t_R g2028 ( 
.A(n_1064),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1226),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1226),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1226),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1234),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1079),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1234),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1067),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1234),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1069),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1234),
.Y(n_2038)
);

CKINVDCx14_ASAP7_75t_R g2039 ( 
.A(n_1659),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1284),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1284),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1284),
.Y(n_2042)
);

CKINVDCx20_ASAP7_75t_R g2043 ( 
.A(n_1079),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1284),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1101),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_1552),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_1128),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1552),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_1081),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1552),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1552),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1914),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1564),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1564),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1253),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1081),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1564),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1564),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1739),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1739),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1739),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1087),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1294),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1087),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1739),
.Y(n_2065)
);

CKINVDCx20_ASAP7_75t_R g2066 ( 
.A(n_1094),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1784),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1343),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1784),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1784),
.Y(n_2070)
);

INVxp33_ASAP7_75t_SL g2071 ( 
.A(n_1413),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1128),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1784),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1825),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1825),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_1450),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1825),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1825),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1912),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1913),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1094),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1068),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_1185),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_1417),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1103),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1073),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1075),
.Y(n_2087)
);

INVxp67_ASAP7_75t_SL g2088 ( 
.A(n_1138),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1901),
.Y(n_2089)
);

INVxp33_ASAP7_75t_SL g2090 ( 
.A(n_1466),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_1103),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1507),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1077),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1577),
.Y(n_2094)
);

CKINVDCx20_ASAP7_75t_R g2095 ( 
.A(n_1112),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_1144),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1085),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1604),
.Y(n_2098)
);

BUFx2_ASAP7_75t_SL g2099 ( 
.A(n_1128),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_1112),
.Y(n_2100)
);

CKINVDCx16_ASAP7_75t_R g2101 ( 
.A(n_1200),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1086),
.Y(n_2102)
);

CKINVDCx20_ASAP7_75t_R g2103 ( 
.A(n_1130),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1089),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1091),
.Y(n_2105)
);

INVxp33_ASAP7_75t_SL g2106 ( 
.A(n_1797),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1900),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1902),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1093),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1096),
.Y(n_2110)
);

INVxp33_ASAP7_75t_SL g2111 ( 
.A(n_1802),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1102),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1200),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_2067),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1952),
.B(n_1197),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_1956),
.A2(n_1833),
.B1(n_1582),
.B2(n_1698),
.Y(n_2116)
);

CKINVDCx6p67_ASAP7_75t_R g2117 ( 
.A(n_1919),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2008),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_1976),
.Y(n_2119)
);

OA21x2_ASAP7_75t_L g2120 ( 
.A1(n_1975),
.A2(n_1147),
.B(n_1133),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2015),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2067),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1963),
.B(n_1965),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2034),
.Y(n_2124)
);

OAI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_1956),
.A2(n_1168),
.B1(n_1065),
.B2(n_1123),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_1989),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2053),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2067),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_1959),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1960),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1994),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1960),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2046),
.B(n_1197),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1966),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1968),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1938),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1970),
.Y(n_2137)
);

BUFx12f_ASAP7_75t_L g2138 ( 
.A(n_1950),
.Y(n_2138)
);

AND2x6_ASAP7_75t_L g2139 ( 
.A(n_1920),
.B(n_1133),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_2035),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2022),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1973),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1974),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1995),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1996),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1918),
.A2(n_1165),
.B(n_1147),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2023),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2024),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_SL g2149 ( 
.A1(n_1944),
.A2(n_1865),
.B1(n_1824),
.B2(n_1194),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2025),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2026),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2029),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2030),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2031),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2113),
.B(n_1964),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1962),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2032),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_2001),
.Y(n_2158)
);

AND2x2_ASAP7_75t_SL g2159 ( 
.A(n_1945),
.B(n_1165),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1999),
.B(n_1218),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1988),
.B(n_1370),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_2003),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2036),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2038),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2040),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_SL g2166 ( 
.A(n_1986),
.B(n_1130),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2088),
.B(n_1218),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2041),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1971),
.Y(n_2169)
);

OAI22x1_ASAP7_75t_L g2170 ( 
.A1(n_1986),
.A2(n_1953),
.B1(n_1927),
.B2(n_1937),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_2004),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2063),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2101),
.B(n_1200),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2042),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_1987),
.A2(n_1869),
.B1(n_1747),
.B2(n_1071),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_2087),
.Y(n_2176)
);

BUFx12f_ASAP7_75t_L g2177 ( 
.A(n_1993),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_2071),
.B(n_1869),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_2044),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2096),
.B(n_1244),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2020),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2037),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_2090),
.B(n_1244),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_2048),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2050),
.Y(n_2185)
);

INVx4_ASAP7_75t_L g2186 ( 
.A(n_2045),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2051),
.Y(n_2187)
);

BUFx3_ASAP7_75t_L g2188 ( 
.A(n_2006),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_2054),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2057),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2058),
.Y(n_2191)
);

OA21x2_ASAP7_75t_L g2192 ( 
.A1(n_1977),
.A2(n_1179),
.B(n_1177),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2007),
.B(n_1331),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_2059),
.Y(n_2194)
);

NAND2xp33_ASAP7_75t_L g2195 ( 
.A(n_2055),
.B(n_1063),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_1940),
.A2(n_1179),
.B(n_1177),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2060),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2010),
.B(n_1331),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_2068),
.B(n_1220),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_SL g2200 ( 
.A(n_1929),
.B(n_1194),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2061),
.Y(n_2201)
);

INVx5_ASAP7_75t_L g2202 ( 
.A(n_1949),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2084),
.B(n_1368),
.Y(n_2203)
);

INVx6_ASAP7_75t_L g2204 ( 
.A(n_2099),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_2092),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_2076),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2065),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_2069),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1958),
.A2(n_1266),
.B(n_1251),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_SL g2210 ( 
.A1(n_1947),
.A2(n_1865),
.B1(n_1824),
.B2(n_1225),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2070),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2073),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_1921),
.A2(n_1266),
.B(n_1251),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2074),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2005),
.B(n_1992),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2075),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2094),
.B(n_2098),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2011),
.B(n_1368),
.Y(n_2218)
);

AND3x1_ASAP7_75t_L g2219 ( 
.A(n_2000),
.B(n_1846),
.C(n_1268),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_2077),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2078),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1922),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_2106),
.B(n_1846),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2079),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1998),
.B(n_1108),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2080),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1924),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2082),
.Y(n_2228)
);

AOI22x1_ASAP7_75t_SL g2229 ( 
.A1(n_2027),
.A2(n_1225),
.B1(n_1239),
.B2(n_1198),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1978),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1983),
.B(n_1220),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2086),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2012),
.B(n_2013),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_1979),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_1980),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2014),
.B(n_1070),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1928),
.Y(n_2237)
);

INVx4_ASAP7_75t_L g2238 ( 
.A(n_1932),
.Y(n_2238)
);

CKINVDCx11_ASAP7_75t_R g2239 ( 
.A(n_2028),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2009),
.A2(n_1065),
.B1(n_1123),
.B2(n_1063),
.Y(n_2240)
);

BUFx8_ASAP7_75t_L g2241 ( 
.A(n_2016),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1933),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1981),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2017),
.B(n_2018),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2089),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2019),
.B(n_1072),
.Y(n_2246)
);

BUFx3_ASAP7_75t_L g2247 ( 
.A(n_2021),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_1923),
.A2(n_1991),
.B1(n_1926),
.B2(n_1930),
.Y(n_2248)
);

BUFx2_ASAP7_75t_L g2249 ( 
.A(n_1961),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_1927),
.B(n_1109),
.Y(n_2250)
);

OA21x2_ASAP7_75t_L g2251 ( 
.A1(n_1934),
.A2(n_1268),
.B(n_1267),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_1967),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_1953),
.B(n_1110),
.Y(n_2253)
);

OA21x2_ASAP7_75t_L g2254 ( 
.A1(n_1935),
.A2(n_1270),
.B(n_1267),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1936),
.B(n_1074),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2093),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_2047),
.B(n_1111),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1982),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1941),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2072),
.B(n_1120),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1943),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_1946),
.Y(n_2262)
);

NAND2xp33_ASAP7_75t_L g2263 ( 
.A(n_2002),
.B(n_1124),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2111),
.B(n_1076),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1948),
.B(n_1078),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1951),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2052),
.B(n_1126),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1954),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1984),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1985),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2083),
.B(n_1270),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_1957),
.A2(n_1327),
.B(n_1289),
.Y(n_2272)
);

BUFx12f_ASAP7_75t_L g2273 ( 
.A(n_2039),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2083),
.B(n_1289),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2033),
.A2(n_1239),
.B1(n_1245),
.B2(n_1198),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1942),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1925),
.B(n_1080),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_1931),
.A2(n_1125),
.B1(n_1129),
.B2(n_1124),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_1969),
.B(n_1134),
.Y(n_2279)
);

BUFx8_ASAP7_75t_SL g2280 ( 
.A(n_2043),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1990),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2097),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2049),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2102),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2056),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2104),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2105),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2107),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2108),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_1939),
.B(n_1082),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_1972),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2109),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2110),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2112),
.B(n_1083),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1955),
.B(n_1327),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_1997),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2062),
.B(n_1340),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2064),
.Y(n_2298)
);

OA21x2_ASAP7_75t_L g2299 ( 
.A1(n_2066),
.A2(n_1361),
.B(n_1340),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2081),
.A2(n_1129),
.B1(n_1135),
.B2(n_1125),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2085),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_L g2302 ( 
.A(n_2091),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2103),
.B(n_1220),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2095),
.Y(n_2304)
);

BUFx12f_ASAP7_75t_L g2305 ( 
.A(n_2100),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2071),
.B(n_1084),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2008),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1994),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1994),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2008),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2008),
.Y(n_2311)
);

OAI21x1_ASAP7_75t_L g2312 ( 
.A1(n_1918),
.A2(n_1389),
.B(n_1361),
.Y(n_2312)
);

INVx4_ASAP7_75t_L g2313 ( 
.A(n_2035),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2067),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2008),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_2067),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1952),
.B(n_1088),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1994),
.Y(n_2318)
);

OAI21x1_ASAP7_75t_L g2319 ( 
.A1(n_1918),
.A2(n_1409),
.B(n_1389),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1994),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_1938),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2008),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_1976),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_1976),
.Y(n_2324)
);

BUFx8_ASAP7_75t_L g2325 ( 
.A(n_1964),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2067),
.Y(n_2326)
);

CKINVDCx6p67_ASAP7_75t_R g2327 ( 
.A(n_1919),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2067),
.Y(n_2328)
);

HB1xp67_ASAP7_75t_L g2329 ( 
.A(n_1959),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_1952),
.B(n_1409),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2113),
.B(n_1136),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_1976),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2008),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_1959),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_1959),
.A2(n_1092),
.B1(n_1095),
.B2(n_1090),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1994),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2067),
.Y(n_2337)
);

OA21x2_ASAP7_75t_L g2338 ( 
.A1(n_1975),
.A2(n_1433),
.B(n_1427),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_2113),
.B(n_1137),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1994),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2113),
.B(n_1139),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_1944),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1994),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2113),
.B(n_1140),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2008),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_1976),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2008),
.Y(n_2347)
);

BUFx8_ASAP7_75t_L g2348 ( 
.A(n_1964),
.Y(n_2348)
);

INVxp33_ASAP7_75t_SL g2349 ( 
.A(n_1938),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2113),
.B(n_1141),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1994),
.Y(n_2351)
);

BUFx8_ASAP7_75t_SL g2352 ( 
.A(n_1938),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1994),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_1952),
.B(n_1427),
.Y(n_2354)
);

BUFx12f_ASAP7_75t_L g2355 ( 
.A(n_1938),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2008),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1952),
.B(n_1097),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_1959),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2113),
.B(n_1146),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2008),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2008),
.Y(n_2361)
);

INVx6_ASAP7_75t_L g2362 ( 
.A(n_2113),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_1976),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_1976),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1952),
.B(n_1433),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1994),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2071),
.B(n_1098),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2067),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_1952),
.B(n_1452),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1952),
.B(n_1099),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1994),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2008),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_2067),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_1959),
.A2(n_1105),
.B1(n_1107),
.B2(n_1104),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_2067),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1952),
.B(n_1452),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2008),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_1976),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2067),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2008),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1994),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1952),
.B(n_1113),
.Y(n_2382)
);

INVx5_ASAP7_75t_L g2383 ( 
.A(n_2067),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_2067),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1952),
.B(n_1115),
.Y(n_2385)
);

INVx4_ASAP7_75t_L g2386 ( 
.A(n_2035),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2101),
.B(n_1232),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2113),
.B(n_1150),
.Y(n_2388)
);

OAI21x1_ASAP7_75t_L g2389 ( 
.A1(n_1918),
.A2(n_1490),
.B(n_1470),
.Y(n_2389)
);

OA21x2_ASAP7_75t_L g2390 ( 
.A1(n_1975),
.A2(n_1490),
.B(n_1470),
.Y(n_2390)
);

AOI22x1_ASAP7_75t_SL g2391 ( 
.A1(n_2027),
.A2(n_1254),
.B1(n_1263),
.B2(n_1245),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2008),
.Y(n_2392)
);

NOR2x1_ASAP7_75t_L g2393 ( 
.A(n_2022),
.B(n_1157),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_1938),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2008),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2008),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_1956),
.A2(n_1142),
.B1(n_1143),
.B2(n_1135),
.Y(n_2397)
);

AND2x2_ASAP7_75t_SL g2398 ( 
.A(n_1945),
.B(n_1531),
.Y(n_2398)
);

OAI22x1_ASAP7_75t_R g2399 ( 
.A1(n_2027),
.A2(n_1263),
.B1(n_1272),
.B2(n_1254),
.Y(n_2399)
);

OA21x2_ASAP7_75t_L g2400 ( 
.A1(n_1975),
.A2(n_1534),
.B(n_1531),
.Y(n_2400)
);

OAI22x1_ASAP7_75t_L g2401 ( 
.A1(n_1956),
.A2(n_1142),
.B1(n_1145),
.B2(n_1143),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2008),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2101),
.B(n_1232),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_1976),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2067),
.Y(n_2405)
);

INVx3_ASAP7_75t_L g2406 ( 
.A(n_1976),
.Y(n_2406)
);

CKINVDCx8_ASAP7_75t_R g2407 ( 
.A(n_2099),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1959),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1994),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2008),
.Y(n_2410)
);

BUFx2_ASAP7_75t_L g2411 ( 
.A(n_1944),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_1956),
.A2(n_1148),
.B1(n_1149),
.B2(n_1145),
.Y(n_2412)
);

BUFx8_ASAP7_75t_L g2413 ( 
.A(n_1964),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2008),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_1938),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2113),
.B(n_1159),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_SL g2417 ( 
.A(n_1956),
.B(n_1272),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1994),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2008),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2008),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_1976),
.Y(n_2421)
);

INVx6_ASAP7_75t_L g2422 ( 
.A(n_2113),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2008),
.Y(n_2423)
);

INVx5_ASAP7_75t_L g2424 ( 
.A(n_2067),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2008),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2067),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_1952),
.B(n_1534),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2008),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1952),
.B(n_1119),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_2113),
.B(n_1163),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2008),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1994),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1994),
.Y(n_2433)
);

NAND2xp33_ASAP7_75t_L g2434 ( 
.A(n_2035),
.B(n_1148),
.Y(n_2434)
);

AND2x6_ASAP7_75t_L g2435 ( 
.A(n_1920),
.B(n_1537),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2067),
.Y(n_2436)
);

INVxp33_ASAP7_75t_SL g2437 ( 
.A(n_1938),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2067),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2008),
.Y(n_2439)
);

NOR2x1_ASAP7_75t_L g2440 ( 
.A(n_2022),
.B(n_1175),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2008),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_1952),
.B(n_1121),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1952),
.B(n_1171),
.Y(n_2443)
);

INVx6_ASAP7_75t_L g2444 ( 
.A(n_2113),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2113),
.B(n_1178),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1994),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2067),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2008),
.Y(n_2448)
);

OA21x2_ASAP7_75t_L g2449 ( 
.A1(n_1975),
.A2(n_1560),
.B(n_1537),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2067),
.Y(n_2450)
);

OAI21x1_ASAP7_75t_L g2451 ( 
.A1(n_1918),
.A2(n_1572),
.B(n_1560),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2008),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1994),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_SL g2454 ( 
.A(n_1956),
.B(n_1279),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1994),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2114),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_2140),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2135),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_2205),
.Y(n_2459)
);

AND2x2_ASAP7_75t_R g2460 ( 
.A(n_2399),
.B(n_2166),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2280),
.Y(n_2461)
);

INVx2_ASAP7_75t_SL g2462 ( 
.A(n_2204),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_R g2463 ( 
.A(n_2136),
.B(n_1172),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2352),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2321),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2394),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2114),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2415),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2273),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2224),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2239),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2276),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2349),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2226),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2437),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_2407),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2228),
.Y(n_2477)
);

CKINVDCx20_ASAP7_75t_R g2478 ( 
.A(n_2117),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2122),
.Y(n_2479)
);

BUFx6f_ASAP7_75t_L g2480 ( 
.A(n_2122),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2232),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2138),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2245),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2256),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2355),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_2305),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2217),
.B(n_1173),
.Y(n_2487)
);

BUFx10_ASAP7_75t_L g2488 ( 
.A(n_2264),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2284),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2327),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2135),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_2324),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2119),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2177),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2286),
.Y(n_2495)
);

CKINVDCx20_ASAP7_75t_R g2496 ( 
.A(n_2249),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2289),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2314),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2252),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2342),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2186),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_2411),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2313),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2386),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2182),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2302),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2293),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2302),
.Y(n_2508)
);

INVxp67_ASAP7_75t_L g2509 ( 
.A(n_2417),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_R g2510 ( 
.A(n_2195),
.B(n_1180),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2144),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_2346),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2283),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2285),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_2325),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2145),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2348),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_R g2518 ( 
.A(n_2434),
.B(n_1181),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2314),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_R g2520 ( 
.A(n_2200),
.B(n_1187),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2413),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2296),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2162),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2296),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2129),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_R g2526 ( 
.A(n_2304),
.B(n_1188),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2181),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2329),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2334),
.Y(n_2529)
);

HB1xp67_ASAP7_75t_L g2530 ( 
.A(n_2323),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2358),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2298),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2188),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2184),
.Y(n_2534)
);

INVxp67_ASAP7_75t_L g2535 ( 
.A(n_2454),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2123),
.B(n_2238),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_2291),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2306),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2247),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2262),
.B(n_1572),
.Y(n_2540)
);

BUFx10_ASAP7_75t_L g2541 ( 
.A(n_2367),
.Y(n_2541)
);

INVxp67_ASAP7_75t_SL g2542 ( 
.A(n_2363),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2378),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2137),
.Y(n_2544)
);

CKINVDCx20_ASAP7_75t_R g2545 ( 
.A(n_2301),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2421),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2137),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2277),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_2248),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2251),
.Y(n_2550)
);

INVxp33_ASAP7_75t_L g2551 ( 
.A(n_2275),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2290),
.Y(n_2552)
);

INVxp67_ASAP7_75t_L g2553 ( 
.A(n_2178),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2362),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2364),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2184),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2422),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_R g2558 ( 
.A(n_2172),
.B(n_1189),
.Y(n_2558)
);

CKINVDCx20_ASAP7_75t_R g2559 ( 
.A(n_2303),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_2444),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2128),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2404),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2406),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2254),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2194),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2131),
.B(n_1191),
.Y(n_2566)
);

CKINVDCx16_ASAP7_75t_R g2567 ( 
.A(n_2231),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2222),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2159),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2227),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2308),
.B(n_1587),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2237),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_R g2573 ( 
.A(n_2172),
.B(n_1193),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2398),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2242),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2194),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2335),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_R g2578 ( 
.A(n_2206),
.B(n_1195),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2374),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2259),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2261),
.Y(n_2581)
);

CKINVDCx20_ASAP7_75t_R g2582 ( 
.A(n_2149),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2408),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2266),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2309),
.B(n_1587),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2268),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2230),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2316),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2295),
.B(n_1232),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2230),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2316),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2126),
.Y(n_2592)
);

HB1xp67_ASAP7_75t_L g2593 ( 
.A(n_2126),
.Y(n_2593)
);

BUFx10_ASAP7_75t_L g2594 ( 
.A(n_2155),
.Y(n_2594)
);

AND3x2_ASAP7_75t_L g2595 ( 
.A(n_2183),
.B(n_1636),
.C(n_1615),
.Y(n_2595)
);

NAND2xp33_ASAP7_75t_R g2596 ( 
.A(n_2299),
.B(n_1149),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2332),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_R g2598 ( 
.A(n_2206),
.B(n_1196),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2234),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2295),
.B(n_1236),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_2332),
.Y(n_2601)
);

CKINVDCx20_ASAP7_75t_R g2602 ( 
.A(n_2210),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_2229),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2318),
.B(n_1615),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2391),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_2300),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2208),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2234),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2223),
.Y(n_2609)
);

INVx2_ASAP7_75t_SL g2610 ( 
.A(n_2215),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2115),
.B(n_1236),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2208),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2220),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2235),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2115),
.B(n_1236),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2320),
.B(n_1202),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2317),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2235),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2357),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2370),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2382),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2243),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_R g2623 ( 
.A(n_2336),
.B(n_1203),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2385),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2429),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_2442),
.Y(n_2626)
);

OR2x6_ASAP7_75t_L g2627 ( 
.A(n_2297),
.B(n_2173),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2243),
.Y(n_2628)
);

BUFx6f_ASAP7_75t_L g2629 ( 
.A(n_2326),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2258),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2220),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2297),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_2326),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_R g2634 ( 
.A(n_2340),
.B(n_1205),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2443),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2258),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2271),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2270),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2270),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2175),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2343),
.Y(n_2641)
);

BUFx10_ASAP7_75t_L g2642 ( 
.A(n_2331),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2351),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_2278),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_2161),
.Y(n_2645)
);

CKINVDCx20_ASAP7_75t_R g2646 ( 
.A(n_2199),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2353),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2240),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_2366),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_2387),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2271),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2371),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2381),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2409),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2418),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2330),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_2432),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2263),
.A2(n_2219),
.B1(n_2267),
.B2(n_2225),
.Y(n_2658)
);

NAND2xp33_ASAP7_75t_SL g2659 ( 
.A(n_2170),
.B(n_1279),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2328),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_R g2661 ( 
.A(n_2433),
.B(n_1206),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2446),
.Y(n_2662)
);

CKINVDCx20_ASAP7_75t_R g2663 ( 
.A(n_2403),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2328),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2453),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2339),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2455),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2241),
.Y(n_2668)
);

HB1xp67_ASAP7_75t_L g2669 ( 
.A(n_2274),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_R g2670 ( 
.A(n_2167),
.B(n_1207),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_2274),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2330),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2170),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_R g2674 ( 
.A(n_2180),
.B(n_1209),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2236),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2282),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2246),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2337),
.Y(n_2678)
);

CKINVDCx20_ASAP7_75t_R g2679 ( 
.A(n_2255),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2397),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2412),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_2203),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2265),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_R g2684 ( 
.A(n_2133),
.B(n_1210),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2294),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2341),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2257),
.B(n_1287),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2287),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2344),
.Y(n_2689)
);

CKINVDCx20_ASAP7_75t_R g2690 ( 
.A(n_2125),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2260),
.B(n_1287),
.Y(n_2691)
);

NAND2xp33_ASAP7_75t_R g2692 ( 
.A(n_2350),
.B(n_1151),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_R g2693 ( 
.A(n_2354),
.B(n_1211),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2359),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_R g2695 ( 
.A(n_2354),
.B(n_1213),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2288),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2388),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2416),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_R g2699 ( 
.A(n_2365),
.B(n_1214),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2430),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2292),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2445),
.B(n_1287),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2116),
.Y(n_2703)
);

NAND2xp33_ASAP7_75t_R g2704 ( 
.A(n_2250),
.B(n_1151),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2337),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2365),
.Y(n_2706)
);

NOR2xp67_ASAP7_75t_L g2707 ( 
.A(n_2202),
.B(n_1215),
.Y(n_2707)
);

NOR2xp67_ASAP7_75t_L g2708 ( 
.A(n_2202),
.B(n_1216),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2369),
.B(n_1636),
.Y(n_2709)
);

CKINVDCx20_ASAP7_75t_R g2710 ( 
.A(n_2369),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2376),
.Y(n_2711)
);

BUFx10_ASAP7_75t_L g2712 ( 
.A(n_2279),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2376),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2368),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2368),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2373),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_2427),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2281),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2373),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2427),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2141),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2401),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2401),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2375),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2253),
.Y(n_2725)
);

CKINVDCx16_ASAP7_75t_R g2726 ( 
.A(n_2160),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2375),
.Y(n_2727)
);

CKINVDCx16_ASAP7_75t_R g2728 ( 
.A(n_2160),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2156),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2147),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2379),
.Y(n_2731)
);

CKINVDCx16_ASAP7_75t_R g2732 ( 
.A(n_2193),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2151),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2193),
.Y(n_2734)
);

NAND2xp33_ASAP7_75t_R g2735 ( 
.A(n_2198),
.B(n_1152),
.Y(n_2735)
);

CKINVDCx5p33_ASAP7_75t_R g2736 ( 
.A(n_2156),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2169),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2169),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2233),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2244),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2218),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2198),
.Y(n_2742)
);

CKINVDCx20_ASAP7_75t_R g2743 ( 
.A(n_2120),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2269),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2379),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2384),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2384),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2405),
.Y(n_2748)
);

CKINVDCx20_ASAP7_75t_R g2749 ( 
.A(n_2192),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2405),
.Y(n_2750)
);

INVxp67_ASAP7_75t_SL g2751 ( 
.A(n_2426),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2426),
.Y(n_2752)
);

CKINVDCx20_ASAP7_75t_R g2753 ( 
.A(n_2338),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2153),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2436),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2154),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2130),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_R g2758 ( 
.A(n_2176),
.B(n_1217),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2157),
.Y(n_2759)
);

INVxp33_ASAP7_75t_L g2760 ( 
.A(n_2393),
.Y(n_2760)
);

CKINVDCx20_ASAP7_75t_R g2761 ( 
.A(n_2390),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2729),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2470),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2568),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2570),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2474),
.Y(n_2766)
);

AOI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_2743),
.A2(n_2435),
.B1(n_2139),
.B2(n_2272),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2477),
.Y(n_2768)
);

OR2x6_ASAP7_75t_L g2769 ( 
.A(n_2610),
.B(n_1317),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2481),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2572),
.Y(n_2771)
);

AND3x1_ASAP7_75t_L g2772 ( 
.A(n_2658),
.B(n_1183),
.C(n_1182),
.Y(n_2772)
);

AND2x6_ASAP7_75t_L g2773 ( 
.A(n_2550),
.B(n_2564),
.Y(n_2773)
);

OR2x6_ASAP7_75t_L g2774 ( 
.A(n_2462),
.B(n_1839),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2553),
.B(n_1114),
.Y(n_2775)
);

NAND3x1_ASAP7_75t_L g2776 ( 
.A(n_2460),
.B(n_1186),
.C(n_1184),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2683),
.B(n_2139),
.Y(n_2777)
);

BUFx10_ASAP7_75t_L g2778 ( 
.A(n_2464),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2483),
.Y(n_2779)
);

OR2x6_ASAP7_75t_L g2780 ( 
.A(n_2492),
.B(n_2440),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2484),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2589),
.B(n_2158),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2617),
.B(n_2139),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2575),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_2457),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2512),
.B(n_2171),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2619),
.B(n_2435),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2489),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2495),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2682),
.B(n_2620),
.Y(n_2790)
);

AO22x2_ASAP7_75t_L g2791 ( 
.A1(n_2509),
.A2(n_1106),
.B1(n_1176),
.B2(n_1122),
.Y(n_2791)
);

BUFx3_ASAP7_75t_L g2792 ( 
.A(n_2736),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2497),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_SL g2794 ( 
.A(n_2621),
.B(n_2436),
.Y(n_2794)
);

AND2x4_ASAP7_75t_L g2795 ( 
.A(n_2656),
.B(n_2164),
.Y(n_2795)
);

BUFx6f_ASAP7_75t_L g2796 ( 
.A(n_2456),
.Y(n_2796)
);

HB1xp67_ASAP7_75t_L g2797 ( 
.A(n_2632),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2624),
.B(n_2435),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2580),
.Y(n_2799)
);

BUFx3_ASAP7_75t_L g2800 ( 
.A(n_2737),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2456),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2587),
.B(n_2185),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2507),
.Y(n_2803)
);

AND2x6_ASAP7_75t_L g2804 ( 
.A(n_2611),
.B(n_1670),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2590),
.B(n_2187),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2721),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2625),
.B(n_2626),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2726),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2600),
.B(n_2728),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2738),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2732),
.B(n_1299),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2730),
.Y(n_2812)
);

AND2x6_ASAP7_75t_L g2813 ( 
.A(n_2615),
.B(n_1670),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2733),
.Y(n_2814)
);

OR2x6_ASAP7_75t_L g2815 ( 
.A(n_2627),
.B(n_1677),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2754),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2581),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2459),
.Y(n_2818)
);

INVx4_ASAP7_75t_L g2819 ( 
.A(n_2554),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2635),
.B(n_2438),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2584),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2536),
.B(n_2400),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2756),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2706),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2734),
.B(n_1299),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2759),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2487),
.B(n_2449),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2685),
.B(n_2739),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2506),
.Y(n_2829)
);

INVx2_ASAP7_75t_SL g2830 ( 
.A(n_2594),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2586),
.Y(n_2831)
);

INVx2_ASAP7_75t_SL g2832 ( 
.A(n_2594),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2599),
.B(n_2191),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2609),
.B(n_2538),
.Y(n_2834)
);

BUFx10_ASAP7_75t_L g2835 ( 
.A(n_2461),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2676),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2675),
.B(n_2118),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2742),
.B(n_1299),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2688),
.Y(n_2839)
);

AND2x6_ASAP7_75t_L g2840 ( 
.A(n_2511),
.B(n_1677),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2548),
.B(n_1212),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2696),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2701),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2718),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2552),
.B(n_1281),
.Y(n_2845)
);

INVx4_ASAP7_75t_L g2846 ( 
.A(n_2557),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2465),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2561),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2740),
.B(n_1304),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2637),
.Y(n_2850)
);

BUFx6f_ASAP7_75t_L g2851 ( 
.A(n_2456),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2651),
.Y(n_2852)
);

BUFx4f_ASAP7_75t_L g2853 ( 
.A(n_2627),
.Y(n_2853)
);

AND2x6_ASAP7_75t_L g2854 ( 
.A(n_2516),
.B(n_1692),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2669),
.Y(n_2855)
);

INVx3_ASAP7_75t_L g2856 ( 
.A(n_2467),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2677),
.B(n_1345),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2608),
.B(n_2214),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2757),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2671),
.Y(n_2860)
);

AND2x6_ASAP7_75t_L g2861 ( 
.A(n_2523),
.B(n_1692),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2672),
.B(n_2121),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2641),
.Y(n_2863)
);

NAND2x1p5_ASAP7_75t_L g2864 ( 
.A(n_2534),
.B(n_2213),
.Y(n_2864)
);

AND2x6_ASAP7_75t_L g2865 ( 
.A(n_2533),
.B(n_1781),
.Y(n_2865)
);

OR2x6_ASAP7_75t_L g2866 ( 
.A(n_2627),
.B(n_1781),
.Y(n_2866)
);

INVx4_ASAP7_75t_L g2867 ( 
.A(n_2560),
.Y(n_2867)
);

INVx4_ASAP7_75t_L g2868 ( 
.A(n_2745),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2643),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2647),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2749),
.A2(n_2221),
.B1(n_2134),
.B2(n_2143),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2654),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2665),
.Y(n_2873)
);

NAND2xp33_ASAP7_75t_R g2874 ( 
.A(n_2569),
.B(n_1152),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2534),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2713),
.B(n_1363),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2710),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2614),
.B(n_2132),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2571),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2556),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2585),
.Y(n_2881)
);

INVx5_ASAP7_75t_L g2882 ( 
.A(n_2467),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_SL g2883 ( 
.A(n_2476),
.B(n_1288),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2720),
.B(n_2124),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2709),
.B(n_2127),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2556),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2712),
.Y(n_2887)
);

NAND2x1p5_ASAP7_75t_L g2888 ( 
.A(n_2666),
.B(n_2146),
.Y(n_2888)
);

OR2x6_ASAP7_75t_L g2889 ( 
.A(n_2697),
.B(n_1790),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2649),
.B(n_1358),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2652),
.B(n_2438),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2508),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2753),
.B(n_2307),
.Y(n_2893)
);

BUFx3_ASAP7_75t_L g2894 ( 
.A(n_2746),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2604),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2618),
.B(n_2310),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2622),
.Y(n_2897)
);

AND3x4_ASAP7_75t_L g2898 ( 
.A(n_2551),
.B(n_1298),
.C(n_1288),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2747),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2761),
.B(n_2311),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2458),
.Y(n_2901)
);

INVx3_ASAP7_75t_L g2902 ( 
.A(n_2467),
.Y(n_2902)
);

AND2x6_ASAP7_75t_L g2903 ( 
.A(n_2539),
.B(n_1790),
.Y(n_2903)
);

INVx4_ASAP7_75t_L g2904 ( 
.A(n_2748),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2491),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2628),
.Y(n_2906)
);

BUFx12f_ASAP7_75t_L g2907 ( 
.A(n_2522),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2479),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2630),
.Y(n_2909)
);

INVx1_ASAP7_75t_SL g2910 ( 
.A(n_2524),
.Y(n_2910)
);

INVx2_ASAP7_75t_SL g2911 ( 
.A(n_2712),
.Y(n_2911)
);

INVx6_ASAP7_75t_L g2912 ( 
.A(n_2479),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2636),
.Y(n_2913)
);

BUFx6f_ASAP7_75t_L g2914 ( 
.A(n_2479),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2638),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2544),
.Y(n_2916)
);

AND2x4_ASAP7_75t_L g2917 ( 
.A(n_2639),
.B(n_2315),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2711),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2664),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2653),
.B(n_1382),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2547),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2542),
.B(n_2322),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2750),
.Y(n_2923)
);

AND2x6_ASAP7_75t_L g2924 ( 
.A(n_2678),
.B(n_1819),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_L g2925 ( 
.A(n_2655),
.B(n_1432),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2657),
.B(n_2333),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_L g2927 ( 
.A(n_2662),
.B(n_1478),
.Y(n_2927)
);

BUFx10_ASAP7_75t_L g2928 ( 
.A(n_2473),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2565),
.Y(n_2929)
);

AND2x6_ASAP7_75t_L g2930 ( 
.A(n_2705),
.B(n_1819),
.Y(n_2930)
);

INVxp33_ASAP7_75t_L g2931 ( 
.A(n_2558),
.Y(n_2931)
);

INVx6_ASAP7_75t_L g2932 ( 
.A(n_2480),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2576),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2714),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2715),
.Y(n_2935)
);

OR2x2_ASAP7_75t_L g2936 ( 
.A(n_2535),
.B(n_1484),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2679),
.A2(n_2142),
.B1(n_2150),
.B2(n_2148),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2667),
.B(n_2345),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2480),
.Y(n_2939)
);

NAND2x1p5_ASAP7_75t_L g2940 ( 
.A(n_2660),
.B(n_2196),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2716),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2744),
.B(n_2592),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2724),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2607),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2593),
.B(n_2597),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2660),
.Y(n_2946)
);

AND2x2_ASAP7_75t_SL g2947 ( 
.A(n_2567),
.B(n_1826),
.Y(n_2947)
);

AND2x6_ASAP7_75t_L g2948 ( 
.A(n_2612),
.B(n_1826),
.Y(n_2948)
);

BUFx3_ASAP7_75t_L g2949 ( 
.A(n_2752),
.Y(n_2949)
);

INVx3_ASAP7_75t_L g2950 ( 
.A(n_2480),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2601),
.B(n_2648),
.Y(n_2951)
);

CKINVDCx16_ASAP7_75t_R g2952 ( 
.A(n_2496),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2573),
.B(n_2447),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2578),
.B(n_2447),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2731),
.Y(n_2955)
);

BUFx3_ASAP7_75t_L g2956 ( 
.A(n_2755),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2598),
.B(n_2450),
.Y(n_2957)
);

BUFx2_ASAP7_75t_L g2958 ( 
.A(n_2717),
.Y(n_2958)
);

INVx2_ASAP7_75t_SL g2959 ( 
.A(n_2693),
.Y(n_2959)
);

HB1xp67_ASAP7_75t_L g2960 ( 
.A(n_2513),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2613),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2566),
.B(n_2616),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2731),
.Y(n_2963)
);

BUFx4f_ASAP7_75t_L g2964 ( 
.A(n_2498),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2695),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2631),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2493),
.B(n_2347),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2699),
.B(n_2356),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2562),
.B(n_1363),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2498),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2563),
.B(n_1363),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_L g2972 ( 
.A(n_2703),
.B(n_1497),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2530),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2680),
.B(n_1503),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2488),
.B(n_2541),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2645),
.B(n_2450),
.Y(n_2976)
);

BUFx3_ASAP7_75t_L g2977 ( 
.A(n_2543),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2540),
.B(n_2360),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2681),
.B(n_1599),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2555),
.Y(n_2980)
);

BUFx6f_ASAP7_75t_L g2981 ( 
.A(n_2498),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2519),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2546),
.B(n_2361),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2488),
.B(n_1366),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2519),
.Y(n_2985)
);

INVxp33_ASAP7_75t_L g2986 ( 
.A(n_2526),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2670),
.B(n_2152),
.Y(n_2987)
);

BUFx10_ASAP7_75t_L g2988 ( 
.A(n_2475),
.Y(n_2988)
);

BUFx4_ASAP7_75t_L g2989 ( 
.A(n_2482),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2519),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2541),
.B(n_2674),
.Y(n_2991)
);

AND2x4_ASAP7_75t_L g2992 ( 
.A(n_2751),
.B(n_2372),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2588),
.Y(n_2993)
);

NAND2x1p5_ASAP7_75t_L g2994 ( 
.A(n_2588),
.B(n_2209),
.Y(n_2994)
);

OR2x6_ASAP7_75t_L g2995 ( 
.A(n_2702),
.B(n_1883),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2588),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2574),
.B(n_1609),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2659),
.A2(n_2319),
.B1(n_2389),
.B2(n_2312),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2591),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2577),
.B(n_1635),
.Y(n_3000)
);

OR2x6_ASAP7_75t_L g3001 ( 
.A(n_2687),
.B(n_1883),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2591),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2591),
.Y(n_3003)
);

NOR2xp33_ASAP7_75t_L g3004 ( 
.A(n_2579),
.B(n_1643),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2499),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2629),
.Y(n_3006)
);

INVx5_ASAP7_75t_L g3007 ( 
.A(n_2629),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2962),
.B(n_2501),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2879),
.B(n_2503),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2881),
.B(n_2504),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2807),
.B(n_2606),
.Y(n_3011)
);

NOR2x1p5_ASAP7_75t_L g3012 ( 
.A(n_2810),
.B(n_2515),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2828),
.B(n_2505),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2895),
.B(n_2684),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2763),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_SL g3016 ( 
.A(n_2945),
.B(n_2510),
.Y(n_3016)
);

OR2x6_ASAP7_75t_L g3017 ( 
.A(n_2907),
.B(n_2691),
.Y(n_3017)
);

OAI22xp5_ASAP7_75t_SL g3018 ( 
.A1(n_2898),
.A2(n_2602),
.B1(n_2582),
.B2(n_2549),
.Y(n_3018)
);

OAI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2972),
.A2(n_2583),
.B1(n_2644),
.B2(n_2673),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2974),
.A2(n_2690),
.B1(n_2518),
.B2(n_2722),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_SL g3021 ( 
.A(n_2790),
.B(n_2809),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2829),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2766),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2768),
.Y(n_3024)
);

INVx4_ASAP7_75t_L g3025 ( 
.A(n_2892),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2849),
.B(n_2623),
.Y(n_3026)
);

INVxp67_ASAP7_75t_L g3027 ( 
.A(n_2936),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2770),
.Y(n_3028)
);

A2O1A1Ixp33_ASAP7_75t_L g3029 ( 
.A1(n_2857),
.A2(n_2760),
.B(n_2451),
.C(n_2723),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2779),
.Y(n_3030)
);

XOR2xp5_ASAP7_75t_L g3031 ( 
.A(n_2785),
.B(n_2471),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2775),
.B(n_2634),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2781),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2782),
.B(n_2661),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2979),
.B(n_2514),
.Y(n_3035)
);

INVxp33_ASAP7_75t_L g3036 ( 
.A(n_3000),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2863),
.B(n_2725),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2959),
.B(n_2525),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2762),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2870),
.B(n_2741),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2872),
.B(n_2532),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2869),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2841),
.B(n_2466),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2845),
.B(n_2595),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_3004),
.B(n_2468),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2873),
.Y(n_3046)
);

INVx2_ASAP7_75t_SL g3047 ( 
.A(n_2786),
.Y(n_3047)
);

INVxp67_ASAP7_75t_L g3048 ( 
.A(n_2890),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2796),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2920),
.B(n_2463),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2925),
.B(n_2686),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2788),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2965),
.B(n_2527),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2927),
.B(n_2689),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2789),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2997),
.B(n_2528),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2834),
.B(n_2472),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2885),
.B(n_2694),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2822),
.A2(n_2700),
.B(n_2698),
.Y(n_3059)
);

A2O1A1Ixp33_ASAP7_75t_L g3060 ( 
.A1(n_2783),
.A2(n_2646),
.B(n_2663),
.C(n_2650),
.Y(n_3060)
);

NOR3x1_ASAP7_75t_L g3061 ( 
.A(n_2877),
.B(n_1192),
.C(n_1190),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2808),
.Y(n_3062)
);

NOR2x1_ASAP7_75t_L g3063 ( 
.A(n_2792),
.B(n_2478),
.Y(n_3063)
);

INVx2_ASAP7_75t_SL g3064 ( 
.A(n_2912),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2931),
.B(n_2529),
.Y(n_3065)
);

INVxp33_ASAP7_75t_L g3066 ( 
.A(n_2960),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2951),
.B(n_2531),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2793),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2803),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2806),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2812),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2837),
.B(n_2707),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2825),
.B(n_2520),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2814),
.Y(n_3074)
);

AOI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2804),
.A2(n_2813),
.B1(n_2798),
.B2(n_2787),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2986),
.B(n_2545),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2816),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2823),
.B(n_2826),
.Y(n_3078)
);

AND2x4_ASAP7_75t_SL g3079 ( 
.A(n_2819),
.B(n_2500),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2827),
.A2(n_2708),
.B(n_2424),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2838),
.B(n_2642),
.Y(n_3081)
);

AOI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2804),
.A2(n_2596),
.B1(n_2640),
.B2(n_2559),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2824),
.B(n_2537),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2910),
.B(n_2502),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2797),
.B(n_2490),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2777),
.B(n_2642),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2862),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2773),
.B(n_2629),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2773),
.B(n_2633),
.Y(n_3089)
);

INVx2_ASAP7_75t_SL g3090 ( 
.A(n_2932),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_2800),
.Y(n_3091)
);

INVx2_ASAP7_75t_SL g3092 ( 
.A(n_2889),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2843),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2848),
.Y(n_3094)
);

AND2x6_ASAP7_75t_SL g3095 ( 
.A(n_2975),
.B(n_1199),
.Y(n_3095)
);

INVx8_ASAP7_75t_L g3096 ( 
.A(n_2882),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2773),
.B(n_2633),
.Y(n_3097)
);

INVx4_ASAP7_75t_L g3098 ( 
.A(n_2818),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2764),
.Y(n_3099)
);

AOI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_2804),
.A2(n_2704),
.B1(n_2735),
.B2(n_2692),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2795),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2942),
.B(n_2517),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2813),
.B(n_2633),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2813),
.B(n_2719),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2978),
.B(n_2719),
.Y(n_3105)
);

AOI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_2893),
.A2(n_1322),
.B1(n_1357),
.B2(n_1298),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2900),
.B(n_2719),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2765),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2926),
.B(n_2727),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2938),
.B(n_2968),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2991),
.B(n_2947),
.Y(n_3111)
);

INVx3_ASAP7_75t_L g3112 ( 
.A(n_2796),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2922),
.B(n_2727),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2853),
.B(n_2494),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_SL g3115 ( 
.A(n_2894),
.Y(n_3115)
);

BUFx3_ASAP7_75t_L g3116 ( 
.A(n_2899),
.Y(n_3116)
);

INVxp67_ASAP7_75t_L g3117 ( 
.A(n_2876),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_L g3118 ( 
.A(n_2883),
.B(n_2521),
.Y(n_3118)
);

OR2x2_ASAP7_75t_L g3119 ( 
.A(n_3005),
.B(n_2486),
.Y(n_3119)
);

AND2x6_ASAP7_75t_SL g3120 ( 
.A(n_2984),
.B(n_1204),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2967),
.B(n_2727),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2871),
.B(n_2758),
.Y(n_3122)
);

AOI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_2772),
.A2(n_2165),
.B1(n_2168),
.B2(n_2163),
.Y(n_3123)
);

INVx2_ASAP7_75t_SL g3124 ( 
.A(n_2983),
.Y(n_3124)
);

NAND2x1_ASAP7_75t_L g3125 ( 
.A(n_2801),
.B(n_2377),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_SL g3126 ( 
.A(n_2847),
.B(n_2485),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2884),
.B(n_2380),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2771),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2850),
.B(n_2469),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2969),
.B(n_2174),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2767),
.B(n_2392),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2784),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2799),
.Y(n_3133)
);

AND3x1_ASAP7_75t_L g3134 ( 
.A(n_2811),
.B(n_1221),
.C(n_1208),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_2852),
.A2(n_2860),
.B1(n_2855),
.B2(n_2840),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2971),
.B(n_2868),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2817),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_2958),
.B(n_1658),
.Y(n_3138)
);

OR2x6_ASAP7_75t_L g3139 ( 
.A(n_2949),
.B(n_1897),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_SL g3140 ( 
.A(n_2904),
.B(n_2190),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2821),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2831),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2836),
.B(n_2395),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2864),
.A2(n_2424),
.B(n_2383),
.Y(n_3144)
);

OAI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2888),
.A2(n_1357),
.B1(n_1411),
.B2(n_1322),
.Y(n_3145)
);

AND2x4_ASAP7_75t_L g3146 ( 
.A(n_2956),
.B(n_2846),
.Y(n_3146)
);

BUFx6f_ASAP7_75t_L g3147 ( 
.A(n_2801),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2998),
.A2(n_2980),
.B1(n_2973),
.B2(n_2815),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2839),
.B(n_2396),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2977),
.B(n_1366),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2842),
.B(n_2844),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2923),
.B(n_1366),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2992),
.B(n_2402),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2840),
.B(n_2410),
.Y(n_3154)
);

A2O1A1Ixp33_ASAP7_75t_L g3155 ( 
.A1(n_2897),
.A2(n_1686),
.B(n_1701),
.C(n_1663),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_SL g3156 ( 
.A(n_2859),
.B(n_2197),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2840),
.B(n_2414),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2866),
.B(n_1388),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2937),
.B(n_2201),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2896),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2917),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2940),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2878),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2906),
.Y(n_3164)
);

A2O1A1Ixp33_ASAP7_75t_L g3165 ( 
.A1(n_2909),
.A2(n_1827),
.B(n_1896),
.C(n_1709),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2854),
.B(n_2419),
.Y(n_3166)
);

INVxp67_ASAP7_75t_L g3167 ( 
.A(n_2918),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2780),
.B(n_1388),
.Y(n_3168)
);

BUFx8_ASAP7_75t_L g3169 ( 
.A(n_2887),
.Y(n_3169)
);

INVx1_ASAP7_75t_SL g3170 ( 
.A(n_2952),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2901),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2905),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2854),
.B(n_2420),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2830),
.B(n_1388),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_2832),
.B(n_1395),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_SL g3176 ( 
.A(n_2964),
.B(n_2882),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2854),
.B(n_2423),
.Y(n_3177)
);

NAND2x1p5_ASAP7_75t_L g3178 ( 
.A(n_2867),
.B(n_2425),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_SL g3179 ( 
.A(n_2928),
.B(n_2668),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2916),
.Y(n_3180)
);

INVxp67_ASAP7_75t_L g3181 ( 
.A(n_2874),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2861),
.B(n_2428),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2861),
.B(n_2431),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_3007),
.B(n_2207),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2913),
.Y(n_3185)
);

AND2x4_ASAP7_75t_L g3186 ( 
.A(n_2875),
.B(n_2439),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2861),
.B(n_2441),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2865),
.B(n_2448),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_SL g3189 ( 
.A(n_3007),
.B(n_2211),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2851),
.B(n_2212),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2794),
.B(n_1411),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2915),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2769),
.B(n_1395),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2865),
.B(n_2452),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2865),
.B(n_2216),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2820),
.B(n_1434),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2903),
.B(n_2179),
.Y(n_3197)
);

OAI221xp5_ASAP7_75t_L g3198 ( 
.A1(n_3001),
.A2(n_1916),
.B1(n_1237),
.B2(n_1240),
.C(n_1230),
.Y(n_3198)
);

OR2x6_ASAP7_75t_L g3199 ( 
.A(n_2911),
.B(n_1897),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2903),
.B(n_2189),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_SL g3201 ( 
.A(n_2778),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_2851),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2903),
.A2(n_1458),
.B1(n_1505),
.B2(n_1434),
.Y(n_3203)
);

AND2x2_ASAP7_75t_L g3204 ( 
.A(n_2988),
.B(n_1395),
.Y(n_3204)
);

NAND3xp33_ASAP7_75t_L g3205 ( 
.A(n_2891),
.B(n_2605),
.C(n_2603),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2921),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_2908),
.B(n_2914),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2908),
.B(n_1458),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3110),
.A2(n_2987),
.B(n_2994),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3015),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3131),
.A2(n_2976),
.B(n_2954),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3072),
.A2(n_2957),
.B(n_2953),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3008),
.B(n_2929),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_3087),
.B(n_2933),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_3062),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3032),
.B(n_3048),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3162),
.A2(n_2886),
.B(n_2880),
.Y(n_3217)
);

BUFx8_ASAP7_75t_L g3218 ( 
.A(n_3115),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3023),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3011),
.A2(n_2955),
.B1(n_2963),
.B2(n_2946),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_3091),
.B(n_2966),
.Y(n_3221)
);

INVx2_ASAP7_75t_SL g3222 ( 
.A(n_3096),
.Y(n_3222)
);

OAI22x1_ASAP7_75t_L g3223 ( 
.A1(n_3100),
.A2(n_2776),
.B1(n_1154),
.B2(n_1155),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3121),
.B(n_2802),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3036),
.B(n_2774),
.Y(n_3225)
);

CKINVDCx10_ASAP7_75t_R g3226 ( 
.A(n_3201),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_3105),
.A2(n_2961),
.B(n_2944),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3024),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3052),
.Y(n_3229)
);

OAI21xp33_ASAP7_75t_L g3230 ( 
.A1(n_3203),
.A2(n_2791),
.B(n_2995),
.Y(n_3230)
);

NOR2x1p5_ASAP7_75t_SL g3231 ( 
.A(n_3042),
.B(n_2970),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_3009),
.B(n_2914),
.Y(n_3232)
);

O2A1O1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_3111),
.A2(n_2934),
.B(n_2935),
.C(n_2919),
.Y(n_3233)
);

OAI21xp33_ASAP7_75t_L g3234 ( 
.A1(n_3045),
.A2(n_1514),
.B(n_1505),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3026),
.B(n_2996),
.Y(n_3235)
);

BUFx3_ASAP7_75t_L g3236 ( 
.A(n_3022),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3050),
.B(n_3043),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3034),
.A2(n_3003),
.B(n_2981),
.Y(n_3238)
);

NOR3xp33_ASAP7_75t_L g3239 ( 
.A(n_3067),
.B(n_2902),
.C(n_2856),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_3098),
.Y(n_3240)
);

INVx4_ASAP7_75t_L g3241 ( 
.A(n_3096),
.Y(n_3241)
);

BUFx6f_ASAP7_75t_L g3242 ( 
.A(n_3049),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_3069),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3127),
.A2(n_2981),
.B(n_2982),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3028),
.Y(n_3245)
);

NOR2xp67_ASAP7_75t_L g3246 ( 
.A(n_3025),
.B(n_2941),
.Y(n_3246)
);

OAI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_3029),
.A2(n_2943),
.B(n_2833),
.Y(n_3247)
);

NAND2xp33_ASAP7_75t_L g3248 ( 
.A(n_3014),
.B(n_2985),
.Y(n_3248)
);

O2A1O1Ixp33_ASAP7_75t_L g3249 ( 
.A1(n_3122),
.A2(n_2993),
.B(n_2999),
.C(n_2990),
.Y(n_3249)
);

OAI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_3075),
.A2(n_2858),
.B(n_2805),
.Y(n_3250)
);

OR2x2_ASAP7_75t_L g3251 ( 
.A(n_3035),
.B(n_3138),
.Y(n_3251)
);

O2A1O1Ixp33_ASAP7_75t_L g3252 ( 
.A1(n_3044),
.A2(n_3006),
.B(n_3002),
.C(n_2950),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3010),
.B(n_2939),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_3046),
.A2(n_2948),
.B1(n_2930),
.B2(n_2924),
.Y(n_3254)
);

BUFx4f_ASAP7_75t_L g3255 ( 
.A(n_3146),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3113),
.A2(n_2383),
.B(n_1241),
.Y(n_3256)
);

A2O1A1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_3191),
.A2(n_1242),
.B(n_1246),
.C(n_1224),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3058),
.B(n_2948),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3078),
.B(n_2948),
.Y(n_3259)
);

OR2x2_ASAP7_75t_L g3260 ( 
.A(n_3027),
.B(n_1153),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_3167),
.Y(n_3261)
);

INVx2_ASAP7_75t_SL g3262 ( 
.A(n_3039),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3094),
.Y(n_3263)
);

NOR2xp67_ASAP7_75t_L g3264 ( 
.A(n_3117),
.B(n_3057),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_3107),
.B(n_2924),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_3049),
.Y(n_3266)
);

OAI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3030),
.A2(n_2930),
.B(n_2924),
.Y(n_3267)
);

INVx2_ASAP7_75t_SL g3268 ( 
.A(n_3116),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3109),
.A2(n_1256),
.B(n_1252),
.Y(n_3269)
);

AO21x1_ASAP7_75t_L g3270 ( 
.A1(n_3148),
.A2(n_1274),
.B(n_1265),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3056),
.B(n_2835),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3033),
.A2(n_2930),
.B(n_1282),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3153),
.A2(n_1285),
.B(n_1275),
.Y(n_3273)
);

AOI21x1_ASAP7_75t_L g3274 ( 
.A1(n_3080),
.A2(n_1296),
.B(n_1290),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_3051),
.B(n_1514),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3055),
.B(n_1219),
.Y(n_3276)
);

A2O1A1Ixp33_ASAP7_75t_L g3277 ( 
.A1(n_3196),
.A2(n_1303),
.B(n_1307),
.C(n_1300),
.Y(n_3277)
);

NOR2x1_ASAP7_75t_L g3278 ( 
.A(n_3073),
.B(n_1529),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_SL g3279 ( 
.A(n_3054),
.B(n_1529),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3068),
.B(n_1222),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3093),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3151),
.A2(n_1309),
.B(n_1308),
.Y(n_3282)
);

CKINVDCx10_ASAP7_75t_R g3283 ( 
.A(n_3017),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_3019),
.B(n_1530),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3070),
.Y(n_3285)
);

AOI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3088),
.A2(n_1318),
.B(n_1314),
.Y(n_3286)
);

NOR3xp33_ASAP7_75t_L g3287 ( 
.A(n_3018),
.B(n_1227),
.C(n_1223),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3071),
.B(n_1228),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3089),
.A2(n_1325),
.B(n_1320),
.Y(n_3289)
);

CKINVDCx5p33_ASAP7_75t_R g3290 ( 
.A(n_3079),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3074),
.B(n_1229),
.Y(n_3291)
);

AO21x1_ASAP7_75t_L g3292 ( 
.A1(n_3159),
.A2(n_1335),
.B(n_1330),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_3097),
.A2(n_1342),
.B(n_1338),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3077),
.B(n_1231),
.Y(n_3294)
);

NAND2x1p5_ASAP7_75t_L g3295 ( 
.A(n_3147),
.B(n_2989),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_3147),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3059),
.A2(n_1359),
.B(n_1348),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_3086),
.A2(n_3041),
.B(n_3021),
.Y(n_3298)
);

AOI21x1_ASAP7_75t_L g3299 ( 
.A1(n_3154),
.A2(n_1371),
.B(n_1362),
.Y(n_3299)
);

AOI21x1_ASAP7_75t_L g3300 ( 
.A1(n_3157),
.A2(n_1381),
.B(n_1375),
.Y(n_3300)
);

NOR2xp33_ASAP7_75t_R g3301 ( 
.A(n_3126),
.B(n_3179),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3108),
.B(n_1233),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3103),
.A2(n_1385),
.B(n_1384),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3040),
.B(n_1530),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3099),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3164),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3132),
.Y(n_3307)
);

AO21x1_ASAP7_75t_L g3308 ( 
.A1(n_3016),
.A2(n_3195),
.B(n_3173),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3128),
.B(n_1235),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3141),
.B(n_1238),
.Y(n_3310)
);

NOR2x1p5_ASAP7_75t_L g3311 ( 
.A(n_3119),
.B(n_1153),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3020),
.A2(n_1597),
.B1(n_1616),
.B2(n_1563),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3104),
.A2(n_1393),
.B(n_1391),
.Y(n_3313)
);

A2O1A1Ixp33_ASAP7_75t_L g3314 ( 
.A1(n_3135),
.A2(n_1396),
.B(n_1401),
.C(n_1394),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3142),
.B(n_1243),
.Y(n_3315)
);

OAI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3185),
.A2(n_3192),
.B(n_3137),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3037),
.B(n_1563),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3133),
.B(n_1247),
.Y(n_3318)
);

NOR3xp33_ASAP7_75t_L g3319 ( 
.A(n_3065),
.B(n_1250),
.C(n_1249),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3082),
.A2(n_1616),
.B1(n_1713),
.B2(n_1597),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3171),
.Y(n_3321)
);

BUFx6f_ASAP7_75t_L g3322 ( 
.A(n_3121),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3081),
.B(n_1255),
.Y(n_3323)
);

CKINVDCx12_ASAP7_75t_R g3324 ( 
.A(n_3017),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3130),
.A2(n_1405),
.B(n_1404),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3143),
.Y(n_3326)
);

A2O1A1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_3172),
.A2(n_1421),
.B(n_1422),
.C(n_1412),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3181),
.B(n_1397),
.Y(n_3328)
);

AOI21xp33_ASAP7_75t_L g3329 ( 
.A1(n_3066),
.A2(n_1714),
.B(n_1713),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3145),
.B(n_3208),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3180),
.A2(n_1725),
.B1(n_1729),
.B2(n_1714),
.Y(n_3331)
);

INVx11_ASAP7_75t_L g3332 ( 
.A(n_3169),
.Y(n_3332)
);

O2A1O1Ixp33_ASAP7_75t_L g3333 ( 
.A1(n_3155),
.A2(n_1425),
.B(n_1428),
.C(n_1426),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3206),
.B(n_1258),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3186),
.B(n_1259),
.Y(n_3335)
);

O2A1O1Ixp33_ASAP7_75t_L g3336 ( 
.A1(n_3165),
.A2(n_1430),
.B(n_1437),
.C(n_1435),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3186),
.B(n_1260),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3106),
.B(n_1154),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_3084),
.B(n_1725),
.Y(n_3339)
);

AOI21xp33_ASAP7_75t_L g3340 ( 
.A1(n_3085),
.A2(n_3129),
.B(n_3124),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3197),
.A2(n_1461),
.B(n_1455),
.Y(n_3341)
);

NAND2x1p5_ASAP7_75t_L g3342 ( 
.A(n_3112),
.B(n_3047),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3200),
.A2(n_1469),
.B(n_1467),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3166),
.A2(n_1480),
.B(n_1473),
.Y(n_3344)
);

BUFx12f_ASAP7_75t_L g3345 ( 
.A(n_3012),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3177),
.A2(n_1485),
.B(n_1482),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3182),
.A2(n_1495),
.B(n_1487),
.Y(n_3347)
);

AO21x1_ASAP7_75t_L g3348 ( 
.A1(n_3183),
.A2(n_1516),
.B(n_1501),
.Y(n_3348)
);

INVxp67_ASAP7_75t_L g3349 ( 
.A(n_3150),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3060),
.A2(n_3101),
.B1(n_3136),
.B2(n_3160),
.Y(n_3350)
);

BUFx12f_ASAP7_75t_L g3351 ( 
.A(n_3095),
.Y(n_3351)
);

OR2x6_ASAP7_75t_L g3352 ( 
.A(n_3092),
.B(n_1915),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3187),
.A2(n_3194),
.B(n_3188),
.Y(n_3353)
);

INVx4_ASAP7_75t_L g3354 ( 
.A(n_3139),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3149),
.A2(n_1524),
.B(n_1517),
.Y(n_3355)
);

AO21x1_ASAP7_75t_L g3356 ( 
.A1(n_3190),
.A2(n_1528),
.B(n_1525),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3207),
.A2(n_1545),
.B(n_1543),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3156),
.Y(n_3358)
);

O2A1O1Ixp5_ASAP7_75t_L g3359 ( 
.A1(n_3125),
.A2(n_1915),
.B(n_1565),
.C(n_1567),
.Y(n_3359)
);

INVx4_ASAP7_75t_L g3360 ( 
.A(n_3255),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3237),
.B(n_3339),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3209),
.A2(n_3140),
.B(n_3013),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_3330),
.A2(n_3102),
.B(n_3118),
.C(n_3152),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3353),
.A2(n_3053),
.B(n_3038),
.Y(n_3364)
);

NAND3xp33_ASAP7_75t_SL g3365 ( 
.A(n_3275),
.B(n_3204),
.C(n_3198),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_R g3366 ( 
.A(n_3290),
.B(n_3170),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3216),
.B(n_3076),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_3284),
.B(n_3083),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3326),
.B(n_3174),
.Y(n_3369)
);

HB1xp67_ASAP7_75t_L g3370 ( 
.A(n_3215),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3264),
.A2(n_3134),
.B1(n_3161),
.B2(n_3163),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3281),
.Y(n_3372)
);

BUFx3_ASAP7_75t_L g3373 ( 
.A(n_3236),
.Y(n_3373)
);

BUFx3_ASAP7_75t_L g3374 ( 
.A(n_3296),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3212),
.A2(n_3176),
.B(n_3144),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3278),
.B(n_3139),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_3234),
.B(n_3031),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3240),
.B(n_3063),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_3261),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3210),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_3247),
.A2(n_3250),
.B(n_3298),
.Y(n_3381)
);

INVx8_ASAP7_75t_L g3382 ( 
.A(n_3242),
.Y(n_3382)
);

NAND3xp33_ASAP7_75t_L g3383 ( 
.A(n_3319),
.B(n_3175),
.C(n_3205),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_3251),
.B(n_3168),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3219),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3262),
.B(n_3064),
.Y(n_3386)
);

BUFx3_ASAP7_75t_L g3387 ( 
.A(n_3242),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3213),
.B(n_3158),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3228),
.Y(n_3389)
);

BUFx8_ASAP7_75t_L g3390 ( 
.A(n_3345),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_L g3391 ( 
.A(n_3279),
.B(n_3312),
.Y(n_3391)
);

NOR3xp33_ASAP7_75t_SL g3392 ( 
.A(n_3230),
.B(n_3114),
.C(n_1156),
.Y(n_3392)
);

BUFx3_ASAP7_75t_L g3393 ( 
.A(n_3242),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3235),
.B(n_3202),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3320),
.B(n_3193),
.Y(n_3395)
);

AOI21x1_ASAP7_75t_L g3396 ( 
.A1(n_3308),
.A2(n_3189),
.B(n_3184),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3328),
.B(n_3199),
.Y(n_3397)
);

INVx5_ASAP7_75t_L g3398 ( 
.A(n_3266),
.Y(n_3398)
);

A2O1A1Ixp33_ASAP7_75t_L g3399 ( 
.A1(n_3211),
.A2(n_3123),
.B(n_1571),
.C(n_1574),
.Y(n_3399)
);

OR2x2_ASAP7_75t_L g3400 ( 
.A(n_3260),
.B(n_3090),
.Y(n_3400)
);

OAI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3245),
.A2(n_3178),
.B1(n_3199),
.B2(n_1737),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_R g3402 ( 
.A(n_3268),
.B(n_3120),
.Y(n_3402)
);

OAI22x1_ASAP7_75t_L g3403 ( 
.A1(n_3317),
.A2(n_1156),
.B1(n_1158),
.B2(n_1155),
.Y(n_3403)
);

OAI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3316),
.A2(n_1576),
.B(n_1553),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3257),
.A2(n_1579),
.B(n_1580),
.C(n_1578),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3271),
.B(n_3061),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3285),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_3266),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3248),
.A2(n_1589),
.B(n_1583),
.Y(n_3409)
);

NOR2x1_ASAP7_75t_SL g3410 ( 
.A(n_3220),
.B(n_1600),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3266),
.Y(n_3411)
);

OR2x2_ASAP7_75t_L g3412 ( 
.A(n_3338),
.B(n_1158),
.Y(n_3412)
);

HB1xp67_ASAP7_75t_L g3413 ( 
.A(n_3322),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3258),
.A2(n_3253),
.B(n_3227),
.Y(n_3414)
);

AOI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_3304),
.A2(n_1737),
.B1(n_1758),
.B2(n_1729),
.Y(n_3415)
);

A2O1A1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_3333),
.A2(n_1607),
.B(n_1610),
.C(n_1603),
.Y(n_3416)
);

NOR3xp33_ASAP7_75t_L g3417 ( 
.A(n_3340),
.B(n_1637),
.C(n_1618),
.Y(n_3417)
);

CKINVDCx5p33_ASAP7_75t_R g3418 ( 
.A(n_3226),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3306),
.Y(n_3419)
);

O2A1O1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_3277),
.A2(n_1614),
.B(n_1623),
.C(n_1622),
.Y(n_3420)
);

O2A1O1Ixp33_ASAP7_75t_L g3421 ( 
.A1(n_3350),
.A2(n_1631),
.B(n_1639),
.C(n_1632),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_3232),
.A2(n_1650),
.B(n_1641),
.Y(n_3422)
);

AOI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3225),
.A2(n_1759),
.B1(n_1764),
.B2(n_1758),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3265),
.A2(n_1656),
.B(n_1651),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_3336),
.A2(n_1666),
.B(n_1672),
.C(n_1668),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3214),
.B(n_1673),
.Y(n_3426)
);

NOR2xp67_ASAP7_75t_SL g3427 ( 
.A(n_3241),
.B(n_1164),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_3224),
.B(n_1674),
.Y(n_3428)
);

OAI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_3229),
.A2(n_3243),
.B1(n_3349),
.B2(n_3259),
.Y(n_3429)
);

O2A1O1Ixp33_ASAP7_75t_L g3430 ( 
.A1(n_3329),
.A2(n_1676),
.B(n_1682),
.C(n_1681),
.Y(n_3430)
);

O2A1O1Ixp5_ASAP7_75t_L g3431 ( 
.A1(n_3270),
.A2(n_1685),
.B(n_1699),
.C(n_1696),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_3233),
.A2(n_1703),
.B(n_1704),
.C(n_1702),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3244),
.A2(n_1712),
.B(n_1705),
.Y(n_3433)
);

BUFx8_ASAP7_75t_SL g3434 ( 
.A(n_3351),
.Y(n_3434)
);

O2A1O1Ixp5_ASAP7_75t_L g3435 ( 
.A1(n_3274),
.A2(n_1716),
.B(n_1718),
.C(n_1717),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3323),
.B(n_1759),
.Y(n_3436)
);

CKINVDCx5p33_ASAP7_75t_R g3437 ( 
.A(n_3301),
.Y(n_3437)
);

OR2x2_ASAP7_75t_L g3438 ( 
.A(n_3335),
.B(n_1164),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3305),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3307),
.B(n_1719),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3224),
.B(n_3287),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3263),
.Y(n_3442)
);

HB1xp67_ASAP7_75t_L g3443 ( 
.A(n_3322),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3238),
.A2(n_1724),
.B(n_1720),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_3322),
.B(n_1764),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3252),
.A2(n_1734),
.B(n_1733),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_3221),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3331),
.B(n_1773),
.Y(n_3448)
);

OA22x2_ASAP7_75t_L g3449 ( 
.A1(n_3223),
.A2(n_3352),
.B1(n_3354),
.B2(n_3221),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3249),
.A2(n_1748),
.B(n_1738),
.Y(n_3450)
);

BUFx4f_ASAP7_75t_L g3451 ( 
.A(n_3295),
.Y(n_3451)
);

BUFx4f_ASAP7_75t_L g3452 ( 
.A(n_3222),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3342),
.Y(n_3453)
);

BUFx6f_ASAP7_75t_L g3454 ( 
.A(n_3352),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3321),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3276),
.B(n_1761),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3246),
.B(n_1773),
.Y(n_3457)
);

OAI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3217),
.A2(n_1767),
.B(n_1765),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_3239),
.B(n_1795),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3272),
.A2(n_1789),
.B(n_1778),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3280),
.B(n_1796),
.Y(n_3461)
);

CKINVDCx11_ASAP7_75t_R g3462 ( 
.A(n_3332),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3288),
.B(n_1795),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3291),
.B(n_1799),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3358),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_3318),
.A2(n_1809),
.B(n_1800),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_L g3467 ( 
.A1(n_3356),
.A2(n_1808),
.B1(n_1812),
.B2(n_1804),
.Y(n_3467)
);

BUFx8_ASAP7_75t_SL g3468 ( 
.A(n_3337),
.Y(n_3468)
);

O2A1O1Ixp33_ASAP7_75t_L g3469 ( 
.A1(n_3327),
.A2(n_1811),
.B(n_1817),
.C(n_1810),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_3294),
.B(n_1804),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3334),
.A2(n_1828),
.B(n_1821),
.Y(n_3471)
);

NOR3xp33_ASAP7_75t_L g3472 ( 
.A(n_3302),
.B(n_1867),
.C(n_1829),
.Y(n_3472)
);

NAND2x1p5_ASAP7_75t_L g3473 ( 
.A(n_3311),
.B(n_1836),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3267),
.A2(n_1861),
.B(n_1860),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3309),
.A2(n_1873),
.B(n_1866),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3299),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3310),
.B(n_1808),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3300),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3286),
.Y(n_3479)
);

BUFx6f_ASAP7_75t_L g3480 ( 
.A(n_3315),
.Y(n_3480)
);

A2O1A1Ixp33_ASAP7_75t_L g3481 ( 
.A1(n_3297),
.A2(n_1895),
.B(n_1898),
.C(n_1888),
.Y(n_3481)
);

NAND2xp33_ASAP7_75t_SL g3482 ( 
.A(n_3254),
.B(n_1812),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3269),
.B(n_1261),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3282),
.B(n_3273),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3314),
.B(n_1262),
.Y(n_3485)
);

INVx2_ASAP7_75t_SL g3486 ( 
.A(n_3283),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3256),
.A2(n_1822),
.B(n_1818),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3359),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3324),
.B(n_1818),
.Y(n_3489)
);

A2O1A1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3289),
.A2(n_1863),
.B(n_1874),
.C(n_1822),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3344),
.B(n_1264),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3292),
.B(n_1863),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3346),
.B(n_1269),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3303),
.A2(n_1886),
.B1(n_1890),
.B2(n_1874),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3231),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3348),
.B(n_1886),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3313),
.A2(n_1891),
.B1(n_1890),
.B2(n_1167),
.Y(n_3497)
);

INVx3_ASAP7_75t_L g3498 ( 
.A(n_3218),
.Y(n_3498)
);

BUFx6f_ASAP7_75t_L g3499 ( 
.A(n_3218),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_3370),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3381),
.A2(n_3347),
.B(n_3343),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3385),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3361),
.B(n_3341),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3389),
.Y(n_3504)
);

OAI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3363),
.A2(n_3293),
.B(n_3325),
.Y(n_3505)
);

AO31x2_ASAP7_75t_L g3506 ( 
.A1(n_3488),
.A2(n_3355),
.A3(n_3357),
.B(n_1584),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3367),
.B(n_1166),
.Y(n_3507)
);

AO31x2_ASAP7_75t_L g3508 ( 
.A1(n_3476),
.A2(n_2),
.A3(n_0),
.B(n_1),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3484),
.A2(n_1891),
.B(n_1273),
.Y(n_3509)
);

AOI221x1_ASAP7_75t_L g3510 ( 
.A1(n_3391),
.A2(n_1504),
.B1(n_1511),
.B2(n_1448),
.C(n_1397),
.Y(n_3510)
);

AOI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_3368),
.A2(n_1276),
.B1(n_1277),
.B2(n_1271),
.Y(n_3511)
);

OAI21x1_ASAP7_75t_L g3512 ( 
.A1(n_3414),
.A2(n_2),
.B(n_3),
.Y(n_3512)
);

OAI21x1_ASAP7_75t_L g3513 ( 
.A1(n_3375),
.A2(n_3),
.B(n_4),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3477),
.B(n_3436),
.Y(n_3514)
);

INVx3_ASAP7_75t_L g3515 ( 
.A(n_3373),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3360),
.B(n_1166),
.Y(n_3516)
);

OAI21x1_ASAP7_75t_L g3517 ( 
.A1(n_3362),
.A2(n_3),
.B(n_5),
.Y(n_3517)
);

OAI21x1_ASAP7_75t_L g3518 ( 
.A1(n_3364),
.A2(n_5),
.B(n_6),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3407),
.Y(n_3519)
);

AOI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3395),
.A2(n_1280),
.B1(n_1283),
.B2(n_1278),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3404),
.A2(n_3369),
.B(n_3388),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3480),
.B(n_1167),
.Y(n_3522)
);

AO31x2_ASAP7_75t_L g3523 ( 
.A1(n_3478),
.A2(n_8),
.A3(n_6),
.B(n_7),
.Y(n_3523)
);

OAI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3365),
.A2(n_1917),
.B(n_1291),
.Y(n_3524)
);

BUFx2_ASAP7_75t_L g3525 ( 
.A(n_3379),
.Y(n_3525)
);

AOI221x1_ASAP7_75t_L g3526 ( 
.A1(n_3482),
.A2(n_1504),
.B1(n_1511),
.B2(n_1448),
.C(n_1397),
.Y(n_3526)
);

OAI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3396),
.A2(n_3479),
.B(n_3495),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3419),
.Y(n_3528)
);

OAI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3433),
.A2(n_6),
.B(n_7),
.Y(n_3529)
);

OAI21xp5_ASAP7_75t_L g3530 ( 
.A1(n_3421),
.A2(n_1292),
.B(n_1286),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3480),
.B(n_1169),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3374),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3383),
.A2(n_1295),
.B(n_1293),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3492),
.B(n_1169),
.Y(n_3534)
);

NOR2xp67_ASAP7_75t_L g3535 ( 
.A(n_3437),
.B(n_7),
.Y(n_3535)
);

AO31x2_ASAP7_75t_L g3536 ( 
.A1(n_3410),
.A2(n_10),
.A3(n_8),
.B(n_9),
.Y(n_3536)
);

AO31x2_ASAP7_75t_L g3537 ( 
.A1(n_3399),
.A2(n_10),
.A3(n_8),
.B(n_9),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3401),
.B(n_3378),
.Y(n_3538)
);

OR2x2_ASAP7_75t_L g3539 ( 
.A(n_3445),
.B(n_1170),
.Y(n_3539)
);

OAI21x1_ASAP7_75t_L g3540 ( 
.A1(n_3444),
.A2(n_9),
.B(n_10),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3394),
.B(n_1170),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3429),
.A2(n_1310),
.B(n_1305),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3397),
.B(n_1448),
.Y(n_3543)
);

OAI21x1_ASAP7_75t_L g3544 ( 
.A1(n_3435),
.A2(n_11),
.B(n_12),
.Y(n_3544)
);

OAI21x1_ASAP7_75t_L g3545 ( 
.A1(n_3474),
.A2(n_11),
.B(n_12),
.Y(n_3545)
);

AOI21x1_ASAP7_75t_L g3546 ( 
.A1(n_3450),
.A2(n_12),
.B(n_15),
.Y(n_3546)
);

INVx5_ASAP7_75t_L g3547 ( 
.A(n_3382),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3456),
.A2(n_1312),
.B(n_1311),
.Y(n_3548)
);

AOI21xp33_ASAP7_75t_L g3549 ( 
.A1(n_3448),
.A2(n_1882),
.B(n_1881),
.Y(n_3549)
);

AO31x2_ASAP7_75t_L g3550 ( 
.A1(n_3432),
.A2(n_3446),
.A3(n_3460),
.B(n_3409),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3463),
.B(n_1881),
.Y(n_3551)
);

AOI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3424),
.A2(n_16),
.B(n_17),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3372),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3386),
.B(n_1882),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_3462),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3461),
.A2(n_1316),
.B(n_1313),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_3382),
.Y(n_3557)
);

O2A1O1Ixp33_ASAP7_75t_SL g3558 ( 
.A1(n_3496),
.A2(n_47),
.B(n_48),
.C(n_46),
.Y(n_3558)
);

BUFx12f_ASAP7_75t_L g3559 ( 
.A(n_3499),
.Y(n_3559)
);

OAI21x1_ASAP7_75t_L g3560 ( 
.A1(n_3458),
.A2(n_16),
.B(n_17),
.Y(n_3560)
);

BUFx6f_ASAP7_75t_L g3561 ( 
.A(n_3398),
.Y(n_3561)
);

INVx1_ASAP7_75t_SL g3562 ( 
.A(n_3400),
.Y(n_3562)
);

INVx1_ASAP7_75t_SL g3563 ( 
.A(n_3366),
.Y(n_3563)
);

O2A1O1Ixp33_ASAP7_75t_L g3564 ( 
.A1(n_3490),
.A2(n_1511),
.B(n_1654),
.C(n_1504),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3464),
.A2(n_1321),
.B(n_1319),
.Y(n_3565)
);

INVx4_ASAP7_75t_L g3566 ( 
.A(n_3398),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3491),
.A2(n_1324),
.B(n_1323),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3493),
.A2(n_1328),
.B(n_1326),
.Y(n_3568)
);

OAI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3431),
.A2(n_3422),
.B(n_3465),
.Y(n_3569)
);

OAI21x1_ASAP7_75t_L g3570 ( 
.A1(n_3466),
.A2(n_16),
.B(n_18),
.Y(n_3570)
);

A2O1A1Ixp33_ASAP7_75t_L g3571 ( 
.A1(n_3472),
.A2(n_1885),
.B(n_1887),
.C(n_1884),
.Y(n_3571)
);

NAND3x1_ASAP7_75t_L g3572 ( 
.A(n_3498),
.B(n_1667),
.C(n_1654),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3470),
.B(n_3447),
.Y(n_3573)
);

OAI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3483),
.A2(n_1332),
.B(n_1329),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3426),
.A2(n_1334),
.B(n_1333),
.Y(n_3575)
);

OR2x2_ASAP7_75t_L g3576 ( 
.A(n_3412),
.B(n_1884),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3377),
.B(n_1885),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3380),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3439),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3455),
.B(n_1887),
.Y(n_3580)
);

OAI21xp5_ASAP7_75t_SL g3581 ( 
.A1(n_3415),
.A2(n_1667),
.B(n_1654),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_SL g3582 ( 
.A1(n_3485),
.A2(n_1893),
.B(n_1892),
.Y(n_3582)
);

OAI21x1_ASAP7_75t_L g3583 ( 
.A1(n_3471),
.A2(n_18),
.B(n_19),
.Y(n_3583)
);

OAI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3475),
.A2(n_3449),
.B(n_3440),
.Y(n_3584)
);

A2O1A1Ixp33_ASAP7_75t_L g3585 ( 
.A1(n_3392),
.A2(n_1893),
.B(n_1894),
.C(n_1892),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3457),
.B(n_1894),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3467),
.B(n_1899),
.Y(n_3587)
);

NOR2xp33_ASAP7_75t_L g3588 ( 
.A(n_3459),
.B(n_1336),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3442),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3384),
.B(n_1899),
.Y(n_3590)
);

OAI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3425),
.A2(n_19),
.B(n_20),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3371),
.A2(n_1339),
.B(n_1337),
.Y(n_3592)
);

OAI21x1_ASAP7_75t_L g3593 ( 
.A1(n_3469),
.A2(n_20),
.B(n_21),
.Y(n_3593)
);

A2O1A1Ixp33_ASAP7_75t_L g3594 ( 
.A1(n_3405),
.A2(n_1904),
.B(n_1905),
.C(n_1903),
.Y(n_3594)
);

AOI21x1_ASAP7_75t_L g3595 ( 
.A1(n_3403),
.A2(n_20),
.B(n_21),
.Y(n_3595)
);

AOI221xp5_ASAP7_75t_L g3596 ( 
.A1(n_3494),
.A2(n_1346),
.B1(n_1347),
.B2(n_1344),
.C(n_1341),
.Y(n_3596)
);

OAI21x1_ASAP7_75t_L g3597 ( 
.A1(n_3420),
.A2(n_22),
.B(n_23),
.Y(n_3597)
);

NOR2xp67_ASAP7_75t_L g3598 ( 
.A(n_3413),
.B(n_22),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3416),
.A2(n_1350),
.B(n_1349),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3443),
.Y(n_3600)
);

O2A1O1Ixp33_ASAP7_75t_L g3601 ( 
.A1(n_3497),
.A2(n_1678),
.B(n_1786),
.C(n_1667),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3441),
.A2(n_1352),
.B(n_1351),
.Y(n_3602)
);

OAI22xp5_ASAP7_75t_L g3603 ( 
.A1(n_3438),
.A2(n_1904),
.B1(n_1905),
.B2(n_1903),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3376),
.B(n_1678),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3398),
.A2(n_1354),
.B(n_1353),
.Y(n_3605)
);

AOI21x1_ASAP7_75t_SL g3606 ( 
.A1(n_3406),
.A2(n_1786),
.B(n_1678),
.Y(n_3606)
);

NOR2x1_ASAP7_75t_L g3607 ( 
.A(n_3387),
.B(n_1786),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3487),
.B(n_1906),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3428),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3417),
.B(n_1906),
.Y(n_3610)
);

AOI221xp5_ASAP7_75t_L g3611 ( 
.A1(n_3549),
.A2(n_3601),
.B1(n_3534),
.B2(n_3564),
.C(n_3581),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3501),
.A2(n_3527),
.B(n_3513),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3514),
.A2(n_3423),
.B1(n_3451),
.B2(n_3489),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_3525),
.B(n_3393),
.Y(n_3614)
);

INVx5_ASAP7_75t_L g3615 ( 
.A(n_3561),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3521),
.B(n_3430),
.Y(n_3616)
);

OAI21x1_ASAP7_75t_L g3617 ( 
.A1(n_3512),
.A2(n_3473),
.B(n_3411),
.Y(n_3617)
);

OAI21xp33_ASAP7_75t_SL g3618 ( 
.A1(n_3584),
.A2(n_3408),
.B(n_3481),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_SL g3619 ( 
.A1(n_3595),
.A2(n_3486),
.B(n_3468),
.Y(n_3619)
);

CKINVDCx6p67_ASAP7_75t_R g3620 ( 
.A(n_3559),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3518),
.A2(n_3427),
.B(n_3453),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3578),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3509),
.A2(n_3452),
.B(n_1356),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3517),
.A2(n_3453),
.B(n_3390),
.Y(n_3624)
);

OA21x2_ASAP7_75t_L g3625 ( 
.A1(n_3505),
.A2(n_1360),
.B(n_1355),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3502),
.B(n_3454),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3504),
.B(n_3454),
.Y(n_3627)
);

OAI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_3503),
.A2(n_1365),
.B(n_1364),
.Y(n_3628)
);

OAI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3538),
.A2(n_3499),
.B1(n_1908),
.B2(n_1909),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_SL g3630 ( 
.A1(n_3587),
.A2(n_3418),
.B1(n_1908),
.B2(n_1909),
.Y(n_3630)
);

INVx1_ASAP7_75t_SL g3631 ( 
.A(n_3562),
.Y(n_3631)
);

OA21x2_ASAP7_75t_L g3632 ( 
.A1(n_3544),
.A2(n_1369),
.B(n_1367),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3577),
.B(n_3434),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3500),
.B(n_3519),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3563),
.B(n_1372),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3569),
.A2(n_3540),
.B(n_3529),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3528),
.B(n_3402),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_3555),
.Y(n_3638)
);

OAI21x1_ASAP7_75t_L g3639 ( 
.A1(n_3546),
.A2(n_22),
.B(n_23),
.Y(n_3639)
);

AND2x4_ASAP7_75t_L g3640 ( 
.A(n_3532),
.B(n_48),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3553),
.Y(n_3641)
);

BUFx5_ASAP7_75t_L g3642 ( 
.A(n_3579),
.Y(n_3642)
);

HB1xp67_ASAP7_75t_L g3643 ( 
.A(n_3600),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3589),
.Y(n_3644)
);

OAI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3524),
.A2(n_1374),
.B(n_1373),
.Y(n_3645)
);

OA21x2_ASAP7_75t_L g3646 ( 
.A1(n_3560),
.A2(n_1377),
.B(n_1376),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3573),
.B(n_1907),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3545),
.A2(n_3583),
.B(n_3570),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3593),
.A2(n_24),
.B(n_25),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3507),
.B(n_1872),
.Y(n_3650)
);

NAND2xp33_ASAP7_75t_SL g3651 ( 
.A(n_3561),
.B(n_1907),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3508),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3515),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3597),
.A2(n_24),
.B(n_26),
.Y(n_3654)
);

AOI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3552),
.A2(n_1383),
.B(n_1380),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3536),
.Y(n_3656)
);

AO21x2_ASAP7_75t_L g3657 ( 
.A1(n_3591),
.A2(n_1911),
.B(n_1910),
.Y(n_3657)
);

AO21x2_ASAP7_75t_L g3658 ( 
.A1(n_3542),
.A2(n_1911),
.B(n_1910),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3606),
.A2(n_24),
.B(n_26),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3510),
.A2(n_1390),
.B(n_1387),
.Y(n_3660)
);

O2A1O1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3571),
.A2(n_3585),
.B(n_3610),
.C(n_3608),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_L g3662 ( 
.A1(n_3533),
.A2(n_26),
.B(n_27),
.Y(n_3662)
);

OAI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_3520),
.A2(n_1399),
.B1(n_1400),
.B2(n_1392),
.Y(n_3663)
);

NAND2x1p5_ASAP7_75t_L g3664 ( 
.A(n_3547),
.B(n_49),
.Y(n_3664)
);

O2A1O1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_3558),
.A2(n_1859),
.B(n_1862),
.C(n_1857),
.Y(n_3665)
);

CKINVDCx5p33_ASAP7_75t_R g3666 ( 
.A(n_3557),
.Y(n_3666)
);

OAI21x1_ASAP7_75t_L g3667 ( 
.A1(n_3602),
.A2(n_27),
.B(n_28),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3508),
.Y(n_3668)
);

NAND2x1p5_ASAP7_75t_L g3669 ( 
.A(n_3547),
.B(n_50),
.Y(n_3669)
);

OAI21x1_ASAP7_75t_L g3670 ( 
.A1(n_3506),
.A2(n_29),
.B(n_30),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3604),
.B(n_51),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3526),
.B(n_3541),
.Y(n_3672)
);

OAI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3530),
.A2(n_1876),
.B1(n_1877),
.B2(n_1875),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_3609),
.Y(n_3674)
);

OAI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3511),
.A2(n_1879),
.B1(n_1878),
.B2(n_1403),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3536),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3588),
.B(n_3539),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3523),
.Y(n_3678)
);

AOI22xp33_ASAP7_75t_SL g3679 ( 
.A1(n_3574),
.A2(n_1406),
.B1(n_1407),
.B2(n_1402),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3551),
.A2(n_3586),
.B1(n_3603),
.B2(n_3543),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3566),
.B(n_51),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3590),
.A2(n_1410),
.B1(n_1415),
.B2(n_1408),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3598),
.B(n_52),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3523),
.Y(n_3684)
);

NAND2x1p5_ASAP7_75t_L g3685 ( 
.A(n_3607),
.B(n_52),
.Y(n_3685)
);

BUFx2_ASAP7_75t_L g3686 ( 
.A(n_3522),
.Y(n_3686)
);

NOR2x1_ASAP7_75t_SL g3687 ( 
.A(n_3652),
.B(n_3531),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3644),
.Y(n_3688)
);

AO31x2_ASAP7_75t_L g3689 ( 
.A1(n_3656),
.A2(n_3594),
.A3(n_3592),
.B(n_3568),
.Y(n_3689)
);

AO21x2_ASAP7_75t_L g3690 ( 
.A1(n_3616),
.A2(n_3567),
.B(n_3575),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3668),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3678),
.Y(n_3692)
);

OA21x2_ASAP7_75t_L g3693 ( 
.A1(n_3670),
.A2(n_3599),
.B(n_3605),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3625),
.A2(n_3582),
.B(n_3550),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3614),
.B(n_3537),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_3625),
.A2(n_3550),
.B(n_3548),
.Y(n_3696)
);

OR2x2_ASAP7_75t_L g3697 ( 
.A(n_3676),
.B(n_3643),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3674),
.B(n_3626),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3622),
.Y(n_3699)
);

AO21x2_ASAP7_75t_L g3700 ( 
.A1(n_3672),
.A2(n_3565),
.B(n_3556),
.Y(n_3700)
);

OR2x6_ASAP7_75t_L g3701 ( 
.A(n_3624),
.B(n_3572),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3634),
.B(n_3537),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3641),
.Y(n_3703)
);

AOI21xp5_ASAP7_75t_L g3704 ( 
.A1(n_3611),
.A2(n_3580),
.B(n_3596),
.Y(n_3704)
);

AOI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3655),
.A2(n_3535),
.B(n_3516),
.Y(n_3705)
);

CKINVDCx11_ASAP7_75t_R g3706 ( 
.A(n_3620),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3653),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3642),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3684),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3631),
.B(n_3576),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3642),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3686),
.B(n_3554),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3628),
.A2(n_3506),
.B(n_1418),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3612),
.A2(n_29),
.B(n_30),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_3636),
.A2(n_30),
.B(n_31),
.Y(n_3715)
);

AO21x2_ASAP7_75t_L g3716 ( 
.A1(n_3639),
.A2(n_32),
.B(n_33),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3677),
.B(n_3627),
.Y(n_3717)
);

OA21x2_ASAP7_75t_L g3718 ( 
.A1(n_3659),
.A2(n_1419),
.B(n_1416),
.Y(n_3718)
);

OAI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3648),
.A2(n_32),
.B(n_33),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3642),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3642),
.Y(n_3721)
);

OAI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3649),
.A2(n_33),
.B(n_34),
.Y(n_3722)
);

OAI21x1_ASAP7_75t_L g3723 ( 
.A1(n_3654),
.A2(n_34),
.B(n_35),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_3661),
.A2(n_1424),
.B(n_1423),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3617),
.Y(n_3725)
);

OAI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3621),
.A2(n_35),
.B(n_36),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3662),
.Y(n_3727)
);

INVx4_ASAP7_75t_L g3728 ( 
.A(n_3615),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3667),
.Y(n_3729)
);

OA21x2_ASAP7_75t_L g3730 ( 
.A1(n_3619),
.A2(n_3623),
.B(n_3660),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3632),
.Y(n_3731)
);

OA21x2_ASAP7_75t_L g3732 ( 
.A1(n_3645),
.A2(n_1431),
.B(n_1429),
.Y(n_3732)
);

OR2x2_ASAP7_75t_L g3733 ( 
.A(n_3657),
.B(n_53),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3646),
.Y(n_3734)
);

BUFx6f_ASAP7_75t_L g3735 ( 
.A(n_3615),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3637),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3618),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_3680),
.B(n_1438),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3681),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3613),
.B(n_3647),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3683),
.Y(n_3741)
);

OA21x2_ASAP7_75t_L g3742 ( 
.A1(n_3650),
.A2(n_1440),
.B(n_1439),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3671),
.B(n_3635),
.Y(n_3743)
);

BUFx2_ASAP7_75t_L g3744 ( 
.A(n_3695),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3697),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3688),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3691),
.Y(n_3747)
);

HB1xp67_ASAP7_75t_L g3748 ( 
.A(n_3697),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3692),
.Y(n_3749)
);

INVx3_ASAP7_75t_L g3750 ( 
.A(n_3703),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3702),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3699),
.Y(n_3752)
);

OR2x6_ASAP7_75t_L g3753 ( 
.A(n_3701),
.B(n_3664),
.Y(n_3753)
);

HB1xp67_ASAP7_75t_L g3754 ( 
.A(n_3727),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3698),
.B(n_3640),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3709),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3711),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3720),
.Y(n_3758)
);

BUFx3_ASAP7_75t_L g3759 ( 
.A(n_3707),
.Y(n_3759)
);

HB1xp67_ASAP7_75t_L g3760 ( 
.A(n_3729),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3708),
.Y(n_3761)
);

HB1xp67_ASAP7_75t_L g3762 ( 
.A(n_3737),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3721),
.Y(n_3763)
);

BUFx2_ASAP7_75t_L g3764 ( 
.A(n_3728),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3725),
.Y(n_3765)
);

AOI21x1_ASAP7_75t_L g3766 ( 
.A1(n_3701),
.A2(n_3629),
.B(n_3682),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3735),
.Y(n_3767)
);

BUFx6f_ASAP7_75t_L g3768 ( 
.A(n_3735),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3687),
.Y(n_3769)
);

OR2x2_ASAP7_75t_L g3770 ( 
.A(n_3717),
.B(n_3685),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3736),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3734),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3710),
.B(n_3658),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3714),
.Y(n_3774)
);

HB1xp67_ASAP7_75t_L g3775 ( 
.A(n_3731),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3741),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3715),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3719),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3696),
.A2(n_3665),
.B(n_3669),
.Y(n_3779)
);

INVxp33_ASAP7_75t_L g3780 ( 
.A(n_3743),
.Y(n_3780)
);

CKINVDCx20_ASAP7_75t_R g3781 ( 
.A(n_3706),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3739),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3712),
.B(n_3633),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3726),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3716),
.Y(n_3785)
);

OA21x2_ASAP7_75t_L g3786 ( 
.A1(n_3694),
.A2(n_1442),
.B(n_1441),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3740),
.B(n_3673),
.Y(n_3787)
);

AOI21x1_ASAP7_75t_L g3788 ( 
.A1(n_3713),
.A2(n_3663),
.B(n_3679),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3704),
.B(n_3666),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3722),
.Y(n_3790)
);

CKINVDCx20_ASAP7_75t_R g3791 ( 
.A(n_3738),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3700),
.B(n_1443),
.Y(n_3792)
);

OAI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3723),
.A2(n_3693),
.B(n_3718),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3733),
.B(n_3651),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3730),
.B(n_3638),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3733),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3742),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3742),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3689),
.Y(n_3799)
);

INVx2_ASAP7_75t_SL g3800 ( 
.A(n_3690),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3689),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_L g3802 ( 
.A1(n_3705),
.A2(n_3675),
.B(n_35),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3772),
.Y(n_3803)
);

BUFx6f_ASAP7_75t_SL g3804 ( 
.A(n_3753),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3747),
.Y(n_3805)
);

OAI21xp33_ASAP7_75t_L g3806 ( 
.A1(n_3787),
.A2(n_3724),
.B(n_1446),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3747),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3793),
.A2(n_3732),
.B(n_36),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3745),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3749),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3744),
.B(n_3732),
.Y(n_3811)
);

OAI21x1_ASAP7_75t_L g3812 ( 
.A1(n_3799),
.A2(n_3801),
.B(n_3779),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3792),
.A2(n_3630),
.B(n_1447),
.Y(n_3813)
);

OAI211xp5_ASAP7_75t_SL g3814 ( 
.A1(n_3789),
.A2(n_1449),
.B(n_1451),
.C(n_1445),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3780),
.B(n_1453),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_L g3816 ( 
.A1(n_3795),
.A2(n_1850),
.B1(n_1851),
.B2(n_1849),
.Y(n_3816)
);

BUFx3_ASAP7_75t_L g3817 ( 
.A(n_3781),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3748),
.B(n_37),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3745),
.B(n_38),
.Y(n_3819)
);

BUFx2_ASAP7_75t_L g3820 ( 
.A(n_3764),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3749),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3796),
.A2(n_3797),
.B1(n_3798),
.B2(n_3791),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3796),
.A2(n_1457),
.B1(n_1463),
.B2(n_1460),
.Y(n_3823)
);

OAI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3773),
.A2(n_1465),
.B1(n_1468),
.B2(n_1464),
.C(n_1454),
.Y(n_3824)
);

OAI22xp33_ASAP7_75t_L g3825 ( 
.A1(n_3788),
.A2(n_1472),
.B1(n_1474),
.B2(n_1471),
.Y(n_3825)
);

NAND2xp33_ASAP7_75t_R g3826 ( 
.A(n_3753),
.B(n_38),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3786),
.A2(n_1844),
.B1(n_1845),
.B2(n_1843),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3763),
.Y(n_3828)
);

AOI22xp33_ASAP7_75t_L g3829 ( 
.A1(n_3786),
.A2(n_1848),
.B1(n_1852),
.B2(n_1847),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3794),
.A2(n_1854),
.B1(n_1855),
.B2(n_1853),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3751),
.B(n_1475),
.Y(n_3831)
);

BUFx6f_ASAP7_75t_L g3832 ( 
.A(n_3768),
.Y(n_3832)
);

OAI211xp5_ASAP7_75t_L g3833 ( 
.A1(n_3785),
.A2(n_1496),
.B(n_1512),
.C(n_1476),
.Y(n_3833)
);

AOI22xp33_ASAP7_75t_L g3834 ( 
.A1(n_3785),
.A2(n_1479),
.B1(n_1481),
.B2(n_1477),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3762),
.B(n_3782),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3771),
.B(n_1488),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3820),
.B(n_3776),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3805),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3807),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3811),
.B(n_3750),
.Y(n_3840)
);

BUFx2_ASAP7_75t_L g3841 ( 
.A(n_3835),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3809),
.B(n_3828),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3810),
.Y(n_3843)
);

INVx2_ASAP7_75t_SL g3844 ( 
.A(n_3832),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3806),
.A2(n_3790),
.B1(n_3784),
.B2(n_3770),
.Y(n_3845)
);

INVxp67_ASAP7_75t_SL g3846 ( 
.A(n_3821),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3803),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3822),
.B(n_3759),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3812),
.Y(n_3849)
);

INVx4_ASAP7_75t_L g3850 ( 
.A(n_3832),
.Y(n_3850)
);

BUFx2_ASAP7_75t_L g3851 ( 
.A(n_3832),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3825),
.A2(n_3790),
.B1(n_3774),
.B2(n_3777),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3818),
.B(n_3769),
.Y(n_3853)
);

AND2x4_ASAP7_75t_SL g3854 ( 
.A(n_3819),
.B(n_3768),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3817),
.B(n_3755),
.Y(n_3855)
);

AOI22xp5_ASAP7_75t_SL g3856 ( 
.A1(n_3826),
.A2(n_3767),
.B1(n_3768),
.B2(n_3783),
.Y(n_3856)
);

BUFx6f_ASAP7_75t_L g3857 ( 
.A(n_3808),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3836),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3831),
.B(n_3750),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3804),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3816),
.B(n_3761),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3815),
.B(n_3757),
.Y(n_3862)
);

HB1xp67_ASAP7_75t_L g3863 ( 
.A(n_3804),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3823),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3830),
.B(n_3758),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3834),
.B(n_3775),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3824),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3833),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3827),
.B(n_3767),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3863),
.B(n_3746),
.Y(n_3870)
);

NOR2x1p5_ASAP7_75t_L g3871 ( 
.A(n_3860),
.B(n_3766),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3860),
.B(n_3754),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3838),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3858),
.B(n_3752),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3838),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3839),
.Y(n_3876)
);

HB1xp67_ASAP7_75t_L g3877 ( 
.A(n_3846),
.Y(n_3877)
);

OR2x2_ASAP7_75t_L g3878 ( 
.A(n_3841),
.B(n_3778),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3851),
.B(n_3760),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3850),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3848),
.B(n_3765),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3839),
.Y(n_3882)
);

INVxp67_ASAP7_75t_SL g3883 ( 
.A(n_3856),
.Y(n_3883)
);

NAND2x1_ASAP7_75t_SL g3884 ( 
.A(n_3849),
.B(n_3778),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3850),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3843),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3844),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3865),
.B(n_3829),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3847),
.Y(n_3889)
);

NOR2xp33_ASAP7_75t_L g3890 ( 
.A(n_3867),
.B(n_3814),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3842),
.Y(n_3891)
);

OR2x2_ASAP7_75t_L g3892 ( 
.A(n_3840),
.B(n_3800),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_L g3893 ( 
.A1(n_3867),
.A2(n_3868),
.B1(n_3864),
.B2(n_3857),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3857),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3859),
.B(n_3756),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3837),
.B(n_3802),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3857),
.B(n_3813),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3854),
.B(n_38),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_3849),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3862),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3853),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3861),
.B(n_3866),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3845),
.B(n_1491),
.Y(n_3903)
);

OR2x2_ASAP7_75t_L g3904 ( 
.A(n_3852),
.B(n_39),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3877),
.Y(n_3905)
);

NOR2xp67_ASAP7_75t_L g3906 ( 
.A(n_3899),
.B(n_3869),
.Y(n_3906)
);

INVx2_ASAP7_75t_SL g3907 ( 
.A(n_3898),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3873),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3883),
.B(n_3855),
.Y(n_3909)
);

AOI211xp5_ASAP7_75t_L g3910 ( 
.A1(n_3890),
.A2(n_1493),
.B(n_1500),
.C(n_1492),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3887),
.B(n_40),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3900),
.B(n_1498),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3881),
.B(n_40),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3902),
.B(n_1502),
.Y(n_3914)
);

OAI31xp33_ASAP7_75t_SL g3915 ( 
.A1(n_3898),
.A2(n_43),
.A3(n_41),
.B(n_42),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3875),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3880),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3885),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3891),
.B(n_41),
.Y(n_3919)
);

INVxp67_ASAP7_75t_SL g3920 ( 
.A(n_3871),
.Y(n_3920)
);

INVxp67_ASAP7_75t_SL g3921 ( 
.A(n_3897),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3876),
.Y(n_3922)
);

BUFx2_ASAP7_75t_L g3923 ( 
.A(n_3895),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3888),
.A2(n_1871),
.B(n_1508),
.Y(n_3924)
);

AND3x1_ASAP7_75t_L g3925 ( 
.A(n_3893),
.B(n_43),
.C(n_44),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3882),
.Y(n_3926)
);

NAND4xp25_ASAP7_75t_L g3927 ( 
.A(n_3904),
.B(n_44),
.C(n_55),
.D(n_54),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3886),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3870),
.B(n_1506),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3903),
.A2(n_1831),
.B(n_1830),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3874),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3901),
.B(n_44),
.Y(n_3932)
);

NAND4xp25_ASAP7_75t_L g3933 ( 
.A(n_3894),
.B(n_1510),
.C(n_1513),
.D(n_1509),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3884),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3879),
.B(n_54),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3895),
.B(n_56),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3884),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3896),
.B(n_57),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3872),
.Y(n_3939)
);

CKINVDCx16_ASAP7_75t_R g3940 ( 
.A(n_3907),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3938),
.B(n_3889),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_R g3942 ( 
.A(n_3935),
.B(n_57),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3909),
.Y(n_3943)
);

AND2x4_ASAP7_75t_L g3944 ( 
.A(n_3905),
.B(n_3878),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3929),
.B(n_3892),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3939),
.B(n_58),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3920),
.B(n_59),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3908),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3921),
.B(n_60),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3916),
.Y(n_3950)
);

AND2x2_ASAP7_75t_L g3951 ( 
.A(n_3923),
.B(n_61),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3917),
.B(n_1515),
.Y(n_3952)
);

INVx1_ASAP7_75t_SL g3953 ( 
.A(n_3913),
.Y(n_3953)
);

AOI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3924),
.A2(n_1519),
.B(n_1518),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3936),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3918),
.B(n_61),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3922),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3906),
.B(n_63),
.Y(n_3958)
);

OR2x2_ASAP7_75t_L g3959 ( 
.A(n_3931),
.B(n_63),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3926),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3906),
.B(n_1520),
.Y(n_3961)
);

INVx1_ASAP7_75t_SL g3962 ( 
.A(n_3911),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3928),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3919),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3932),
.B(n_3925),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3925),
.B(n_64),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3915),
.B(n_1521),
.Y(n_3967)
);

BUFx2_ASAP7_75t_L g3968 ( 
.A(n_3934),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3914),
.B(n_1526),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3912),
.B(n_64),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3910),
.B(n_1527),
.Y(n_3971)
);

OR2x2_ASAP7_75t_L g3972 ( 
.A(n_3927),
.B(n_65),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_3933),
.B(n_1532),
.Y(n_3973)
);

INVx1_ASAP7_75t_SL g3974 ( 
.A(n_3937),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3933),
.B(n_66),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3910),
.B(n_66),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3930),
.B(n_1535),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3909),
.B(n_67),
.Y(n_3978)
);

OAI33xp33_ASAP7_75t_L g3979 ( 
.A1(n_3928),
.A2(n_1540),
.A3(n_1538),
.B1(n_1541),
.B2(n_1539),
.B3(n_1536),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3909),
.B(n_67),
.Y(n_3980)
);

NOR2xp33_ASAP7_75t_L g3981 ( 
.A(n_3907),
.B(n_1542),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3909),
.B(n_68),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3905),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3909),
.B(n_68),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3905),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3940),
.A2(n_1835),
.B1(n_1837),
.B2(n_1834),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3983),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3943),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3953),
.B(n_69),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3962),
.B(n_3964),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3965),
.B(n_1546),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3947),
.B(n_1547),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3985),
.B(n_69),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3955),
.B(n_1548),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3983),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3963),
.Y(n_3996)
);

OR2x2_ASAP7_75t_L g3997 ( 
.A(n_3949),
.B(n_70),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3963),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3968),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3978),
.B(n_71),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3941),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3966),
.B(n_1549),
.Y(n_4002)
);

INVx2_ASAP7_75t_SL g4003 ( 
.A(n_3944),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3958),
.B(n_1550),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3944),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3948),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3974),
.B(n_72),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3950),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3951),
.B(n_1551),
.Y(n_4009)
);

INVx4_ASAP7_75t_L g4010 ( 
.A(n_3956),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3980),
.B(n_72),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3957),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3960),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3982),
.B(n_74),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3984),
.B(n_1554),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3945),
.B(n_74),
.Y(n_4016)
);

INVxp67_ASAP7_75t_L g4017 ( 
.A(n_3981),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3946),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3970),
.B(n_75),
.Y(n_4019)
);

OR2x2_ASAP7_75t_L g4020 ( 
.A(n_3961),
.B(n_76),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3959),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3976),
.B(n_3967),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3952),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3972),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3969),
.Y(n_4025)
);

NOR2xp33_ASAP7_75t_L g4026 ( 
.A(n_3975),
.B(n_1556),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_L g4027 ( 
.A(n_3942),
.B(n_1557),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3977),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3973),
.B(n_3971),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3954),
.B(n_77),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3979),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3940),
.B(n_78),
.Y(n_4032)
);

INVxp67_ASAP7_75t_L g4033 ( 
.A(n_3965),
.Y(n_4033)
);

OR2x2_ASAP7_75t_L g4034 ( 
.A(n_3953),
.B(n_78),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3940),
.B(n_80),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3940),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3940),
.B(n_81),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3965),
.B(n_1558),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3940),
.B(n_81),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3983),
.Y(n_4040)
);

INVxp67_ASAP7_75t_L g4041 ( 
.A(n_3965),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3940),
.B(n_82),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3983),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3983),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3940),
.B(n_83),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3983),
.Y(n_4046)
);

OR2x2_ASAP7_75t_L g4047 ( 
.A(n_3953),
.B(n_84),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3983),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3983),
.Y(n_4049)
);

INVxp67_ASAP7_75t_L g4050 ( 
.A(n_3965),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3983),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_4036),
.Y(n_4052)
);

OAI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_4003),
.A2(n_1562),
.B1(n_1566),
.B2(n_1561),
.Y(n_4053)
);

OAI221xp5_ASAP7_75t_L g4054 ( 
.A1(n_4033),
.A2(n_1840),
.B1(n_1813),
.B2(n_1573),
.C(n_1575),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_4041),
.B(n_1568),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_4051),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_L g4057 ( 
.A(n_4010),
.B(n_1569),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_4051),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_4050),
.B(n_4032),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3990),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3989),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3987),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3995),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_4035),
.B(n_1581),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_4037),
.B(n_1585),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_4039),
.B(n_1586),
.Y(n_4066)
);

INVxp67_ASAP7_75t_L g4067 ( 
.A(n_4042),
.Y(n_4067)
);

NAND4xp25_ASAP7_75t_L g4068 ( 
.A(n_4024),
.B(n_86),
.C(n_84),
.D(n_85),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_4005),
.A2(n_1591),
.B1(n_1592),
.B2(n_1590),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4040),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4043),
.Y(n_4071)
);

OAI221xp5_ASAP7_75t_L g4072 ( 
.A1(n_4001),
.A2(n_1832),
.B1(n_1805),
.B2(n_1596),
.C(n_1598),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_3999),
.B(n_87),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4045),
.B(n_1593),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4010),
.A2(n_1601),
.B1(n_1602),
.B2(n_1594),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4044),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_4029),
.B(n_1605),
.Y(n_4077)
);

INVx1_ASAP7_75t_SL g4078 ( 
.A(n_4034),
.Y(n_4078)
);

INVxp67_ASAP7_75t_L g4079 ( 
.A(n_4007),
.Y(n_4079)
);

OAI32xp33_ASAP7_75t_L g4080 ( 
.A1(n_4049),
.A2(n_1611),
.A3(n_1612),
.B1(n_1608),
.B2(n_1606),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4046),
.Y(n_4081)
);

OAI221xp5_ASAP7_75t_L g4082 ( 
.A1(n_4021),
.A2(n_1620),
.B1(n_1621),
.B2(n_1619),
.C(n_1613),
.Y(n_4082)
);

OAI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_4022),
.A2(n_4031),
.B(n_3991),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_4018),
.B(n_1624),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_4047),
.Y(n_4085)
);

OAI21xp5_ASAP7_75t_SL g4086 ( 
.A1(n_3986),
.A2(n_91),
.B(n_89),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4048),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3993),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4026),
.B(n_4016),
.Y(n_4089)
);

OAI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3988),
.A2(n_1626),
.B1(n_1627),
.B2(n_1625),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_4017),
.B(n_1628),
.Y(n_4091)
);

NAND2x1p5_ASAP7_75t_L g4092 ( 
.A(n_4000),
.B(n_88),
.Y(n_4092)
);

OAI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_4038),
.A2(n_1630),
.B1(n_1633),
.B2(n_1629),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3996),
.Y(n_4094)
);

NAND3xp33_ASAP7_75t_L g4095 ( 
.A(n_4023),
.B(n_1642),
.C(n_1640),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3998),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_4028),
.B(n_1644),
.Y(n_4097)
);

OAI221xp5_ASAP7_75t_L g4098 ( 
.A1(n_4025),
.A2(n_1820),
.B1(n_1798),
.B2(n_1647),
.C(n_1648),
.Y(n_4098)
);

OAI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_4006),
.A2(n_1646),
.B1(n_1649),
.B2(n_1645),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3997),
.Y(n_4100)
);

AND2x4_ASAP7_75t_L g4101 ( 
.A(n_4008),
.B(n_92),
.Y(n_4101)
);

NOR2xp67_ASAP7_75t_L g4102 ( 
.A(n_4012),
.B(n_91),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4011),
.Y(n_4103)
);

NAND2x1p5_ASAP7_75t_L g4104 ( 
.A(n_4014),
.B(n_94),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4013),
.Y(n_4105)
);

INVxp67_ASAP7_75t_SL g4106 ( 
.A(n_4027),
.Y(n_4106)
);

OR2x2_ASAP7_75t_L g4107 ( 
.A(n_4020),
.B(n_94),
.Y(n_4107)
);

NAND2x1_ASAP7_75t_L g4108 ( 
.A(n_4019),
.B(n_95),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4002),
.B(n_1652),
.Y(n_4109)
);

OAI32xp33_ASAP7_75t_L g4110 ( 
.A1(n_3994),
.A2(n_1657),
.A3(n_1661),
.B1(n_1655),
.B2(n_1653),
.Y(n_4110)
);

INVx1_ASAP7_75t_SL g4111 ( 
.A(n_4030),
.Y(n_4111)
);

AOI322xp5_ASAP7_75t_L g4112 ( 
.A1(n_4004),
.A2(n_1665),
.A3(n_1662),
.B1(n_1669),
.B2(n_1671),
.C1(n_1664),
.C2(n_1660),
.Y(n_4112)
);

AOI211x1_ASAP7_75t_SL g4113 ( 
.A1(n_3992),
.A2(n_98),
.B(n_95),
.C(n_96),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_4009),
.A2(n_1823),
.B(n_1816),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4015),
.B(n_1679),
.Y(n_4115)
);

OA22x2_ASAP7_75t_L g4116 ( 
.A1(n_4033),
.A2(n_1683),
.B1(n_1684),
.B2(n_1680),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4036),
.B(n_1687),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_4033),
.A2(n_1721),
.B(n_1735),
.C(n_1695),
.Y(n_4118)
);

NAND2x1p5_ASAP7_75t_L g4119 ( 
.A(n_4032),
.B(n_99),
.Y(n_4119)
);

INVx1_ASAP7_75t_SL g4120 ( 
.A(n_4032),
.Y(n_4120)
);

AOI222xp33_ASAP7_75t_L g4121 ( 
.A1(n_4033),
.A2(n_1691),
.B1(n_1689),
.B2(n_1693),
.C1(n_1690),
.C2(n_1688),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4033),
.B(n_1694),
.Y(n_4122)
);

OAI33xp33_ASAP7_75t_L g4123 ( 
.A1(n_4033),
.A2(n_1707),
.A3(n_1700),
.B1(n_1708),
.B2(n_1706),
.B3(n_1697),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_4036),
.Y(n_4124)
);

OAI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_4033),
.A2(n_1715),
.B(n_1710),
.Y(n_4125)
);

OAI21xp33_ASAP7_75t_L g4126 ( 
.A1(n_4036),
.A2(n_1726),
.B(n_1722),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_4033),
.B(n_1727),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_4033),
.B(n_99),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_4051),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_4036),
.Y(n_4130)
);

INVx4_ASAP7_75t_L g4131 ( 
.A(n_4032),
.Y(n_4131)
);

NAND2x1p5_ASAP7_75t_L g4132 ( 
.A(n_4032),
.B(n_100),
.Y(n_4132)
);

INVx1_ASAP7_75t_SL g4133 ( 
.A(n_4032),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_4033),
.B(n_1728),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4033),
.B(n_1730),
.Y(n_4135)
);

OAI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_4003),
.A2(n_1732),
.B1(n_1736),
.B2(n_1731),
.Y(n_4136)
);

OR2x2_ASAP7_75t_L g4137 ( 
.A(n_4033),
.B(n_100),
.Y(n_4137)
);

OR2x2_ASAP7_75t_L g4138 ( 
.A(n_4033),
.B(n_101),
.Y(n_4138)
);

OAI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_4033),
.A2(n_1741),
.B1(n_1742),
.B2(n_1740),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_4131),
.B(n_1743),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4102),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4131),
.B(n_1744),
.Y(n_4142)
);

AOI21xp33_ASAP7_75t_SL g4143 ( 
.A1(n_4067),
.A2(n_102),
.B(n_103),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4060),
.Y(n_4144)
);

CKINVDCx20_ASAP7_75t_R g4145 ( 
.A(n_4120),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4119),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4056),
.Y(n_4147)
);

OAI21xp33_ASAP7_75t_L g4148 ( 
.A1(n_4052),
.A2(n_1749),
.B(n_1746),
.Y(n_4148)
);

OAI322xp33_ASAP7_75t_L g4149 ( 
.A1(n_4062),
.A2(n_1753),
.A3(n_1751),
.B1(n_1754),
.B2(n_1755),
.C1(n_1752),
.C2(n_1750),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4058),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4129),
.Y(n_4151)
);

INVxp33_ASAP7_75t_L g4152 ( 
.A(n_4132),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_4133),
.B(n_1756),
.Y(n_4153)
);

OAI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_4068),
.A2(n_1762),
.B1(n_1763),
.B2(n_1757),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4124),
.B(n_4130),
.Y(n_4155)
);

NAND4xp75_ASAP7_75t_L g4156 ( 
.A(n_4059),
.B(n_105),
.C(n_103),
.D(n_104),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4065),
.B(n_4066),
.Y(n_4157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4158 ( 
.A1(n_4061),
.A2(n_107),
.B(n_104),
.C(n_106),
.D(n_108),
.Y(n_4158)
);

INVx3_ASAP7_75t_SL g4159 ( 
.A(n_4073),
.Y(n_4159)
);

AOI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_4083),
.A2(n_1769),
.B(n_1766),
.Y(n_4160)
);

HB1xp67_ASAP7_75t_L g4161 ( 
.A(n_4108),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4103),
.Y(n_4162)
);

AOI31xp33_ASAP7_75t_L g4163 ( 
.A1(n_4078),
.A2(n_1771),
.A3(n_1772),
.B(n_1770),
.Y(n_4163)
);

AOI22xp5_ASAP7_75t_L g4164 ( 
.A1(n_4111),
.A2(n_1775),
.B1(n_1776),
.B2(n_1774),
.Y(n_4164)
);

NAND4xp25_ASAP7_75t_L g4165 ( 
.A(n_4100),
.B(n_4079),
.C(n_4085),
.D(n_4089),
.Y(n_4165)
);

OAI22xp33_ASAP7_75t_SL g4166 ( 
.A1(n_4088),
.A2(n_1815),
.B1(n_1838),
.B2(n_1814),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_4092),
.B(n_1777),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4107),
.Y(n_4168)
);

AOI21xp5_ASAP7_75t_L g4169 ( 
.A1(n_4057),
.A2(n_1782),
.B(n_1780),
.Y(n_4169)
);

AOI221xp5_ASAP7_75t_L g4170 ( 
.A1(n_4063),
.A2(n_1787),
.B1(n_1788),
.B2(n_1785),
.C(n_1783),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4128),
.Y(n_4171)
);

HB1xp67_ASAP7_75t_L g4172 ( 
.A(n_4104),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_4137),
.B(n_1792),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4138),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4117),
.B(n_1793),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4101),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4101),
.Y(n_4177)
);

AOI221xp5_ASAP7_75t_L g4178 ( 
.A1(n_4070),
.A2(n_1803),
.B1(n_1806),
.B2(n_1801),
.C(n_1794),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4097),
.B(n_1807),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4106),
.Y(n_4180)
);

AOI21xp5_ASAP7_75t_L g4181 ( 
.A1(n_4077),
.A2(n_1856),
.B(n_1841),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4071),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4084),
.B(n_1864),
.Y(n_4183)
);

OR2x2_ASAP7_75t_L g4184 ( 
.A(n_4055),
.B(n_106),
.Y(n_4184)
);

OAI32xp33_ASAP7_75t_L g4185 ( 
.A1(n_4113),
.A2(n_1868),
.A3(n_110),
.B1(n_112),
.B2(n_109),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4076),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4116),
.B(n_108),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_SL g4188 ( 
.A(n_4053),
.B(n_111),
.Y(n_4188)
);

OR2x2_ASAP7_75t_L g4189 ( 
.A(n_4122),
.B(n_111),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4086),
.B(n_112),
.Y(n_4190)
);

INVxp67_ASAP7_75t_L g4191 ( 
.A(n_4064),
.Y(n_4191)
);

OAI21xp5_ASAP7_75t_SL g4192 ( 
.A1(n_4121),
.A2(n_1052),
.B(n_1051),
.Y(n_4192)
);

OR2x2_ASAP7_75t_L g4193 ( 
.A(n_4127),
.B(n_113),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4081),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_4074),
.A2(n_4069),
.B1(n_4135),
.B2(n_4134),
.Y(n_4195)
);

NOR2xp33_ASAP7_75t_L g4196 ( 
.A(n_4123),
.B(n_113),
.Y(n_4196)
);

OAI22xp5_ASAP7_75t_L g4197 ( 
.A1(n_4087),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_4105),
.A2(n_117),
.B1(n_114),
.B2(n_115),
.Y(n_4198)
);

AOI21xp33_ASAP7_75t_L g4199 ( 
.A1(n_4136),
.A2(n_1055),
.B(n_1054),
.Y(n_4199)
);

NAND2x1_ASAP7_75t_L g4200 ( 
.A(n_4094),
.B(n_1056),
.Y(n_4200)
);

AOI322xp5_ASAP7_75t_L g4201 ( 
.A1(n_4096),
.A2(n_126),
.A3(n_125),
.B1(n_122),
.B2(n_117),
.C1(n_121),
.C2(n_124),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_4126),
.B(n_122),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4091),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4112),
.B(n_126),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4125),
.B(n_127),
.Y(n_4205)
);

OAI22xp5_ASAP7_75t_L g4206 ( 
.A1(n_4095),
.A2(n_4054),
.B1(n_4072),
.B2(n_4109),
.Y(n_4206)
);

OAI221xp5_ASAP7_75t_L g4207 ( 
.A1(n_4118),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.C(n_132),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4115),
.B(n_131),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_4098),
.B(n_132),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4139),
.Y(n_4210)
);

INVxp33_ASAP7_75t_L g4211 ( 
.A(n_4082),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4075),
.Y(n_4212)
);

OAI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4093),
.A2(n_133),
.B(n_134),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4080),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4090),
.B(n_133),
.Y(n_4215)
);

INVxp67_ASAP7_75t_SL g4216 ( 
.A(n_4099),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4110),
.B(n_4114),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4102),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4102),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4102),
.Y(n_4220)
);

XNOR2x1_ASAP7_75t_L g4221 ( 
.A(n_4120),
.B(n_134),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4131),
.B(n_135),
.Y(n_4222)
);

AOI22xp33_ASAP7_75t_SL g4223 ( 
.A1(n_4131),
.A2(n_141),
.B1(n_136),
.B2(n_139),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4102),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_4131),
.B(n_139),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_4052),
.A2(n_146),
.B1(n_142),
.B2(n_144),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4131),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4131),
.B(n_142),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_L g4229 ( 
.A1(n_4052),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_4229)
);

NAND2x1_ASAP7_75t_L g4230 ( 
.A(n_4131),
.B(n_1062),
.Y(n_4230)
);

OR2x2_ASAP7_75t_L g4231 ( 
.A(n_4120),
.B(n_147),
.Y(n_4231)
);

XNOR2xp5_ASAP7_75t_L g4232 ( 
.A(n_4120),
.B(n_1041),
.Y(n_4232)
);

OA222x2_ASAP7_75t_L g4233 ( 
.A1(n_4056),
.A2(n_150),
.B1(n_152),
.B2(n_148),
.C1(n_149),
.C2(n_151),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4083),
.A2(n_150),
.B(n_151),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4102),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4102),
.Y(n_4236)
);

NAND4xp25_ASAP7_75t_SL g4237 ( 
.A(n_4120),
.B(n_154),
.C(n_152),
.D(n_153),
.Y(n_4237)
);

AOI322xp5_ASAP7_75t_L g4238 ( 
.A1(n_4120),
.A2(n_161),
.A3(n_158),
.B1(n_155),
.B2(n_153),
.C1(n_154),
.C2(n_157),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_4131),
.B(n_161),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_L g4240 ( 
.A(n_4131),
.B(n_162),
.Y(n_4240)
);

AOI221xp5_ASAP7_75t_L g4241 ( 
.A1(n_4083),
.A2(n_184),
.B1(n_194),
.B2(n_173),
.C(n_162),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4102),
.Y(n_4242)
);

OR2x2_ASAP7_75t_L g4243 ( 
.A(n_4120),
.B(n_163),
.Y(n_4243)
);

INVx1_ASAP7_75t_SL g4244 ( 
.A(n_4120),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_4131),
.A2(n_167),
.B1(n_164),
.B2(n_166),
.Y(n_4245)
);

HB1xp67_ASAP7_75t_L g4246 ( 
.A(n_4102),
.Y(n_4246)
);

AOI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_4052),
.A2(n_171),
.B1(n_167),
.B2(n_169),
.Y(n_4247)
);

OR2x2_ASAP7_75t_L g4248 ( 
.A(n_4120),
.B(n_171),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4052),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_4249)
);

AOI322xp5_ASAP7_75t_L g4250 ( 
.A1(n_4120),
.A2(n_178),
.A3(n_177),
.B1(n_175),
.B2(n_172),
.C1(n_174),
.C2(n_176),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4131),
.B(n_177),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4131),
.B(n_179),
.Y(n_4252)
);

OAI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_4131),
.A2(n_186),
.B1(n_180),
.B2(n_184),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4102),
.Y(n_4254)
);

OAI221xp5_ASAP7_75t_L g4255 ( 
.A1(n_4083),
.A2(n_187),
.B1(n_180),
.B2(n_186),
.C(n_188),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_4052),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4102),
.Y(n_4257)
);

AOI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_4052),
.A2(n_194),
.B1(n_191),
.B2(n_192),
.Y(n_4258)
);

OAI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_4131),
.A2(n_196),
.B1(n_191),
.B2(n_195),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4131),
.A2(n_199),
.B1(n_195),
.B2(n_197),
.Y(n_4260)
);

NAND2x1_ASAP7_75t_L g4261 ( 
.A(n_4131),
.B(n_1052),
.Y(n_4261)
);

AOI211x1_ASAP7_75t_L g4262 ( 
.A1(n_4083),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_4262)
);

OAI21xp33_ASAP7_75t_SL g4263 ( 
.A1(n_4131),
.A2(n_203),
.B(n_204),
.Y(n_4263)
);

AOI31xp33_ASAP7_75t_L g4264 ( 
.A1(n_4120),
.A2(n_205),
.A3(n_203),
.B(n_204),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4131),
.B(n_206),
.Y(n_4265)
);

NOR2xp33_ASAP7_75t_SL g4266 ( 
.A(n_4131),
.B(n_207),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_SL g4267 ( 
.A(n_4131),
.B(n_207),
.Y(n_4267)
);

OR2x2_ASAP7_75t_L g4268 ( 
.A(n_4120),
.B(n_208),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4102),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4083),
.A2(n_208),
.B(n_209),
.Y(n_4270)
);

NOR2xp33_ASAP7_75t_L g4271 ( 
.A(n_4131),
.B(n_209),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4131),
.B(n_210),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4102),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4102),
.Y(n_4274)
);

BUFx2_ASAP7_75t_L g4275 ( 
.A(n_4131),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4131),
.B(n_210),
.Y(n_4276)
);

NAND2xp33_ASAP7_75t_SL g4277 ( 
.A(n_4108),
.B(n_212),
.Y(n_4277)
);

OAI211xp5_ASAP7_75t_SL g4278 ( 
.A1(n_4083),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_4102),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4120),
.B(n_211),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4131),
.B(n_214),
.Y(n_4281)
);

OAI22xp5_ASAP7_75t_L g4282 ( 
.A1(n_4131),
.A2(n_220),
.B1(n_215),
.B2(n_218),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4102),
.Y(n_4283)
);

XNOR2xp5_ASAP7_75t_L g4284 ( 
.A(n_4120),
.B(n_1057),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4102),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_4131),
.B(n_218),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4131),
.B(n_221),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4131),
.B(n_222),
.Y(n_4288)
);

OAI22xp33_ASAP7_75t_L g4289 ( 
.A1(n_4120),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_4289)
);

OAI21xp33_ASAP7_75t_SL g4290 ( 
.A1(n_4131),
.A2(n_223),
.B(n_225),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4244),
.B(n_226),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4275),
.B(n_227),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4145),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4230),
.Y(n_4294)
);

HB1xp67_ASAP7_75t_L g4295 ( 
.A(n_4246),
.Y(n_4295)
);

AOI221xp5_ASAP7_75t_SL g4296 ( 
.A1(n_4185),
.A2(n_4270),
.B1(n_4234),
.B2(n_4264),
.C(n_4144),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4279),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4161),
.B(n_227),
.Y(n_4298)
);

OAI22xp5_ASAP7_75t_L g4299 ( 
.A1(n_4152),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_4299)
);

AOI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4277),
.A2(n_1048),
.B1(n_1050),
.B2(n_1047),
.Y(n_4300)
);

INVxp67_ASAP7_75t_SL g4301 ( 
.A(n_4261),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_4227),
.B(n_230),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4141),
.Y(n_4303)
);

AOI21xp33_ASAP7_75t_SL g4304 ( 
.A1(n_4159),
.A2(n_4221),
.B(n_4163),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4218),
.Y(n_4305)
);

OR2x2_ASAP7_75t_L g4306 ( 
.A(n_4219),
.B(n_232),
.Y(n_4306)
);

OAI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_4155),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4220),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4224),
.Y(n_4309)
);

AOI322xp5_ASAP7_75t_L g4310 ( 
.A1(n_4216),
.A2(n_239),
.A3(n_238),
.B1(n_236),
.B2(n_234),
.C1(n_235),
.C2(n_237),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4235),
.Y(n_4311)
);

AOI22xp5_ASAP7_75t_L g4312 ( 
.A1(n_4146),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.Y(n_4312)
);

O2A1O1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_4158),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_4165),
.A2(n_1042),
.B1(n_1043),
.B2(n_1040),
.Y(n_4314)
);

AOI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4172),
.A2(n_1044),
.B1(n_1045),
.B2(n_1042),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_4236),
.B(n_241),
.Y(n_4316)
);

NAND3xp33_ASAP7_75t_L g4317 ( 
.A(n_4242),
.B(n_243),
.C(n_244),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_SL g4318 ( 
.A1(n_4254),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4176),
.B(n_246),
.Y(n_4319)
);

AO22x1_ASAP7_75t_L g4320 ( 
.A1(n_4257),
.A2(n_256),
.B1(n_265),
.B2(n_248),
.Y(n_4320)
);

NOR4xp25_ASAP7_75t_SL g4321 ( 
.A(n_4269),
.B(n_251),
.C(n_252),
.D(n_250),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4273),
.Y(n_4322)
);

AOI221xp5_ASAP7_75t_L g4323 ( 
.A1(n_4262),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_253),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4274),
.B(n_249),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4283),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4177),
.B(n_253),
.Y(n_4326)
);

AOI21xp33_ASAP7_75t_SL g4327 ( 
.A1(n_4285),
.A2(n_1037),
.B(n_1036),
.Y(n_4327)
);

AOI321xp33_ASAP7_75t_L g4328 ( 
.A1(n_4180),
.A2(n_1044),
.A3(n_1038),
.B1(n_1045),
.B2(n_1039),
.C(n_1037),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4251),
.B(n_254),
.Y(n_4329)
);

O2A1O1Ixp33_ASAP7_75t_SL g4330 ( 
.A1(n_4200),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4168),
.B(n_255),
.Y(n_4331)
);

HB1xp67_ASAP7_75t_L g4332 ( 
.A(n_4265),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4272),
.B(n_257),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4287),
.B(n_257),
.Y(n_4334)
);

NOR2xp33_ASAP7_75t_L g4335 ( 
.A(n_4266),
.B(n_258),
.Y(n_4335)
);

AOI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4278),
.A2(n_1061),
.B1(n_261),
.B2(n_259),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4222),
.Y(n_4337)
);

NAND2x1p5_ASAP7_75t_L g4338 ( 
.A(n_4167),
.B(n_260),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4231),
.B(n_259),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4228),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4171),
.B(n_263),
.Y(n_4341)
);

NOR3xp33_ASAP7_75t_L g4342 ( 
.A(n_4157),
.B(n_264),
.C(n_267),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4239),
.Y(n_4343)
);

AOI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_4192),
.A2(n_1032),
.B1(n_1033),
.B2(n_1031),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4255),
.A2(n_270),
.B1(n_267),
.B2(n_269),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4252),
.Y(n_4346)
);

OAI21xp33_ASAP7_75t_L g4347 ( 
.A1(n_4211),
.A2(n_270),
.B(n_271),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4262),
.B(n_4232),
.Y(n_4348)
);

OAI221xp5_ASAP7_75t_SL g4349 ( 
.A1(n_4241),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.C(n_275),
.Y(n_4349)
);

OAI221xp5_ASAP7_75t_L g4350 ( 
.A1(n_4162),
.A2(n_1053),
.B1(n_1059),
.B2(n_1051),
.C(n_1048),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4243),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4248),
.B(n_272),
.Y(n_4352)
);

AO22x1_ASAP7_75t_L g4353 ( 
.A1(n_4233),
.A2(n_283),
.B1(n_294),
.B2(n_274),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4284),
.B(n_275),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4276),
.Y(n_4355)
);

INVxp67_ASAP7_75t_L g4356 ( 
.A(n_4240),
.Y(n_4356)
);

OAI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4226),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_4357)
);

OAI32xp33_ASAP7_75t_L g4358 ( 
.A1(n_4263),
.A2(n_297),
.A3(n_307),
.B1(n_288),
.B2(n_277),
.Y(n_4358)
);

OAI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_4190),
.A2(n_281),
.B1(n_278),
.B2(n_280),
.Y(n_4359)
);

AOI221x1_ASAP7_75t_L g4360 ( 
.A1(n_4166),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.C(n_283),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4281),
.Y(n_4361)
);

INVx1_ASAP7_75t_SL g4362 ( 
.A(n_4268),
.Y(n_4362)
);

AOI21xp33_ASAP7_75t_L g4363 ( 
.A1(n_4212),
.A2(n_4210),
.B(n_4174),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4143),
.B(n_282),
.Y(n_4364)
);

OAI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_4229),
.A2(n_288),
.B1(n_285),
.B2(n_287),
.Y(n_4365)
);

AOI21xp33_ASAP7_75t_L g4366 ( 
.A1(n_4195),
.A2(n_285),
.B(n_287),
.Y(n_4366)
);

OAI22xp5_ASAP7_75t_L g4367 ( 
.A1(n_4256),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_4290),
.B(n_293),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4288),
.Y(n_4369)
);

OAI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4223),
.A2(n_4198),
.B1(n_4204),
.B2(n_4214),
.Y(n_4370)
);

OAI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_4247),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4371)
);

OAI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4249),
.A2(n_298),
.B1(n_295),
.B2(n_296),
.Y(n_4372)
);

AND2x2_ASAP7_75t_L g4373 ( 
.A(n_4217),
.B(n_296),
.Y(n_4373)
);

OAI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4258),
.A2(n_301),
.B1(n_298),
.B2(n_300),
.Y(n_4374)
);

OA21x2_ASAP7_75t_L g4375 ( 
.A1(n_4147),
.A2(n_301),
.B(n_303),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4280),
.Y(n_4376)
);

OAI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4207),
.A2(n_4289),
.B1(n_4215),
.B2(n_4164),
.Y(n_4377)
);

OAI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4245),
.A2(n_4259),
.B1(n_4260),
.B2(n_4253),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4271),
.Y(n_4379)
);

OAI22xp33_ASAP7_75t_L g4380 ( 
.A1(n_4282),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_4160),
.A2(n_304),
.B(n_306),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4286),
.Y(n_4382)
);

INVxp67_ASAP7_75t_L g4383 ( 
.A(n_4225),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4237),
.B(n_307),
.Y(n_4384)
);

AOI221xp5_ASAP7_75t_L g4385 ( 
.A1(n_4182),
.A2(n_1035),
.B1(n_1039),
.B2(n_1034),
.C(n_1032),
.Y(n_4385)
);

AOI22xp5_ASAP7_75t_L g4386 ( 
.A1(n_4188),
.A2(n_1059),
.B1(n_1060),
.B2(n_1053),
.Y(n_4386)
);

AOI222xp33_ASAP7_75t_L g4387 ( 
.A1(n_4267),
.A2(n_310),
.B1(n_312),
.B2(n_308),
.C1(n_309),
.C2(n_311),
.Y(n_4387)
);

OAI21xp33_ASAP7_75t_SL g4388 ( 
.A1(n_4150),
.A2(n_308),
.B(n_309),
.Y(n_4388)
);

INVxp67_ASAP7_75t_L g4389 ( 
.A(n_4156),
.Y(n_4389)
);

INVx2_ASAP7_75t_SL g4390 ( 
.A(n_4186),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4184),
.Y(n_4391)
);

OAI31xp33_ASAP7_75t_L g4392 ( 
.A1(n_4197),
.A2(n_314),
.A3(n_310),
.B(n_313),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4189),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4193),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_4187),
.B(n_313),
.Y(n_4395)
);

OAI211xp5_ASAP7_75t_SL g4396 ( 
.A1(n_4191),
.A2(n_317),
.B(n_314),
.C(n_315),
.Y(n_4396)
);

NAND4xp25_ASAP7_75t_SL g4397 ( 
.A(n_4238),
.B(n_318),
.C(n_315),
.D(n_317),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4153),
.B(n_318),
.Y(n_4398)
);

OAI31xp33_ASAP7_75t_L g4399 ( 
.A1(n_4154),
.A2(n_323),
.A3(n_319),
.B(n_322),
.Y(n_4399)
);

NOR3xp33_ASAP7_75t_L g4400 ( 
.A(n_4206),
.B(n_319),
.C(n_322),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4196),
.B(n_323),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4203),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_4402)
);

NOR3xp33_ASAP7_75t_L g4403 ( 
.A(n_4148),
.B(n_326),
.C(n_327),
.Y(n_4403)
);

INVxp67_ASAP7_75t_L g4404 ( 
.A(n_4173),
.Y(n_4404)
);

BUFx2_ASAP7_75t_L g4405 ( 
.A(n_4194),
.Y(n_4405)
);

AOI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4209),
.A2(n_1061),
.B1(n_330),
.B2(n_328),
.Y(n_4406)
);

NAND2x1_ASAP7_75t_L g4407 ( 
.A(n_4151),
.B(n_328),
.Y(n_4407)
);

INVx1_ASAP7_75t_SL g4408 ( 
.A(n_4205),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4175),
.A2(n_332),
.B1(n_329),
.B2(n_331),
.Y(n_4409)
);

AOI22xp5_ASAP7_75t_L g4410 ( 
.A1(n_4202),
.A2(n_1022),
.B1(n_1023),
.B2(n_1021),
.Y(n_4410)
);

OAI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_4313),
.A2(n_4250),
.B(n_4213),
.Y(n_4411)
);

AOI321xp33_ASAP7_75t_L g4412 ( 
.A1(n_4297),
.A2(n_4199),
.A3(n_4142),
.B1(n_4140),
.B2(n_4178),
.C(n_4170),
.Y(n_4412)
);

OAI21xp33_ASAP7_75t_L g4413 ( 
.A1(n_4293),
.A2(n_4208),
.B(n_4179),
.Y(n_4413)
);

AOI211xp5_ASAP7_75t_SL g4414 ( 
.A1(n_4363),
.A2(n_4301),
.B(n_4389),
.C(n_4383),
.Y(n_4414)
);

NAND4xp25_ASAP7_75t_L g4415 ( 
.A(n_4296),
.B(n_4201),
.C(n_4183),
.D(n_4181),
.Y(n_4415)
);

AOI221xp5_ASAP7_75t_L g4416 ( 
.A1(n_4370),
.A2(n_4149),
.B1(n_4169),
.B2(n_335),
.C(n_333),
.Y(n_4416)
);

AOI221xp5_ASAP7_75t_L g4417 ( 
.A1(n_4378),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_4417)
);

AOI322xp5_ASAP7_75t_L g4418 ( 
.A1(n_4348),
.A2(n_1034),
.A3(n_1023),
.B1(n_342),
.B2(n_338),
.C1(n_340),
.C2(n_336),
.Y(n_4418)
);

AOI221x1_ASAP7_75t_L g4419 ( 
.A1(n_4304),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.C(n_342),
.Y(n_4419)
);

AOI21xp5_ASAP7_75t_L g4420 ( 
.A1(n_4353),
.A2(n_337),
.B(n_344),
.Y(n_4420)
);

AOI211xp5_ASAP7_75t_L g4421 ( 
.A1(n_4377),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_4421)
);

INVxp67_ASAP7_75t_L g4422 ( 
.A(n_4295),
.Y(n_4422)
);

AOI221xp5_ASAP7_75t_L g4423 ( 
.A1(n_4397),
.A2(n_348),
.B1(n_345),
.B2(n_347),
.C(n_349),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_4294),
.B(n_351),
.Y(n_4424)
);

NOR3xp33_ASAP7_75t_L g4425 ( 
.A(n_4356),
.B(n_354),
.C(n_356),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4320),
.B(n_4332),
.Y(n_4426)
);

OAI21xp5_ASAP7_75t_L g4427 ( 
.A1(n_4388),
.A2(n_357),
.B(n_359),
.Y(n_4427)
);

OAI211xp5_ASAP7_75t_L g4428 ( 
.A1(n_4328),
.A2(n_362),
.B(n_359),
.C(n_361),
.Y(n_4428)
);

AOI21xp5_ASAP7_75t_L g4429 ( 
.A1(n_4401),
.A2(n_361),
.B(n_362),
.Y(n_4429)
);

OAI22xp5_ASAP7_75t_L g4430 ( 
.A1(n_4344),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4292),
.Y(n_4431)
);

OAI221xp5_ASAP7_75t_L g4432 ( 
.A1(n_4303),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.C(n_370),
.Y(n_4432)
);

AOI31xp33_ASAP7_75t_L g4433 ( 
.A1(n_4362),
.A2(n_373),
.A3(n_371),
.B(n_372),
.Y(n_4433)
);

OAI21xp33_ASAP7_75t_L g4434 ( 
.A1(n_4408),
.A2(n_371),
.B(n_373),
.Y(n_4434)
);

AOI211xp5_ASAP7_75t_L g4435 ( 
.A1(n_4358),
.A2(n_1020),
.B(n_1021),
.C(n_1019),
.Y(n_4435)
);

NAND3xp33_ASAP7_75t_L g4436 ( 
.A(n_4305),
.B(n_4309),
.C(n_4308),
.Y(n_4436)
);

OAI221xp5_ASAP7_75t_L g4437 ( 
.A1(n_4311),
.A2(n_379),
.B1(n_376),
.B2(n_377),
.C(n_382),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_4330),
.A2(n_379),
.B(n_382),
.Y(n_4438)
);

OAI21xp5_ASAP7_75t_SL g4439 ( 
.A1(n_4373),
.A2(n_384),
.B(n_385),
.Y(n_4439)
);

O2A1O1Ixp33_ASAP7_75t_SL g4440 ( 
.A1(n_4407),
.A2(n_388),
.B(n_386),
.C(n_387),
.Y(n_4440)
);

OAI221xp5_ASAP7_75t_L g4441 ( 
.A1(n_4322),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.C(n_391),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4319),
.B(n_390),
.Y(n_4442)
);

NOR2xp33_ASAP7_75t_L g4443 ( 
.A(n_4368),
.B(n_393),
.Y(n_4443)
);

AOI211xp5_ASAP7_75t_L g4444 ( 
.A1(n_4349),
.A2(n_1016),
.B(n_1018),
.C(n_1015),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_4298),
.A2(n_396),
.B(n_397),
.Y(n_4445)
);

OR2x2_ASAP7_75t_L g4446 ( 
.A(n_4325),
.B(n_396),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4326),
.B(n_398),
.Y(n_4447)
);

AOI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_4400),
.A2(n_402),
.B1(n_399),
.B2(n_400),
.Y(n_4448)
);

AOI211xp5_ASAP7_75t_L g4449 ( 
.A1(n_4323),
.A2(n_1022),
.B(n_1024),
.C(n_1020),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4316),
.A2(n_399),
.B(n_400),
.Y(n_4450)
);

AOI221xp5_ASAP7_75t_L g4451 ( 
.A1(n_4405),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.C(n_405),
.Y(n_4451)
);

OAI221xp5_ASAP7_75t_SL g4452 ( 
.A1(n_4310),
.A2(n_1031),
.B1(n_1030),
.B2(n_1028),
.C(n_406),
.Y(n_4452)
);

NAND4xp25_ASAP7_75t_L g4453 ( 
.A(n_4376),
.B(n_406),
.C(n_403),
.D(n_405),
.Y(n_4453)
);

NOR4xp25_ASAP7_75t_L g4454 ( 
.A(n_4390),
.B(n_411),
.C(n_407),
.D(n_409),
.Y(n_4454)
);

HB1xp67_ASAP7_75t_L g4455 ( 
.A(n_4375),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_4327),
.B(n_407),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4291),
.B(n_409),
.Y(n_4457)
);

OAI21xp33_ASAP7_75t_L g4458 ( 
.A1(n_4393),
.A2(n_411),
.B(n_412),
.Y(n_4458)
);

AOI311xp33_ASAP7_75t_L g4459 ( 
.A1(n_4337),
.A2(n_414),
.A3(n_412),
.B(n_413),
.C(n_415),
.Y(n_4459)
);

AOI22xp5_ASAP7_75t_L g4460 ( 
.A1(n_4342),
.A2(n_416),
.B1(n_413),
.B2(n_415),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4314),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4318),
.B(n_418),
.Y(n_4462)
);

AOI322xp5_ASAP7_75t_L g4463 ( 
.A1(n_4359),
.A2(n_1025),
.A3(n_426),
.B1(n_423),
.B2(n_425),
.C1(n_421),
.C2(n_422),
.Y(n_4463)
);

AOI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_4345),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4464)
);

AOI211xp5_ASAP7_75t_SL g4465 ( 
.A1(n_4379),
.A2(n_427),
.B(n_424),
.C(n_426),
.Y(n_4465)
);

OAI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_4336),
.A2(n_431),
.B1(n_428),
.B2(n_429),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4324),
.A2(n_428),
.B(n_431),
.Y(n_4467)
);

NAND3xp33_ASAP7_75t_SL g4468 ( 
.A(n_4321),
.B(n_435),
.C(n_433),
.Y(n_4468)
);

O2A1O1Ixp33_ASAP7_75t_L g4469 ( 
.A1(n_4396),
.A2(n_435),
.B(n_432),
.C(n_433),
.Y(n_4469)
);

A2O1A1Ixp33_ASAP7_75t_L g4470 ( 
.A1(n_4392),
.A2(n_445),
.B(n_454),
.C(n_432),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4381),
.A2(n_436),
.B(n_437),
.Y(n_4471)
);

AOI211xp5_ASAP7_75t_SL g4472 ( 
.A1(n_4382),
.A2(n_441),
.B(n_436),
.C(n_440),
.Y(n_4472)
);

OAI321xp33_ASAP7_75t_L g4473 ( 
.A1(n_4340),
.A2(n_443),
.A3(n_445),
.B1(n_441),
.B2(n_442),
.C(n_444),
.Y(n_4473)
);

OAI31xp33_ASAP7_75t_L g4474 ( 
.A1(n_4371),
.A2(n_446),
.A3(n_442),
.B(n_443),
.Y(n_4474)
);

AO21x1_ASAP7_75t_L g4475 ( 
.A1(n_4384),
.A2(n_1016),
.B(n_1006),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4300),
.B(n_446),
.Y(n_4476)
);

OAI221xp5_ASAP7_75t_L g4477 ( 
.A1(n_4399),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.C(n_451),
.Y(n_4477)
);

OAI222xp33_ASAP7_75t_L g4478 ( 
.A1(n_4351),
.A2(n_1018),
.B1(n_1013),
.B2(n_1019),
.C1(n_1014),
.C2(n_1012),
.Y(n_4478)
);

AOI211xp5_ASAP7_75t_L g4479 ( 
.A1(n_4366),
.A2(n_1014),
.B(n_1025),
.C(n_1013),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4306),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_4386),
.A2(n_453),
.B1(n_448),
.B2(n_452),
.Y(n_4481)
);

NOR2xp67_ASAP7_75t_L g4482 ( 
.A(n_4317),
.B(n_452),
.Y(n_4482)
);

AOI222xp33_ASAP7_75t_L g4483 ( 
.A1(n_4343),
.A2(n_455),
.B1(n_457),
.B2(n_453),
.C1(n_454),
.C2(n_456),
.Y(n_4483)
);

OAI21xp33_ASAP7_75t_L g4484 ( 
.A1(n_4404),
.A2(n_4394),
.B(n_4391),
.Y(n_4484)
);

AOI222xp33_ASAP7_75t_L g4485 ( 
.A1(n_4346),
.A2(n_458),
.B1(n_460),
.B2(n_455),
.C1(n_457),
.C2(n_459),
.Y(n_4485)
);

OAI221xp5_ASAP7_75t_L g4486 ( 
.A1(n_4347),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.C(n_461),
.Y(n_4486)
);

OAI21xp33_ASAP7_75t_SL g4487 ( 
.A1(n_4355),
.A2(n_462),
.B(n_463),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4375),
.Y(n_4488)
);

AOI321xp33_ASAP7_75t_L g4489 ( 
.A1(n_4361),
.A2(n_466),
.A3(n_468),
.B1(n_464),
.B2(n_465),
.C(n_467),
.Y(n_4489)
);

AOI22xp5_ASAP7_75t_L g4490 ( 
.A1(n_4403),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_4490)
);

NAND3xp33_ASAP7_75t_L g4491 ( 
.A(n_4360),
.B(n_470),
.C(n_471),
.Y(n_4491)
);

AOI22xp5_ASAP7_75t_L g4492 ( 
.A1(n_4331),
.A2(n_474),
.B1(n_470),
.B2(n_473),
.Y(n_4492)
);

OAI221xp5_ASAP7_75t_SL g4493 ( 
.A1(n_4369),
.A2(n_1001),
.B1(n_1002),
.B2(n_998),
.C(n_997),
.Y(n_4493)
);

OA22x2_ASAP7_75t_L g4494 ( 
.A1(n_4406),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_4494)
);

OAI221xp5_ASAP7_75t_L g4495 ( 
.A1(n_4385),
.A2(n_478),
.B1(n_475),
.B2(n_476),
.C(n_480),
.Y(n_4495)
);

OAI21xp5_ASAP7_75t_SL g4496 ( 
.A1(n_4387),
.A2(n_481),
.B(n_482),
.Y(n_4496)
);

AOI22xp5_ASAP7_75t_L g4497 ( 
.A1(n_4341),
.A2(n_4357),
.B1(n_4367),
.B2(n_4365),
.Y(n_4497)
);

AOI22xp5_ASAP7_75t_L g4498 ( 
.A1(n_4372),
.A2(n_488),
.B1(n_484),
.B2(n_485),
.Y(n_4498)
);

OR2x2_ASAP7_75t_L g4499 ( 
.A(n_4339),
.B(n_489),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_4395),
.A2(n_490),
.B(n_491),
.Y(n_4500)
);

AOI221x1_ASAP7_75t_L g4501 ( 
.A1(n_4299),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.C(n_495),
.Y(n_4501)
);

O2A1O1Ixp33_ASAP7_75t_L g4502 ( 
.A1(n_4307),
.A2(n_497),
.B(n_493),
.C(n_496),
.Y(n_4502)
);

AOI322xp5_ASAP7_75t_L g4503 ( 
.A1(n_4335),
.A2(n_1012),
.A3(n_998),
.B1(n_501),
.B2(n_498),
.C1(n_500),
.C2(n_496),
.Y(n_4503)
);

AOI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_4364),
.A2(n_497),
.B(n_499),
.Y(n_4504)
);

NAND2x1_ASAP7_75t_SL g4505 ( 
.A(n_4315),
.B(n_499),
.Y(n_4505)
);

NOR2xp33_ASAP7_75t_L g4506 ( 
.A(n_4329),
.B(n_500),
.Y(n_4506)
);

AOI211xp5_ASAP7_75t_L g4507 ( 
.A1(n_4380),
.A2(n_1026),
.B(n_1027),
.C(n_1011),
.Y(n_4507)
);

NOR3xp33_ASAP7_75t_L g4508 ( 
.A(n_4398),
.B(n_501),
.C(n_502),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4338),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4410),
.A2(n_506),
.B1(n_503),
.B2(n_504),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4352),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4333),
.B(n_503),
.Y(n_4512)
);

OAI22xp5_ASAP7_75t_L g4513 ( 
.A1(n_4312),
.A2(n_507),
.B1(n_504),
.B2(n_506),
.Y(n_4513)
);

AOI221xp5_ASAP7_75t_L g4514 ( 
.A1(n_4374),
.A2(n_4409),
.B1(n_4350),
.B2(n_4402),
.C(n_4354),
.Y(n_4514)
);

O2A1O1Ixp33_ASAP7_75t_L g4515 ( 
.A1(n_4302),
.A2(n_512),
.B(n_507),
.C(n_509),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4334),
.B(n_509),
.Y(n_4516)
);

AOI222xp33_ASAP7_75t_L g4517 ( 
.A1(n_4370),
.A2(n_515),
.B1(n_518),
.B2(n_513),
.C1(n_514),
.C2(n_516),
.Y(n_4517)
);

AOI221xp5_ASAP7_75t_L g4518 ( 
.A1(n_4370),
.A2(n_518),
.B1(n_513),
.B2(n_516),
.C(n_522),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4353),
.B(n_522),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_SL g4520 ( 
.A(n_4294),
.B(n_524),
.Y(n_4520)
);

AOI221xp5_ASAP7_75t_L g4521 ( 
.A1(n_4370),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.C(n_527),
.Y(n_4521)
);

NAND4xp25_ASAP7_75t_SL g4522 ( 
.A(n_4313),
.B(n_528),
.C(n_525),
.D(n_526),
.Y(n_4522)
);

AOI221xp5_ASAP7_75t_L g4523 ( 
.A1(n_4370),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.C(n_531),
.Y(n_4523)
);

AOI322xp5_ASAP7_75t_L g4524 ( 
.A1(n_4296),
.A2(n_537),
.A3(n_536),
.B1(n_534),
.B2(n_532),
.C1(n_533),
.C2(n_535),
.Y(n_4524)
);

NAND4xp25_ASAP7_75t_L g4525 ( 
.A(n_4363),
.B(n_1028),
.C(n_534),
.D(n_532),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4353),
.B(n_533),
.Y(n_4526)
);

OAI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_4313),
.A2(n_535),
.B(n_536),
.Y(n_4527)
);

AOI322xp5_ASAP7_75t_L g4528 ( 
.A1(n_4296),
.A2(n_1027),
.A3(n_543),
.B1(n_540),
.B2(n_542),
.C1(n_538),
.C2(n_539),
.Y(n_4528)
);

OAI22xp33_ASAP7_75t_L g4529 ( 
.A1(n_4293),
.A2(n_546),
.B1(n_538),
.B2(n_541),
.Y(n_4529)
);

AOI21xp5_ASAP7_75t_L g4530 ( 
.A1(n_4313),
.A2(n_541),
.B(n_546),
.Y(n_4530)
);

NOR3xp33_ASAP7_75t_L g4531 ( 
.A(n_4304),
.B(n_547),
.C(n_548),
.Y(n_4531)
);

AOI221xp5_ASAP7_75t_L g4532 ( 
.A1(n_4370),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.C(n_550),
.Y(n_4532)
);

NAND4xp25_ASAP7_75t_L g4533 ( 
.A(n_4363),
.B(n_1011),
.C(n_553),
.D(n_551),
.Y(n_4533)
);

AOI22xp5_ASAP7_75t_L g4534 ( 
.A1(n_4293),
.A2(n_554),
.B1(n_551),
.B2(n_552),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_L g4535 ( 
.A1(n_4293),
.A2(n_558),
.B1(n_552),
.B2(n_555),
.Y(n_4535)
);

NAND3xp33_ASAP7_75t_SL g4536 ( 
.A(n_4313),
.B(n_555),
.C(n_558),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4353),
.B(n_559),
.Y(n_4537)
);

AOI211xp5_ASAP7_75t_L g4538 ( 
.A1(n_4353),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_4538)
);

AOI22xp5_ASAP7_75t_L g4539 ( 
.A1(n_4293),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_4539)
);

O2A1O1Ixp33_ASAP7_75t_L g4540 ( 
.A1(n_4313),
.A2(n_564),
.B(n_562),
.C(n_563),
.Y(n_4540)
);

AOI21xp5_ASAP7_75t_L g4541 ( 
.A1(n_4313),
.A2(n_564),
.B(n_565),
.Y(n_4541)
);

OAI221xp5_ASAP7_75t_L g4542 ( 
.A1(n_4313),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.C(n_568),
.Y(n_4542)
);

AOI221xp5_ASAP7_75t_L g4543 ( 
.A1(n_4370),
.A2(n_569),
.B1(n_566),
.B2(n_568),
.C(n_570),
.Y(n_4543)
);

AOI21xp33_ASAP7_75t_SL g4544 ( 
.A1(n_4353),
.A2(n_569),
.B(n_570),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4353),
.B(n_571),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4353),
.B(n_572),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4313),
.A2(n_572),
.B(n_573),
.Y(n_4547)
);

OAI221xp5_ASAP7_75t_L g4548 ( 
.A1(n_4313),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.C(n_577),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4353),
.B(n_574),
.Y(n_4549)
);

INVx1_ASAP7_75t_SL g4550 ( 
.A(n_4294),
.Y(n_4550)
);

A2O1A1Ixp33_ASAP7_75t_L g4551 ( 
.A1(n_4313),
.A2(n_578),
.B(n_575),
.C(n_576),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4353),
.B(n_579),
.Y(n_4552)
);

OAI21xp33_ASAP7_75t_L g4553 ( 
.A1(n_4293),
.A2(n_579),
.B(n_581),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4353),
.B(n_581),
.Y(n_4554)
);

NOR2xp33_ASAP7_75t_L g4555 ( 
.A(n_4293),
.B(n_582),
.Y(n_4555)
);

O2A1O1Ixp33_ASAP7_75t_L g4556 ( 
.A1(n_4313),
.A2(n_584),
.B(n_582),
.C(n_583),
.Y(n_4556)
);

OAI22xp33_ASAP7_75t_L g4557 ( 
.A1(n_4293),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4293),
.Y(n_4558)
);

OAI211xp5_ASAP7_75t_SL g4559 ( 
.A1(n_4363),
.A2(n_588),
.B(n_585),
.C(n_586),
.Y(n_4559)
);

AOI21xp5_ASAP7_75t_L g4560 ( 
.A1(n_4313),
.A2(n_589),
.B(n_590),
.Y(n_4560)
);

OAI211xp5_ASAP7_75t_L g4561 ( 
.A1(n_4524),
.A2(n_593),
.B(n_589),
.C(n_591),
.Y(n_4561)
);

NOR3x1_ASAP7_75t_L g4562 ( 
.A(n_4542),
.B(n_591),
.C(n_593),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4455),
.Y(n_4563)
);

AOI221xp5_ASAP7_75t_SL g4564 ( 
.A1(n_4530),
.A2(n_4541),
.B1(n_4560),
.B2(n_4411),
.C(n_4422),
.Y(n_4564)
);

NAND3xp33_ASAP7_75t_L g4565 ( 
.A(n_4544),
.B(n_1009),
.C(n_596),
.Y(n_4565)
);

NOR3xp33_ASAP7_75t_L g4566 ( 
.A(n_4484),
.B(n_1009),
.C(n_596),
.Y(n_4566)
);

NAND4xp25_ASAP7_75t_L g4567 ( 
.A(n_4414),
.B(n_599),
.C(n_597),
.D(n_598),
.Y(n_4567)
);

O2A1O1Ixp5_ASAP7_75t_SL g4568 ( 
.A1(n_4488),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_4568)
);

AOI32xp33_ASAP7_75t_L g4569 ( 
.A1(n_4559),
.A2(n_604),
.A3(n_600),
.B1(n_603),
.B2(n_605),
.Y(n_4569)
);

AOI21xp33_ASAP7_75t_SL g4570 ( 
.A1(n_4491),
.A2(n_603),
.B(n_604),
.Y(n_4570)
);

OAI222xp33_ASAP7_75t_L g4571 ( 
.A1(n_4550),
.A2(n_608),
.B1(n_610),
.B2(n_605),
.C1(n_606),
.C2(n_609),
.Y(n_4571)
);

BUFx6f_ASAP7_75t_L g4572 ( 
.A(n_4558),
.Y(n_4572)
);

AOI322xp5_ASAP7_75t_L g4573 ( 
.A1(n_4536),
.A2(n_614),
.A3(n_612),
.B1(n_610),
.B2(n_606),
.C1(n_609),
.C2(n_611),
.Y(n_4573)
);

AOI22xp5_ASAP7_75t_L g4574 ( 
.A1(n_4522),
.A2(n_4531),
.B1(n_4428),
.B2(n_4468),
.Y(n_4574)
);

NAND3xp33_ASAP7_75t_L g4575 ( 
.A(n_4528),
.B(n_612),
.C(n_615),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4499),
.Y(n_4576)
);

OAI21xp5_ASAP7_75t_L g4577 ( 
.A1(n_4551),
.A2(n_4556),
.B(n_4540),
.Y(n_4577)
);

AOI321xp33_ASAP7_75t_L g4578 ( 
.A1(n_4426),
.A2(n_1008),
.A3(n_618),
.B1(n_620),
.B2(n_615),
.C(n_616),
.Y(n_4578)
);

OAI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_4548),
.A2(n_622),
.B1(n_619),
.B2(n_621),
.Y(n_4579)
);

NOR2x1_ASAP7_75t_L g4580 ( 
.A(n_4519),
.B(n_622),
.Y(n_4580)
);

NOR3xp33_ASAP7_75t_L g4581 ( 
.A(n_4415),
.B(n_1007),
.C(n_623),
.Y(n_4581)
);

OAI22xp5_ASAP7_75t_SL g4582 ( 
.A1(n_4454),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4420),
.B(n_626),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_4440),
.A2(n_627),
.B(n_629),
.Y(n_4584)
);

A2O1A1Ixp33_ASAP7_75t_L g4585 ( 
.A1(n_4469),
.A2(n_1007),
.B(n_632),
.C(n_629),
.Y(n_4585)
);

A2O1A1Ixp33_ASAP7_75t_L g4586 ( 
.A1(n_4527),
.A2(n_4547),
.B(n_4538),
.C(n_4465),
.Y(n_4586)
);

AOI221xp5_ASAP7_75t_L g4587 ( 
.A1(n_4417),
.A2(n_1005),
.B1(n_633),
.B2(n_630),
.C(n_632),
.Y(n_4587)
);

OAI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4438),
.A2(n_634),
.B(n_635),
.Y(n_4588)
);

AOI211xp5_ASAP7_75t_L g4589 ( 
.A1(n_4475),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4457),
.Y(n_4590)
);

NOR2x1_ASAP7_75t_L g4591 ( 
.A(n_4526),
.B(n_636),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_SL g4592 ( 
.A(n_4423),
.B(n_638),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_SL g4593 ( 
.A1(n_4509),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4446),
.Y(n_4594)
);

OAI22xp33_ASAP7_75t_L g4595 ( 
.A1(n_4433),
.A2(n_643),
.B1(n_639),
.B2(n_642),
.Y(n_4595)
);

OAI221xp5_ASAP7_75t_L g4596 ( 
.A1(n_4496),
.A2(n_4427),
.B1(n_4497),
.B2(n_4514),
.C(n_4412),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4537),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4512),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4545),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_SL g4600 ( 
.A(n_4487),
.B(n_642),
.Y(n_4600)
);

OAI21xp33_ASAP7_75t_L g4601 ( 
.A1(n_4413),
.A2(n_4416),
.B(n_4505),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4546),
.Y(n_4602)
);

AOI221x1_ASAP7_75t_L g4603 ( 
.A1(n_4525),
.A2(n_648),
.B1(n_644),
.B2(n_646),
.C(n_649),
.Y(n_4603)
);

AOI21xp33_ASAP7_75t_L g4604 ( 
.A1(n_4431),
.A2(n_4480),
.B(n_4511),
.Y(n_4604)
);

AOI22xp5_ASAP7_75t_L g4605 ( 
.A1(n_4482),
.A2(n_650),
.B1(n_644),
.B2(n_648),
.Y(n_4605)
);

AOI32xp33_ASAP7_75t_L g4606 ( 
.A1(n_4459),
.A2(n_4421),
.A3(n_4444),
.B1(n_4521),
.B2(n_4518),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4549),
.Y(n_4607)
);

AOI221xp5_ASAP7_75t_L g4608 ( 
.A1(n_4452),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.C(n_653),
.Y(n_4608)
);

AOI221xp5_ASAP7_75t_L g4609 ( 
.A1(n_4436),
.A2(n_4523),
.B1(n_4543),
.B2(n_4532),
.C(n_4533),
.Y(n_4609)
);

OAI21xp33_ASAP7_75t_L g4610 ( 
.A1(n_4552),
.A2(n_651),
.B(n_652),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4554),
.Y(n_4611)
);

AOI222xp33_ASAP7_75t_L g4612 ( 
.A1(n_4456),
.A2(n_655),
.B1(n_657),
.B2(n_653),
.C1(n_654),
.C2(n_656),
.Y(n_4612)
);

AOI21xp33_ASAP7_75t_L g4613 ( 
.A1(n_4443),
.A2(n_1004),
.B(n_654),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4490),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_4614)
);

AOI22xp5_ASAP7_75t_L g4615 ( 
.A1(n_4555),
.A2(n_662),
.B1(n_659),
.B2(n_661),
.Y(n_4615)
);

NOR2xp33_ASAP7_75t_L g4616 ( 
.A(n_4439),
.B(n_662),
.Y(n_4616)
);

AOI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_4508),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_4617)
);

OAI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4448),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_4618)
);

OAI221xp5_ASAP7_75t_L g4619 ( 
.A1(n_4474),
.A2(n_669),
.B1(n_667),
.B2(n_668),
.C(n_670),
.Y(n_4619)
);

AOI22xp5_ASAP7_75t_L g4620 ( 
.A1(n_4466),
.A2(n_671),
.B1(n_667),
.B2(n_669),
.Y(n_4620)
);

O2A1O1Ixp33_ASAP7_75t_SL g4621 ( 
.A1(n_4478),
.A2(n_673),
.B(n_671),
.C(n_672),
.Y(n_4621)
);

OAI21x1_ASAP7_75t_L g4622 ( 
.A1(n_4419),
.A2(n_1004),
.B(n_673),
.Y(n_4622)
);

OAI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_4464),
.A2(n_4460),
.B1(n_4498),
.B2(n_4486),
.Y(n_4623)
);

OAI321xp33_ASAP7_75t_L g4624 ( 
.A1(n_4489),
.A2(n_677),
.A3(n_679),
.B1(n_674),
.B2(n_675),
.C(n_678),
.Y(n_4624)
);

AOI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4424),
.A2(n_678),
.B(n_679),
.Y(n_4625)
);

AOI222xp33_ASAP7_75t_L g4626 ( 
.A1(n_4451),
.A2(n_682),
.B1(n_685),
.B2(n_680),
.C1(n_681),
.C2(n_684),
.Y(n_4626)
);

OAI21xp5_ASAP7_75t_L g4627 ( 
.A1(n_4504),
.A2(n_680),
.B(n_684),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4442),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4447),
.Y(n_4629)
);

NAND3xp33_ASAP7_75t_SL g4630 ( 
.A(n_4435),
.B(n_686),
.C(n_687),
.Y(n_4630)
);

OAI21xp5_ASAP7_75t_SL g4631 ( 
.A1(n_4517),
.A2(n_686),
.B(n_687),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4516),
.Y(n_4632)
);

OAI221xp5_ASAP7_75t_L g4633 ( 
.A1(n_4449),
.A2(n_691),
.B1(n_688),
.B2(n_690),
.C(n_693),
.Y(n_4633)
);

AOI22xp33_ASAP7_75t_L g4634 ( 
.A1(n_4494),
.A2(n_696),
.B1(n_693),
.B2(n_694),
.Y(n_4634)
);

A2O1A1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4472),
.A2(n_1002),
.B(n_697),
.C(n_694),
.Y(n_4635)
);

AOI211xp5_ASAP7_75t_SL g4636 ( 
.A1(n_4473),
.A2(n_701),
.B(n_696),
.C(n_699),
.Y(n_4636)
);

AOI21xp33_ASAP7_75t_SL g4637 ( 
.A1(n_4520),
.A2(n_701),
.B(n_702),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4462),
.Y(n_4638)
);

OAI21xp5_ASAP7_75t_SL g4639 ( 
.A1(n_4429),
.A2(n_702),
.B(n_703),
.Y(n_4639)
);

OAI211xp5_ASAP7_75t_L g4640 ( 
.A1(n_4501),
.A2(n_706),
.B(n_703),
.C(n_705),
.Y(n_4640)
);

A2O1A1Ixp33_ASAP7_75t_L g4641 ( 
.A1(n_4502),
.A2(n_708),
.B(n_706),
.C(n_707),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4492),
.Y(n_4642)
);

AO21x1_ASAP7_75t_L g4643 ( 
.A1(n_4445),
.A2(n_707),
.B(n_708),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4506),
.Y(n_4644)
);

OAI22xp5_ASAP7_75t_L g4645 ( 
.A1(n_4477),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4479),
.B(n_710),
.Y(n_4646)
);

INVxp67_ASAP7_75t_L g4647 ( 
.A(n_4483),
.Y(n_4647)
);

AOI322xp5_ASAP7_75t_L g4648 ( 
.A1(n_4425),
.A2(n_711),
.A3(n_712),
.B1(n_713),
.B2(n_715),
.C1(n_717),
.C2(n_719),
.Y(n_4648)
);

INVx2_ASAP7_75t_SL g4649 ( 
.A(n_4572),
.Y(n_4649)
);

OAI22xp33_ASAP7_75t_L g4650 ( 
.A1(n_4636),
.A2(n_4495),
.B1(n_4476),
.B2(n_4453),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_SL g4651 ( 
.A(n_4572),
.B(n_4507),
.Y(n_4651)
);

INVx4_ASAP7_75t_L g4652 ( 
.A(n_4572),
.Y(n_4652)
);

OAI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4565),
.A2(n_4470),
.B(n_4500),
.Y(n_4653)
);

OAI21xp5_ASAP7_75t_SL g4654 ( 
.A1(n_4574),
.A2(n_4471),
.B(n_4515),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4563),
.Y(n_4655)
);

AOI211xp5_ASAP7_75t_L g4656 ( 
.A1(n_4621),
.A2(n_4461),
.B(n_4493),
.C(n_4430),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4643),
.Y(n_4657)
);

AOI22xp5_ASAP7_75t_L g4658 ( 
.A1(n_4581),
.A2(n_4434),
.B1(n_4553),
.B2(n_4481),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4580),
.Y(n_4659)
);

OAI221xp5_ASAP7_75t_L g4660 ( 
.A1(n_4631),
.A2(n_4458),
.B1(n_4467),
.B2(n_4450),
.C(n_4535),
.Y(n_4660)
);

OA22x2_ASAP7_75t_L g4661 ( 
.A1(n_4582),
.A2(n_4539),
.B1(n_4534),
.B2(n_4513),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4590),
.B(n_4576),
.Y(n_4662)
);

AOI21xp5_ASAP7_75t_L g4663 ( 
.A1(n_4600),
.A2(n_4510),
.B(n_4529),
.Y(n_4663)
);

AOI221xp5_ASAP7_75t_L g4664 ( 
.A1(n_4596),
.A2(n_4557),
.B1(n_4437),
.B2(n_4441),
.C(n_4432),
.Y(n_4664)
);

BUFx2_ASAP7_75t_L g4665 ( 
.A(n_4591),
.Y(n_4665)
);

NOR2xp67_ASAP7_75t_L g4666 ( 
.A(n_4640),
.B(n_713),
.Y(n_4666)
);

INVx1_ASAP7_75t_SL g4667 ( 
.A(n_4583),
.Y(n_4667)
);

AOI22xp5_ASAP7_75t_L g4668 ( 
.A1(n_4647),
.A2(n_4485),
.B1(n_4463),
.B2(n_4418),
.Y(n_4668)
);

NOR3xp33_ASAP7_75t_L g4669 ( 
.A(n_4604),
.B(n_4503),
.C(n_721),
.Y(n_4669)
);

AOI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4584),
.A2(n_721),
.B(n_722),
.Y(n_4670)
);

NOR3xp33_ASAP7_75t_L g4671 ( 
.A(n_4601),
.B(n_722),
.C(n_723),
.Y(n_4671)
);

AOI221xp5_ASAP7_75t_L g4672 ( 
.A1(n_4567),
.A2(n_4570),
.B1(n_4609),
.B2(n_4575),
.C(n_4606),
.Y(n_4672)
);

OAI321xp33_ASAP7_75t_L g4673 ( 
.A1(n_4577),
.A2(n_725),
.A3(n_727),
.B1(n_723),
.B2(n_724),
.C(n_726),
.Y(n_4673)
);

AOI322xp5_ASAP7_75t_L g4674 ( 
.A1(n_4564),
.A2(n_724),
.A3(n_727),
.B1(n_729),
.B2(n_730),
.C1(n_731),
.C2(n_733),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_L g4675 ( 
.A1(n_4586),
.A2(n_4588),
.B(n_4595),
.Y(n_4675)
);

HB1xp67_ASAP7_75t_L g4676 ( 
.A(n_4622),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4573),
.B(n_729),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4646),
.Y(n_4678)
);

INVxp67_ASAP7_75t_L g4679 ( 
.A(n_4616),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4597),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4599),
.Y(n_4681)
);

OAI22xp33_ASAP7_75t_SL g4682 ( 
.A1(n_4592),
.A2(n_734),
.B1(n_731),
.B2(n_733),
.Y(n_4682)
);

AOI22xp33_ASAP7_75t_L g4683 ( 
.A1(n_4630),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.Y(n_4683)
);

XNOR2xp5_ASAP7_75t_L g4684 ( 
.A(n_4623),
.B(n_735),
.Y(n_4684)
);

OAI21xp5_ASAP7_75t_L g4685 ( 
.A1(n_4585),
.A2(n_736),
.B(n_737),
.Y(n_4685)
);

AOI22xp5_ASAP7_75t_L g4686 ( 
.A1(n_4566),
.A2(n_740),
.B1(n_737),
.B2(n_738),
.Y(n_4686)
);

AOI321xp33_ASAP7_75t_L g4687 ( 
.A1(n_4602),
.A2(n_742),
.A3(n_744),
.B1(n_738),
.B2(n_741),
.C(n_743),
.Y(n_4687)
);

NAND3xp33_ASAP7_75t_L g4688 ( 
.A(n_4589),
.B(n_744),
.C(n_745),
.Y(n_4688)
);

AOI221xp5_ASAP7_75t_L g4689 ( 
.A1(n_4624),
.A2(n_748),
.B1(n_746),
.B2(n_747),
.C(n_749),
.Y(n_4689)
);

NAND2xp33_ASAP7_75t_R g4690 ( 
.A(n_4637),
.B(n_746),
.Y(n_4690)
);

OAI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4635),
.A2(n_747),
.B(n_749),
.Y(n_4691)
);

AO21x1_ASAP7_75t_L g4692 ( 
.A1(n_4639),
.A2(n_750),
.B(n_751),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4625),
.A2(n_752),
.B(n_754),
.Y(n_4693)
);

OAI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4634),
.A2(n_756),
.B1(n_752),
.B2(n_755),
.Y(n_4694)
);

AOI22xp5_ASAP7_75t_L g4695 ( 
.A1(n_4561),
.A2(n_757),
.B1(n_755),
.B2(n_756),
.Y(n_4695)
);

AOI22xp5_ASAP7_75t_L g4696 ( 
.A1(n_4607),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_4696)
);

OAI221xp5_ASAP7_75t_L g4697 ( 
.A1(n_4569),
.A2(n_761),
.B1(n_758),
.B2(n_760),
.C(n_762),
.Y(n_4697)
);

INVx1_ASAP7_75t_SL g4698 ( 
.A(n_4593),
.Y(n_4698)
);

NAND4xp75_ASAP7_75t_L g4699 ( 
.A(n_4562),
.B(n_762),
.C(n_760),
.D(n_761),
.Y(n_4699)
);

OAI211xp5_ASAP7_75t_SL g4700 ( 
.A1(n_4611),
.A2(n_765),
.B(n_763),
.C(n_764),
.Y(n_4700)
);

AOI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4608),
.A2(n_766),
.B1(n_763),
.B2(n_765),
.Y(n_4701)
);

AOI22x1_ASAP7_75t_L g4702 ( 
.A1(n_4578),
.A2(n_770),
.B1(n_766),
.B2(n_769),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4648),
.B(n_769),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4605),
.Y(n_4704)
);

OAI21xp33_ASAP7_75t_SL g4705 ( 
.A1(n_4594),
.A2(n_771),
.B(n_772),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4610),
.Y(n_4706)
);

NAND4xp75_ASAP7_75t_L g4707 ( 
.A(n_4649),
.B(n_4638),
.C(n_4632),
.D(n_4644),
.Y(n_4707)
);

NOR2x1p5_ASAP7_75t_L g4708 ( 
.A(n_4699),
.B(n_4598),
.Y(n_4708)
);

AOI221xp5_ASAP7_75t_SL g4709 ( 
.A1(n_4650),
.A2(n_4642),
.B1(n_4633),
.B2(n_4629),
.C(n_4628),
.Y(n_4709)
);

AOI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4669),
.A2(n_4645),
.B1(n_4579),
.B2(n_4587),
.Y(n_4710)
);

AOI321xp33_ASAP7_75t_L g4711 ( 
.A1(n_4651),
.A2(n_4619),
.A3(n_4614),
.B1(n_4618),
.B2(n_4641),
.C(n_4617),
.Y(n_4711)
);

AOI22xp5_ASAP7_75t_L g4712 ( 
.A1(n_4698),
.A2(n_4612),
.B1(n_4626),
.B2(n_4620),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4666),
.B(n_4603),
.Y(n_4713)
);

A2O1A1Ixp33_ASAP7_75t_L g4714 ( 
.A1(n_4674),
.A2(n_4627),
.B(n_4613),
.C(n_4615),
.Y(n_4714)
);

AOI322xp5_ASAP7_75t_L g4715 ( 
.A1(n_4672),
.A2(n_4568),
.A3(n_4571),
.B1(n_775),
.B2(n_776),
.C1(n_778),
.C2(n_779),
.Y(n_4715)
);

AOI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_4662),
.A2(n_779),
.B1(n_772),
.B2(n_774),
.Y(n_4716)
);

OAI21xp5_ASAP7_75t_L g4717 ( 
.A1(n_4670),
.A2(n_780),
.B(n_781),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4665),
.Y(n_4718)
);

AOI211xp5_ASAP7_75t_L g4719 ( 
.A1(n_4682),
.A2(n_783),
.B(n_780),
.C(n_782),
.Y(n_4719)
);

OAI22xp33_ASAP7_75t_L g4720 ( 
.A1(n_4657),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_4720)
);

AOI22xp33_ASAP7_75t_L g4721 ( 
.A1(n_4671),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.Y(n_4721)
);

HB1xp67_ASAP7_75t_L g4722 ( 
.A(n_4659),
.Y(n_4722)
);

O2A1O1Ixp33_ASAP7_75t_L g4723 ( 
.A1(n_4676),
.A2(n_787),
.B(n_785),
.C(n_786),
.Y(n_4723)
);

OAI21xp5_ASAP7_75t_SL g4724 ( 
.A1(n_4668),
.A2(n_787),
.B(n_789),
.Y(n_4724)
);

INVx2_ASAP7_75t_SL g4725 ( 
.A(n_4652),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4652),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4655),
.B(n_789),
.Y(n_4727)
);

AOI22xp5_ASAP7_75t_L g4728 ( 
.A1(n_4654),
.A2(n_792),
.B1(n_790),
.B2(n_791),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4695),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.Y(n_4729)
);

OAI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_4705),
.A2(n_794),
.B(n_795),
.Y(n_4730)
);

OAI22xp5_ASAP7_75t_L g4731 ( 
.A1(n_4683),
.A2(n_797),
.B1(n_794),
.B2(n_796),
.Y(n_4731)
);

OAI21xp33_ASAP7_75t_L g4732 ( 
.A1(n_4658),
.A2(n_799),
.B(n_801),
.Y(n_4732)
);

O2A1O1Ixp33_ASAP7_75t_SL g4733 ( 
.A1(n_4656),
.A2(n_803),
.B(n_799),
.C(n_801),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4653),
.B(n_804),
.Y(n_4734)
);

O2A1O1Ixp33_ASAP7_75t_SL g4735 ( 
.A1(n_4677),
.A2(n_808),
.B(n_804),
.C(n_805),
.Y(n_4735)
);

OAI211xp5_ASAP7_75t_L g4736 ( 
.A1(n_4702),
.A2(n_810),
.B(n_805),
.C(n_809),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4684),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4689),
.B(n_809),
.Y(n_4738)
);

NAND3xp33_ASAP7_75t_SL g4739 ( 
.A(n_4692),
.B(n_810),
.C(n_811),
.Y(n_4739)
);

OR2x2_ASAP7_75t_L g4740 ( 
.A(n_4703),
.B(n_812),
.Y(n_4740)
);

NOR2xp33_ASAP7_75t_L g4741 ( 
.A(n_4697),
.B(n_812),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4722),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4734),
.B(n_4708),
.Y(n_4743)
);

AOI22xp5_ASAP7_75t_L g4744 ( 
.A1(n_4724),
.A2(n_4661),
.B1(n_4690),
.B2(n_4664),
.Y(n_4744)
);

AOI22xp5_ASAP7_75t_L g4745 ( 
.A1(n_4718),
.A2(n_4706),
.B1(n_4704),
.B2(n_4694),
.Y(n_4745)
);

NOR2x1_ASAP7_75t_L g4746 ( 
.A(n_4739),
.B(n_4700),
.Y(n_4746)
);

NOR2x1_ASAP7_75t_L g4747 ( 
.A(n_4720),
.B(n_4688),
.Y(n_4747)
);

BUFx2_ASAP7_75t_L g4748 ( 
.A(n_4730),
.Y(n_4748)
);

NOR2xp33_ASAP7_75t_L g4749 ( 
.A(n_4736),
.B(n_4660),
.Y(n_4749)
);

NOR2xp67_ASAP7_75t_L g4750 ( 
.A(n_4725),
.B(n_4673),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4713),
.Y(n_4751)
);

OR2x2_ASAP7_75t_L g4752 ( 
.A(n_4727),
.B(n_4667),
.Y(n_4752)
);

NOR2xp67_ASAP7_75t_L g4753 ( 
.A(n_4726),
.B(n_4663),
.Y(n_4753)
);

AOI211xp5_ASAP7_75t_L g4754 ( 
.A1(n_4733),
.A2(n_4675),
.B(n_4691),
.C(n_4685),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4717),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4715),
.B(n_4686),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4707),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4740),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4723),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4742),
.Y(n_4760)
);

AOI22xp5_ASAP7_75t_L g4761 ( 
.A1(n_4753),
.A2(n_4741),
.B1(n_4712),
.B2(n_4710),
.Y(n_4761)
);

NOR2x1_ASAP7_75t_L g4762 ( 
.A(n_4750),
.B(n_4748),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4754),
.B(n_4719),
.Y(n_4763)
);

XNOR2x1_ASAP7_75t_L g4764 ( 
.A(n_4746),
.B(n_4737),
.Y(n_4764)
);

NAND4xp75_ASAP7_75t_L g4765 ( 
.A(n_4747),
.B(n_4709),
.C(n_4680),
.D(n_4681),
.Y(n_4765)
);

AND5x1_ASAP7_75t_L g4766 ( 
.A(n_4749),
.B(n_4711),
.C(n_4714),
.D(n_4735),
.E(n_4701),
.Y(n_4766)
);

AO22x2_ASAP7_75t_L g4767 ( 
.A1(n_4759),
.A2(n_4731),
.B1(n_4678),
.B2(n_4693),
.Y(n_4767)
);

NOR2x1_ASAP7_75t_L g4768 ( 
.A(n_4743),
.B(n_4757),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4752),
.Y(n_4769)
);

NOR2x1p5_ASAP7_75t_L g4770 ( 
.A(n_4756),
.B(n_4738),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4744),
.Y(n_4771)
);

NOR3xp33_ASAP7_75t_L g4772 ( 
.A(n_4762),
.B(n_4751),
.C(n_4679),
.Y(n_4772)
);

XNOR2xp5_ASAP7_75t_L g4773 ( 
.A(n_4764),
.B(n_4745),
.Y(n_4773)
);

O2A1O1Ixp33_ASAP7_75t_L g4774 ( 
.A1(n_4771),
.A2(n_4755),
.B(n_4758),
.C(n_4732),
.Y(n_4774)
);

AND4x1_ASAP7_75t_L g4775 ( 
.A(n_4768),
.B(n_4721),
.C(n_4728),
.D(n_4716),
.Y(n_4775)
);

OAI211xp5_ASAP7_75t_SL g4776 ( 
.A1(n_4761),
.A2(n_4729),
.B(n_4687),
.C(n_4696),
.Y(n_4776)
);

AND4x1_ASAP7_75t_L g4777 ( 
.A(n_4760),
.B(n_816),
.C(n_814),
.D(n_815),
.Y(n_4777)
);

AND2x4_ASAP7_75t_L g4778 ( 
.A(n_4769),
.B(n_815),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4765),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_4779)
);

NOR3xp33_ASAP7_75t_L g4780 ( 
.A(n_4763),
.B(n_818),
.C(n_819),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_SL g4781 ( 
.A(n_4779),
.B(n_4766),
.Y(n_4781)
);

AND2x4_ASAP7_75t_L g4782 ( 
.A(n_4772),
.B(n_4770),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4778),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4778),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4783),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4784),
.B(n_4780),
.Y(n_4786)
);

OAI22xp5_ASAP7_75t_SL g4787 ( 
.A1(n_4782),
.A2(n_4773),
.B1(n_4775),
.B2(n_4777),
.Y(n_4787)
);

AO22x2_ASAP7_75t_L g4788 ( 
.A1(n_4785),
.A2(n_4781),
.B1(n_4774),
.B2(n_4776),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_SL g4789 ( 
.A1(n_4788),
.A2(n_4786),
.B(n_4767),
.Y(n_4789)
);

CKINVDCx20_ASAP7_75t_R g4790 ( 
.A(n_4789),
.Y(n_4790)
);

OAI22xp33_ASAP7_75t_L g4791 ( 
.A1(n_4790),
.A2(n_4787),
.B1(n_821),
.B2(n_819),
.Y(n_4791)
);

OAI21x1_ASAP7_75t_L g4792 ( 
.A1(n_4790),
.A2(n_820),
.B(n_822),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4791),
.B(n_822),
.Y(n_4793)
);

OAI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4792),
.A2(n_825),
.B1(n_823),
.B2(n_824),
.Y(n_4794)
);

AOI222xp33_ASAP7_75t_SL g4795 ( 
.A1(n_4794),
.A2(n_4793),
.B1(n_825),
.B2(n_826),
.C1(n_827),
.C2(n_828),
.Y(n_4795)
);

AOI222xp33_ASAP7_75t_SL g4796 ( 
.A1(n_4794),
.A2(n_996),
.B1(n_826),
.B2(n_827),
.C1(n_829),
.C2(n_830),
.Y(n_4796)
);

AOI22xp33_ASAP7_75t_L g4797 ( 
.A1(n_4795),
.A2(n_830),
.B1(n_824),
.B2(n_829),
.Y(n_4797)
);

OAI22xp33_ASAP7_75t_L g4798 ( 
.A1(n_4796),
.A2(n_833),
.B1(n_831),
.B2(n_832),
.Y(n_4798)
);

OA21x2_ASAP7_75t_L g4799 ( 
.A1(n_4797),
.A2(n_831),
.B(n_833),
.Y(n_4799)
);

AOI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_4798),
.A2(n_834),
.B(n_835),
.Y(n_4800)
);

AOI22xp5_ASAP7_75t_L g4801 ( 
.A1(n_4799),
.A2(n_4800),
.B1(n_837),
.B2(n_834),
.Y(n_4801)
);

AOI211xp5_ASAP7_75t_L g4802 ( 
.A1(n_4801),
.A2(n_839),
.B(n_836),
.C(n_838),
.Y(n_4802)
);


endmodule