module fake_netlist_6_3657_n_16 (n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_16);

input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_16;

wire n_7;
wire n_12;
wire n_15;
wire n_14;
wire n_13;
wire n_9;
wire n_11;
wire n_8;
wire n_10;

CKINVDCx5p33_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_8),
.B1(n_10),
.B2(n_7),
.Y(n_12)
);

XNOR2x1_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_0),
.Y(n_13)
);

OAI221xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_7),
.B1(n_8),
.B2(n_2),
.C(n_1),
.Y(n_14)
);

INVxp33_ASAP7_75t_SL g15 ( 
.A(n_14),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);


endmodule