module fake_jpeg_23872_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_45),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_37),
.B1(n_27),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_56),
.B1(n_66),
.B2(n_71),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_24),
.B1(n_47),
.B2(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_17),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_37),
.B1(n_28),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_78),
.B1(n_33),
.B2(n_22),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_31),
.B1(n_29),
.B2(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_7),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_22),
.C(n_31),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_31),
.B1(n_29),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_95)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_84),
.B(n_86),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_18),
.B1(n_26),
.B2(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_87),
.Y(n_143)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_89),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_69),
.C(n_62),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_60),
.Y(n_137)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_95),
.A2(n_115),
.B1(n_61),
.B2(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_39),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_117),
.B1(n_36),
.B2(n_21),
.Y(n_135)
);

BUFx6f_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_101),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_113),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_110),
.B1(n_21),
.B2(n_20),
.Y(n_144)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_23),
.B1(n_36),
.B2(n_35),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_30),
.B1(n_36),
.B2(n_18),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_68),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_48),
.B1(n_19),
.B2(n_20),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_147),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_96),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_60),
.A3(n_61),
.B1(n_39),
.B2(n_38),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_113),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_133),
.B1(n_151),
.B2(n_97),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_67),
.B1(n_61),
.B2(n_65),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_135),
.B(n_145),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_139),
.Y(n_164)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_150),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_91),
.B1(n_116),
.B2(n_87),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_80),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_80),
.B(n_10),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_92),
.A2(n_48),
.B1(n_39),
.B2(n_38),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_94),
.B(n_50),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_157),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_100),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_156),
.B(n_167),
.C(n_183),
.Y(n_194)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_159),
.Y(n_214)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_91),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_165),
.C(n_171),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_170),
.B1(n_179),
.B2(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_127),
.B1(n_136),
.B2(n_149),
.Y(n_189)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_168),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_81),
.C(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_116),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_124),
.C(n_152),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_101),
.C(n_108),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_83),
.C(n_148),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_117),
.B1(n_102),
.B2(n_116),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_99),
.B1(n_104),
.B2(n_82),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_103),
.B(n_91),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_131),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_197),
.B(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_188),
.B(n_193),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_7),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_151),
.B1(n_149),
.B2(n_106),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_206),
.B1(n_207),
.B2(n_48),
.Y(n_232)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_162),
.A2(n_112),
.B1(n_123),
.B2(n_121),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_38),
.B1(n_48),
.B2(n_89),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_121),
.B1(n_148),
.B2(n_142),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_158),
.B1(n_139),
.B2(n_163),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_160),
.C(n_165),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_50),
.B(n_38),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_216),
.B(n_1),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

OR2x4_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_50),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_230),
.C(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_178),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_237),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_233),
.B1(n_207),
.B2(n_206),
.Y(n_246)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_238),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_168),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_231),
.B(n_232),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_178),
.C(n_154),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_50),
.B(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_105),
.B1(n_50),
.B2(n_180),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_177),
.C(n_105),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_208),
.B1(n_189),
.B2(n_209),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_7),
.B(n_14),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_1),
.C(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_244),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_249),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_186),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_201),
.B1(n_187),
.B2(n_203),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_187),
.B1(n_196),
.B2(n_186),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_202),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

BUFx4f_ASAP7_75t_SL g267 ( 
.A(n_261),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_193),
.B1(n_212),
.B2(n_188),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_217),
.C(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_268),
.C(n_275),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_253),
.B1(n_261),
.B2(n_229),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_222),
.B1(n_255),
.B2(n_205),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_224),
.C(n_227),
.Y(n_268)
);

OAI31xp33_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_238),
.A3(n_227),
.B(n_223),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_250),
.B(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_239),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_242),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_212),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_246),
.A2(n_229),
.B1(n_226),
.B2(n_195),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_200),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_1),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_294),
.B1(n_267),
.B2(n_272),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_199),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_210),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_200),
.B(n_257),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_291),
.B(n_295),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_8),
.C(n_12),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_293),
.C(n_275),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_274),
.Y(n_297)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_5),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_16),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_6),
.Y(n_295)
);

AO221x1_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_267),
.B1(n_281),
.B2(n_266),
.C(n_278),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_268),
.C(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_305),
.C(n_282),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_269),
.C(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_294),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_6),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_282),
.C(n_288),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_291),
.B(n_289),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_299),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_307),
.B(n_306),
.C(n_10),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_318),
.A2(n_11),
.B(n_3),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_321),
.B(n_315),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.C(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_4),
.B1(n_11),
.B2(n_324),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_4),
.Y(n_327)
);


endmodule