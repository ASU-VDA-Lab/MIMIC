module real_aes_1751_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g91 ( .A1(n_0), .A2(n_56), .B1(n_92), .B2(n_93), .Y(n_91) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_1), .A2(n_52), .B1(n_124), .B2(n_127), .Y(n_123) );
INVx1_ASAP7_75t_L g196 ( .A(n_2), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_3), .A2(n_175), .B1(n_176), .B2(n_182), .Y(n_174) );
INVx1_ASAP7_75t_L g182 ( .A(n_3), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_4), .B(n_239), .Y(n_333) );
INVx1_ASAP7_75t_L g173 ( .A(n_5), .Y(n_173) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_6), .A2(n_19), .B1(n_92), .B2(n_96), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_7), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_8), .A2(n_27), .B1(n_165), .B2(n_167), .Y(n_164) );
INVx2_ASAP7_75t_L g212 ( .A(n_9), .Y(n_212) );
INVx1_ASAP7_75t_L g342 ( .A(n_10), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_11), .A2(n_75), .B1(n_179), .B2(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_11), .Y(n_179) );
INVx1_ASAP7_75t_L g339 ( .A(n_12), .Y(n_339) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_13), .A2(n_170), .B1(n_171), .B2(n_184), .Y(n_169) );
INVx1_ASAP7_75t_SL g184 ( .A(n_13), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_14), .B(n_227), .Y(n_325) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_15), .A2(n_177), .B1(n_178), .B2(n_181), .Y(n_176) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_15), .Y(n_181) );
AOI33xp33_ASAP7_75t_L g276 ( .A1(n_16), .A2(n_40), .A3(n_217), .B1(n_225), .B2(n_277), .B3(n_278), .Y(n_276) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_16), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_17), .A2(n_37), .B1(n_148), .B2(n_152), .Y(n_147) );
INVx1_ASAP7_75t_L g256 ( .A(n_18), .Y(n_256) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_19), .A2(n_56), .B1(n_59), .B2(n_189), .C(n_191), .Y(n_188) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_20), .A2(n_70), .B(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g240 ( .A(n_20), .B(n_70), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_21), .B(n_235), .Y(n_302) );
INVx3_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_23), .A2(n_73), .B1(n_156), .B2(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_24), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_SL g100 ( .A(n_25), .Y(n_100) );
INVx1_ASAP7_75t_L g198 ( .A(n_26), .Y(n_198) );
AND2x2_ASAP7_75t_L g233 ( .A(n_26), .B(n_196), .Y(n_233) );
AND2x2_ASAP7_75t_L g238 ( .A(n_26), .B(n_219), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_28), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_29), .A2(n_44), .B1(n_140), .B2(n_144), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_30), .B(n_235), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_31), .A2(n_210), .B1(n_239), .B2(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_32), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_33), .B(n_227), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_34), .B(n_245), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_35), .B(n_227), .Y(n_248) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_36), .A2(n_59), .B1(n_92), .B2(n_104), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_38), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g86 ( .A1(n_39), .A2(n_66), .B1(n_87), .B2(n_105), .Y(n_86) );
INVx1_ASAP7_75t_L g561 ( .A(n_40), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_41), .B(n_227), .Y(n_288) );
INVx1_ASAP7_75t_L g221 ( .A(n_42), .Y(n_221) );
INVx1_ASAP7_75t_L g229 ( .A(n_42), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_43), .A2(n_65), .B1(n_112), .B2(n_119), .Y(n_111) );
AND2x2_ASAP7_75t_L g289 ( .A(n_45), .B(n_290), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_46), .A2(n_60), .B1(n_215), .B2(n_235), .C(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_47), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g101 ( .A(n_48), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_49), .B(n_210), .Y(n_266) );
INVx1_ASAP7_75t_L g82 ( .A(n_50), .Y(n_82) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_51), .A2(n_215), .B(n_222), .Y(n_214) );
INVx1_ASAP7_75t_L g336 ( .A(n_53), .Y(n_336) );
INVx1_ASAP7_75t_L g287 ( .A(n_54), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_55), .A2(n_215), .B(n_286), .Y(n_285) );
INVxp33_ASAP7_75t_L g193 ( .A(n_56), .Y(n_193) );
INVx1_ASAP7_75t_L g219 ( .A(n_57), .Y(n_219) );
INVx1_ASAP7_75t_L g231 ( .A(n_57), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_58), .B(n_235), .Y(n_279) );
INVxp67_ASAP7_75t_L g192 ( .A(n_59), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_61), .A2(n_83), .B1(n_84), .B2(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_61), .Y(n_552) );
AND2x2_ASAP7_75t_L g306 ( .A(n_62), .B(n_209), .Y(n_306) );
INVx1_ASAP7_75t_L g337 ( .A(n_63), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_64), .A2(n_215), .B(n_304), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_67), .A2(n_215), .B(n_271), .C(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_68), .B(n_209), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_69), .A2(n_215), .B1(n_274), .B2(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g223 ( .A(n_71), .Y(n_223) );
AND2x2_ASAP7_75t_L g280 ( .A(n_72), .B(n_209), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_74), .A2(n_254), .B(n_255), .C(n_258), .Y(n_253) );
INVx1_ASAP7_75t_L g180 ( .A(n_75), .Y(n_180) );
BUFx2_ASAP7_75t_SL g190 ( .A(n_76), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_77), .B(n_227), .Y(n_226) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_185), .B1(n_199), .B2(n_539), .C(n_541), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_169), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_83), .A2(n_84), .B1(n_543), .B2(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
OR2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_138), .Y(n_84) );
NAND4xp25_ASAP7_75t_L g85 ( .A(n_86), .B(n_111), .C(n_123), .D(n_132), .Y(n_85) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_97), .Y(n_89) );
AND2x4_ASAP7_75t_L g146 ( .A(n_90), .B(n_143), .Y(n_146) );
AND2x2_ASAP7_75t_L g159 ( .A(n_90), .B(n_117), .Y(n_159) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
INVx2_ASAP7_75t_L g116 ( .A(n_91), .Y(n_116) );
AND2x2_ASAP7_75t_L g130 ( .A(n_91), .B(n_95), .Y(n_130) );
INVx1_ASAP7_75t_L g93 ( .A(n_92), .Y(n_93) );
INVx2_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
OAI22x1_ASAP7_75t_L g98 ( .A1(n_92), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_92), .Y(n_99) );
INVx1_ASAP7_75t_L g104 ( .A(n_92), .Y(n_104) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_94), .Y(n_110) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x4_ASAP7_75t_L g115 ( .A(n_95), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
AND2x2_ASAP7_75t_L g126 ( .A(n_97), .B(n_115), .Y(n_126) );
AND2x4_ASAP7_75t_L g166 ( .A(n_97), .B(n_136), .Y(n_166) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_102), .Y(n_97) );
AND2x2_ASAP7_75t_L g108 ( .A(n_98), .B(n_103), .Y(n_108) );
INVx2_ASAP7_75t_L g118 ( .A(n_98), .Y(n_118) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
AND2x4_ASAP7_75t_L g143 ( .A(n_102), .B(n_118), .Y(n_143) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g117 ( .A(n_103), .B(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g163 ( .A(n_103), .Y(n_163) );
BUFx6f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x4_ASAP7_75t_L g121 ( .A(n_108), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g135 ( .A(n_108), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND2x4_ASAP7_75t_L g154 ( .A(n_115), .B(n_143), .Y(n_154) );
INVxp67_ASAP7_75t_L g122 ( .A(n_116), .Y(n_122) );
AND2x4_ASAP7_75t_L g136 ( .A(n_116), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g151 ( .A(n_117), .B(n_136), .Y(n_151) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx6_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx12f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x4_ASAP7_75t_L g162 ( .A(n_130), .B(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g168 ( .A(n_130), .B(n_143), .Y(n_168) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx6_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g142 ( .A(n_136), .B(n_143), .Y(n_142) );
NAND4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_147), .C(n_155), .D(n_164), .Y(n_138) );
INVx3_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx8_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx8_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx5_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_174), .B2(n_183), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_173), .A2(n_224), .B(n_232), .C(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_174), .Y(n_183) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g304 ( .A1(n_184), .A2(n_224), .B(n_232), .C(n_305), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
AND3x1_ASAP7_75t_SL g187 ( .A(n_188), .B(n_194), .C(n_197), .Y(n_187) );
INVxp67_ASAP7_75t_L g550 ( .A(n_188), .Y(n_550) );
CKINVDCx8_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_194), .Y(n_548) );
AO21x1_ASAP7_75t_SL g558 ( .A1(n_194), .A2(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g236 ( .A(n_195), .B(n_225), .Y(n_236) );
OR2x2_ASAP7_75t_SL g555 ( .A(n_195), .B(n_197), .Y(n_555) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g220 ( .A(n_196), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_197), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g216 ( .A(n_198), .B(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND3x1_ASAP7_75t_L g201 ( .A(n_202), .B(n_429), .C(n_494), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_383), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_328), .B(n_356), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_292), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_241), .Y(n_205) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_206), .A2(n_431), .B(n_442), .Y(n_430) );
AND2x2_ASAP7_75t_SL g465 ( .A(n_206), .B(n_372), .Y(n_465) );
AND2x2_ASAP7_75t_L g480 ( .A(n_206), .B(n_481), .Y(n_480) );
OR2x6_ASAP7_75t_L g490 ( .A(n_206), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g492 ( .A(n_206), .B(n_482), .Y(n_492) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g366 ( .A(n_207), .Y(n_366) );
AND2x2_ASAP7_75t_L g379 ( .A(n_207), .B(n_380), .Y(n_379) );
INVx4_ASAP7_75t_L g398 ( .A(n_207), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_207), .B(n_317), .Y(n_401) );
NOR2x1_ASAP7_75t_SL g404 ( .A(n_207), .B(n_332), .Y(n_404) );
AND2x4_ASAP7_75t_L g416 ( .A(n_207), .B(n_414), .Y(n_416) );
OR2x2_ASAP7_75t_L g426 ( .A(n_207), .B(n_299), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_207), .B(n_438), .Y(n_443) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_213), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_209), .A2(n_253), .B1(n_259), .B2(n_260), .Y(n_252) );
INVx3_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_210), .B(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
BUFx4f_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
AND2x4_ASAP7_75t_L g239 ( .A(n_212), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_212), .B(n_240), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_234), .B(n_239), .Y(n_213) );
INVxp67_ASAP7_75t_L g265 ( .A(n_215), .Y(n_265) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_216), .Y(n_559) );
INVx1_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x6_ASAP7_75t_L g224 ( .A(n_218), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x6_ASAP7_75t_L g341 ( .A(n_219), .B(n_228), .Y(n_341) );
INVx2_ASAP7_75t_L g225 ( .A(n_221), .Y(n_225) );
AND2x4_ASAP7_75t_L g344 ( .A(n_221), .B(n_230), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_226), .C(n_232), .Y(n_222) );
INVxp67_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_224), .A2(n_232), .B(n_287), .C(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g327 ( .A(n_224), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_224), .A2(n_257), .B1(n_336), .B2(n_337), .Y(n_335) );
INVxp33_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_225), .Y(n_560) );
INVx1_ASAP7_75t_L g257 ( .A(n_227), .Y(n_257) );
AND2x4_ASAP7_75t_L g540 ( .A(n_227), .B(n_233), .Y(n_540) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g274 ( .A(n_232), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_232), .A2(n_325), .B(n_326), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_232), .B(n_239), .Y(n_345) );
INVx5_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
INVx1_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g320 ( .A(n_236), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_237), .Y(n_321) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_241), .A2(n_372), .B1(n_467), .B2(n_468), .Y(n_466) );
INVx1_ASAP7_75t_SL g510 ( .A(n_241), .Y(n_510) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_268), .Y(n_241) );
INVx2_ASAP7_75t_L g441 ( .A(n_242), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_242), .B(n_387), .Y(n_513) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_250), .Y(n_242) );
BUFx3_ASAP7_75t_L g359 ( .A(n_243), .Y(n_359) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g352 ( .A(n_244), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_244), .B(n_270), .Y(n_374) );
AND2x4_ASAP7_75t_L g391 ( .A(n_244), .B(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g407 ( .A(n_244), .Y(n_407) );
INVx2_ASAP7_75t_L g464 ( .A(n_244), .Y(n_464) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_249), .Y(n_244) );
INVx2_ASAP7_75t_SL g271 ( .A(n_245), .Y(n_271) );
AND2x2_ASAP7_75t_L g382 ( .A(n_250), .B(n_348), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g428 ( .A(n_250), .B(n_351), .Y(n_428) );
AND2x2_ASAP7_75t_L g447 ( .A(n_250), .B(n_351), .Y(n_447) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g309 ( .A(n_251), .Y(n_309) );
INVx1_ASAP7_75t_L g390 ( .A(n_251), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_251), .B(n_282), .Y(n_409) );
AND2x4_ASAP7_75t_L g463 ( .A(n_251), .B(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_261), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_260), .A2(n_283), .B(n_289), .Y(n_282) );
AO21x2_ASAP7_75t_L g351 ( .A1(n_260), .A2(n_283), .B(n_289), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B1(n_266), .B2(n_267), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g422 ( .A(n_268), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_268), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_281), .Y(n_268) );
AND2x2_ASAP7_75t_L g406 ( .A(n_269), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g446 ( .A(n_269), .Y(n_446) );
AND2x2_ASAP7_75t_L g451 ( .A(n_269), .B(n_351), .Y(n_451) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_270), .B(n_282), .Y(n_311) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_280), .Y(n_270) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_271), .A2(n_272), .B(n_280), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_279), .Y(n_272) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g387 ( .A(n_281), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_281), .B(n_359), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_281), .B(n_309), .Y(n_526) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_282), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_290), .Y(n_300) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_307), .B(n_312), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_295), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g364 ( .A(n_296), .Y(n_364) );
AND2x2_ASAP7_75t_L g378 ( .A(n_296), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g412 ( .A(n_296), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g478 ( .A(n_296), .B(n_396), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_296), .B(n_525), .C(n_526), .Y(n_524) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g371 ( .A(n_299), .Y(n_371) );
AND2x2_ASAP7_75t_L g377 ( .A(n_299), .B(n_332), .Y(n_377) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_299), .Y(n_388) );
AND2x2_ASAP7_75t_L g433 ( .A(n_299), .B(n_331), .Y(n_433) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_299), .Y(n_456) );
INVx1_ASAP7_75t_L g473 ( .A(n_299), .Y(n_473) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_306), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g515 ( .A(n_307), .Y(n_515) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_308), .B(n_386), .Y(n_487) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g349 ( .A(n_309), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI211x1_ASAP7_75t_L g383 ( .A1(n_313), .A2(n_384), .B(n_393), .C(n_410), .Y(n_383) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_314), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g436 ( .A(n_314), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g372 ( .A(n_316), .B(n_331), .Y(n_372) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g330 ( .A(n_317), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_317), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_317), .Y(n_414) );
AND2x2_ASAP7_75t_L g482 ( .A(n_317), .B(n_332), .Y(n_482) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_323), .Y(n_317) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .C(n_322), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_346), .B(n_353), .Y(n_328) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_329), .B(n_398), .Y(n_501) );
INVx2_ASAP7_75t_L g533 ( .A(n_329), .Y(n_533) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g365 ( .A(n_330), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g438 ( .A(n_331), .Y(n_438) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .B(n_345), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_342), .B2(n_343), .Y(n_338) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
OR2x2_ASAP7_75t_L g440 ( .A(n_347), .B(n_441), .Y(n_440) );
NAND2x1_ASAP7_75t_SL g462 ( .A(n_347), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g362 ( .A(n_348), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
INVx1_ASAP7_75t_L g516 ( .A(n_349), .Y(n_516) );
AND2x2_ASAP7_75t_L g381 ( .A(n_350), .B(n_382), .Y(n_381) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g363 ( .A(n_351), .Y(n_363) );
INVxp33_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g420 ( .A(n_355), .B(n_413), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_367), .C(n_375), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g444 ( .A(n_358), .B(n_445), .Y(n_444) );
NOR2xp67_ASAP7_75t_SL g449 ( .A(n_358), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_359), .B(n_446), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_365), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
AND2x2_ASAP7_75t_L g493 ( .A(n_362), .B(n_463), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g511 ( .A1(n_365), .A2(n_512), .B1(n_514), .B2(n_517), .C1(n_518), .C2(n_521), .Y(n_511) );
INVx1_ASAP7_75t_L g475 ( .A(n_366), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_373), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_371), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g491 ( .A(n_372), .Y(n_491) );
AND2x2_ASAP7_75t_L g536 ( .A(n_372), .B(n_388), .Y(n_536) );
AND2x2_ASAP7_75t_L g417 ( .A(n_373), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g530 ( .A(n_374), .B(n_409), .Y(n_530) );
OAI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_378), .B(n_381), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_376), .A2(n_396), .B(n_437), .Y(n_497) );
AND2x2_ASAP7_75t_L g521 ( .A(n_377), .B(n_398), .Y(n_521) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_377), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g469 ( .A(n_380), .Y(n_469) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_380), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g504 ( .A(n_382), .Y(n_504) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AND2x2_ASAP7_75t_L g507 ( .A(n_387), .B(n_391), .Y(n_507) );
BUFx2_ASAP7_75t_L g395 ( .A(n_388), .Y(n_395) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g418 ( .A(n_390), .Y(n_418) );
INVx2_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
AND2x2_ASAP7_75t_L g460 ( .A(n_390), .B(n_451), .Y(n_460) );
AND2x4_ASAP7_75t_L g427 ( .A(n_391), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g467 ( .A(n_391), .B(n_424), .Y(n_467) );
AND2x2_ASAP7_75t_L g518 ( .A(n_391), .B(n_519), .Y(n_518) );
AOI31xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .A3(n_403), .B(n_405), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g415 ( .A(n_395), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x4_ASAP7_75t_L g413 ( .A(n_398), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_401), .A2(n_453), .B1(n_484), .B2(n_487), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_401), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g538 ( .A(n_401), .B(n_454), .Y(n_538) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_454), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
AND2x2_ASAP7_75t_L g476 ( .A(n_406), .B(n_447), .Y(n_476) );
INVx1_ASAP7_75t_L g486 ( .A(n_408), .Y(n_486) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_419), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g509 ( .A(n_412), .Y(n_509) );
AND2x2_ASAP7_75t_L g517 ( .A(n_413), .B(n_469), .Y(n_517) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_413), .Y(n_523) );
AND2x2_ASAP7_75t_L g468 ( .A(n_416), .B(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B1(n_425), .B2(n_427), .Y(n_419) );
NOR2xp33_ASAP7_75t_SL g421 ( .A(n_422), .B(n_423), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_422), .A2(n_441), .B1(n_535), .B2(n_537), .Y(n_534) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g434 ( .A(n_427), .Y(n_434) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_457), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_433), .A2(n_436), .B(n_439), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_436), .A2(n_460), .B1(n_461), .B2(n_465), .Y(n_459) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_448), .B2(n_452), .Y(n_442) );
INVx1_ASAP7_75t_L g477 ( .A(n_445), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_458), .B(n_470), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_462), .B(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g485 ( .A(n_463), .Y(n_485) );
INVx3_ASAP7_75t_L g499 ( .A(n_467), .Y(n_499) );
INVxp67_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_479), .C(n_483), .D(n_488), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x2_ASAP7_75t_L g481 ( .A(n_473), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
NAND2xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_486), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_493), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND3x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_511), .C(n_522), .Y(n_494) );
AOI221x1_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_498), .B1(n_500), .B2(n_502), .C(n_508), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g502 ( .A(n_503), .B(n_506), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
NAND2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_527), .C(n_534), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_527) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI222xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B1(n_551), .B2(n_553), .C1(n_556), .C2(n_561), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_543), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
endmodule