module fake_jpeg_17627_n_346 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_32),
.B1(n_22),
.B2(n_36),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_58),
.B1(n_63),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_32),
.B1(n_36),
.B2(n_33),
.Y(n_58)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_20),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_68),
.B1(n_46),
.B2(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_23),
.B1(n_35),
.B2(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_23),
.B1(n_20),
.B2(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_74),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_45),
.Y(n_83)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_87),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_98),
.B1(n_77),
.B2(n_50),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_46),
.B1(n_50),
.B2(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_107),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_48),
.Y(n_98)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_48),
.B(n_56),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_37),
.C(n_18),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_75),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_37),
.C(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_43),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_134),
.B1(n_90),
.B2(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_123),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_130),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_75),
.B1(n_55),
.B2(n_29),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_98),
.B1(n_86),
.B2(n_89),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_58),
.B1(n_67),
.B2(n_41),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_87),
.B1(n_91),
.B2(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_41),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_66),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_143),
.B(n_28),
.CI(n_26),
.CON(n_187),
.SN(n_187)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_64),
.B1(n_90),
.B2(n_82),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_126),
.B(n_112),
.Y(n_174)
);

AO21x1_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_99),
.B(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_107),
.B1(n_99),
.B2(n_66),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_81),
.B1(n_97),
.B2(n_94),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_156),
.B1(n_158),
.B2(n_125),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_95),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_160),
.C(n_130),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_92),
.B1(n_82),
.B2(n_102),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_37),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_124),
.C(n_110),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_28),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_114),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_182),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_131),
.A3(n_135),
.B1(n_111),
.B2(n_109),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_162),
.B(n_153),
.C(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_175),
.B(n_181),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_187),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_174),
.B1(n_184),
.B2(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_135),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_162),
.C(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_120),
.Y(n_210)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.C(n_198),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_145),
.B(n_162),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_194),
.A2(n_202),
.B1(n_204),
.B2(n_208),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_140),
.B(n_145),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_200),
.Y(n_241)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_73),
.B1(n_72),
.B2(n_60),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_150),
.B1(n_117),
.B2(n_139),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_117),
.B1(n_137),
.B2(n_122),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_216),
.B1(n_178),
.B2(n_167),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_118),
.B1(n_121),
.B2(n_120),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_159),
.B(n_121),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_115),
.B1(n_64),
.B2(n_21),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_28),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_176),
.B1(n_177),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_186),
.C(n_187),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_220),
.C(n_223),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_187),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_170),
.B1(n_189),
.B2(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_239),
.B1(n_199),
.B2(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_168),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_228),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_182),
.C(n_118),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_237),
.C(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_113),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_18),
.B(n_115),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_236),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_201),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_235),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_19),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_234),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_194),
.B(n_26),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_27),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_19),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_19),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_195),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_208),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_209),
.C(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_263),
.C(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_201),
.B1(n_217),
.B2(n_227),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_255),
.B(n_247),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_201),
.C(n_205),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_201),
.B1(n_191),
.B2(n_234),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_274),
.B1(n_3),
.B2(n_4),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_265),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_220),
.A3(n_237),
.B1(n_191),
.B2(n_26),
.C1(n_31),
.C2(n_60),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_248),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.C(n_273),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_31),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_11),
.B(n_17),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_31),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_24),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_4),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_251),
.C(n_254),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_262),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_243),
.B(n_252),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_4),
.B(n_5),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_259),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_290),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_31),
.C(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_254),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_3),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_3),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_21),
.B(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_73),
.C(n_72),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_277),
.C(n_60),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_277),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_269),
.B1(n_278),
.B2(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_292),
.B1(n_297),
.B2(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_282),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_308),
.C(n_312),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_5),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_284),
.B1(n_6),
.B2(n_7),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_308),
.B1(n_10),
.B2(n_12),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_6),
.Y(n_316)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_7),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_14),
.C(n_15),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_8),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_310),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_9),
.Y(n_329)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_303),
.B(n_312),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_330),
.B(n_15),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_324),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_10),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_317),
.C(n_320),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_335),
.A2(n_337),
.B(n_338),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_313),
.C(n_323),
.Y(n_338)
);

NAND4xp25_ASAP7_75t_SL g342 ( 
.A(n_339),
.B(n_333),
.C(n_332),
.D(n_329),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_318),
.B(n_320),
.Y(n_341)
);

AOI211xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_342),
.B(n_334),
.C(n_16),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_340),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_15),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_17),
.Y(n_346)
);


endmodule