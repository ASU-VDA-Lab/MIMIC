module fake_jpeg_31473_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g167 ( 
.A(n_53),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_89),
.Y(n_126)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_9),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_86),
.Y(n_117)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_9),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_94),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_20),
.B(n_10),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_10),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_99),
.Y(n_119)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_35),
.Y(n_129)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_107),
.A2(n_111),
.B1(n_120),
.B2(n_127),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_23),
.B1(n_44),
.B2(n_49),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_132),
.B1(n_154),
.B2(n_0),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_35),
.B1(n_19),
.B2(n_38),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_27),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_142),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_59),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_102),
.B1(n_96),
.B2(n_78),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_93),
.A2(n_35),
.B1(n_19),
.B2(n_38),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_138),
.A2(n_141),
.B1(n_33),
.B2(n_32),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_63),
.A2(n_35),
.B1(n_19),
.B2(n_38),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_54),
.B(n_46),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_83),
.C(n_104),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_149),
.C(n_45),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_46),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_27),
.C(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_54),
.B(n_49),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_53),
.B(n_51),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_151),
.B(n_164),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_69),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_33),
.B1(n_32),
.B2(n_87),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_50),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_88),
.B1(n_80),
.B2(n_65),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_169),
.A2(n_182),
.B1(n_224),
.B2(n_225),
.Y(n_241)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_124),
.A3(n_122),
.B1(n_108),
.B2(n_117),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_170),
.A2(n_172),
.B(n_135),
.C(n_159),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_48),
.B(n_47),
.C(n_45),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_47),
.B(n_33),
.C(n_45),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_173),
.B(n_184),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_47),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_201),
.Y(n_231)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_167),
.Y(n_180)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_57),
.Y(n_184)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_188),
.A2(n_216),
.B1(n_230),
.B2(n_109),
.Y(n_274)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_189),
.Y(n_247)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_84),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_221),
.B(n_186),
.Y(n_253)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_32),
.B1(n_87),
.B2(n_2),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_7),
.B1(n_17),
.B2(n_2),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_205),
.B1(n_162),
.B2(n_159),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_197),
.B(n_206),
.Y(n_273)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_7),
.B1(n_17),
.B2(n_2),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_199),
.A2(n_204),
.B1(n_210),
.B2(n_5),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_11),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_11),
.B1(n_17),
.B2(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_119),
.B(n_11),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_134),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_219),
.Y(n_235)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_18),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_217),
.Y(n_248)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_218),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_222),
.Y(n_236)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_121),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_111),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_226),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_134),
.A2(n_6),
.B1(n_16),
.B2(n_3),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_120),
.A2(n_6),
.B1(n_16),
.B2(n_3),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_135),
.Y(n_226)
);

BUFx6f_ASAP7_75t_SL g227 ( 
.A(n_106),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_105),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_0),
.Y(n_280)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_156),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_156),
.A2(n_115),
.B1(n_133),
.B2(n_160),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_234),
.B(n_263),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_254),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_130),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_260),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_184),
.B1(n_225),
.B2(n_169),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_174),
.B(n_131),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_230),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_253),
.B(n_180),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_115),
.B1(n_131),
.B2(n_155),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_179),
.B(n_130),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_106),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_269),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_268),
.Y(n_284)
);

AOI32xp33_ASAP7_75t_L g268 ( 
.A1(n_211),
.A2(n_109),
.A3(n_135),
.B1(n_116),
.B2(n_143),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_173),
.B(n_166),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_176),
.B(n_166),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_282),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_274),
.B(n_278),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_192),
.A2(n_116),
.B1(n_14),
.B2(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_205),
.B1(n_195),
.B2(n_171),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_184),
.B(n_0),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_316),
.B1(n_317),
.B2(n_278),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_231),
.B(n_172),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_306),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_187),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_309),
.Y(n_347)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_244),
.A2(n_212),
.B(n_216),
.C(n_182),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_292),
.A2(n_232),
.B(n_249),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_259),
.C(n_249),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_294),
.A2(n_296),
.B1(n_300),
.B2(n_261),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_216),
.B1(n_191),
.B2(n_177),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_175),
.C(n_181),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_299),
.C(n_325),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_242),
.B(n_229),
.C(n_207),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_242),
.A2(n_216),
.B1(n_206),
.B2(n_194),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_252),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_197),
.C(n_214),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_220),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_314),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_180),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_310),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_274),
.A2(n_193),
.B1(n_200),
.B2(n_227),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_311),
.A2(n_247),
.B(n_233),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_236),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_315),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_263),
.B(n_209),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_276),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_241),
.A2(n_202),
.B1(n_218),
.B2(n_217),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_241),
.A2(n_202),
.B1(n_213),
.B2(n_178),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_234),
.B(n_222),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_320),
.B(n_279),
.Y(n_345)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_322),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_203),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_324),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_248),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_242),
.B(n_208),
.C(n_190),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_329),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_252),
.B(n_189),
.C(n_228),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_254),
.C(n_266),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_270),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_330),
.A2(n_359),
.B(n_314),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_331),
.A2(n_335),
.B1(n_337),
.B2(n_341),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_333),
.A2(n_360),
.B1(n_365),
.B2(n_298),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_291),
.A2(n_274),
.B(n_282),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_272),
.B1(n_274),
.B2(n_260),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_339),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_275),
.B1(n_266),
.B2(n_247),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_344),
.A2(n_302),
.B(n_312),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_345),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_306),
.B(n_251),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_369),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_285),
.B(n_198),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_351),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_251),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_286),
.C(n_329),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_313),
.B(n_264),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_303),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_320),
.A2(n_279),
.B(n_259),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_292),
.B1(n_283),
.B2(n_317),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g361 ( 
.A(n_291),
.B(n_312),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_289),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_265),
.B1(n_232),
.B2(n_243),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_366),
.B1(n_297),
.B2(n_315),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_292),
.A2(n_265),
.B1(n_243),
.B2(n_237),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_300),
.A2(n_237),
.B1(n_258),
.B2(n_267),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_369),
.Y(n_371)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_364),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_372),
.B(n_379),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_307),
.B1(n_296),
.B2(n_284),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_374),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_347),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_356),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_378),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_364),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_381),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_382),
.A2(n_393),
.B(n_339),
.Y(n_407)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_301),
.B1(n_312),
.B2(n_321),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_365),
.A2(n_289),
.B1(n_308),
.B2(n_328),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_390),
.B(n_395),
.Y(n_417)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_391),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_333),
.A2(n_325),
.B1(n_295),
.B2(n_299),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_345),
.A2(n_316),
.B1(n_286),
.B2(n_326),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_398),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_288),
.B1(n_290),
.B2(n_305),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_399),
.A2(n_350),
.B1(n_354),
.B2(n_353),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_362),
.A2(n_319),
.B1(n_318),
.B2(n_323),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_267),
.B1(n_258),
.B2(n_240),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_402),
.A2(n_367),
.B1(n_346),
.B2(n_370),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_353),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_403),
.Y(n_426)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_405),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_337),
.A2(n_255),
.B1(n_310),
.B2(n_245),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_407),
.A2(n_393),
.B(n_382),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_336),
.C(n_392),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_410),
.C(n_420),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_336),
.C(n_332),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_435),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_338),
.C(n_349),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_374),
.C(n_390),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_427),
.C(n_433),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_424),
.A2(n_430),
.B1(n_432),
.B2(n_396),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_342),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_342),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_431),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_350),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_399),
.A2(n_331),
.B1(n_361),
.B2(n_359),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_354),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_348),
.C(n_330),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_366),
.C(n_400),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_343),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_384),
.C(n_382),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_438),
.B(n_461),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_439),
.A2(n_464),
.B1(n_423),
.B2(n_411),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_406),
.B(n_381),
.Y(n_442)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_426),
.Y(n_443)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_444),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_403),
.Y(n_447)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_415),
.B(n_371),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_449),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_379),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_453),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_438),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_434),
.A2(n_384),
.B(n_373),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_SL g469 ( 
.A1(n_452),
.A2(n_422),
.B(n_429),
.C(n_409),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_432),
.A2(n_405),
.B(n_363),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_418),
.Y(n_454)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_413),
.A2(n_358),
.B(n_373),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_409),
.Y(n_471)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_458),
.B1(n_459),
.B2(n_462),
.Y(n_478)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_383),
.B1(n_380),
.B2(n_394),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_460),
.A2(n_459),
.B1(n_424),
.B2(n_464),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_437),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_398),
.C(n_391),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_420),
.C(n_417),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_437),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_469),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_453),
.A2(n_433),
.B1(n_431),
.B2(n_427),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_466),
.A2(n_481),
.B1(n_439),
.B2(n_448),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_486),
.C(n_445),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_477),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_417),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_480),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_475),
.A2(n_476),
.B1(n_462),
.B2(n_449),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_460),
.A2(n_414),
.B1(n_413),
.B2(n_412),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_410),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_480),
.B(n_482),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_412),
.B1(n_386),
.B2(n_404),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_438),
.B(n_343),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_423),
.C(n_401),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_467),
.Y(n_489)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_489),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_443),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_491),
.A2(n_355),
.B(n_352),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_445),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_495),
.C(n_496),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_445),
.C(n_461),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_452),
.C(n_446),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_497),
.A2(n_500),
.B1(n_502),
.B2(n_450),
.Y(n_511)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_499),
.Y(n_512)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_483),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_485),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_446),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_504),
.C(n_476),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_465),
.C(n_482),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_442),
.B(n_451),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_5),
.B(n_12),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_493),
.A2(n_478),
.B1(n_469),
.B2(n_484),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_509),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_494),
.Y(n_525)
);

OAI321xp33_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_447),
.A3(n_472),
.B1(n_455),
.B2(n_441),
.C(n_475),
.Y(n_513)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_513),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_502),
.A2(n_469),
.B1(n_441),
.B2(n_456),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_515),
.B1(n_503),
.B2(n_367),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_493),
.A2(n_469),
.B1(n_458),
.B2(n_454),
.Y(n_515)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_495),
.A2(n_440),
.B1(n_421),
.B2(n_355),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_519),
.B1(n_501),
.B2(n_487),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_496),
.A2(n_490),
.B1(n_440),
.B2(n_503),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_507),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_508),
.Y(n_523)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_523),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_525),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_370),
.C(n_255),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_529),
.C(n_509),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_343),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_528),
.B(n_530),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_1),
.C(n_5),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_505),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_531),
.A2(n_514),
.B(n_527),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_533),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_529),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_537),
.B(n_520),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_540),
.C(n_541),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_534),
.B(n_510),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_520),
.C(n_535),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_543),
.B(n_533),
.Y(n_545)
);

AOI321xp33_ASAP7_75t_SL g544 ( 
.A1(n_542),
.A2(n_523),
.A3(n_512),
.B1(n_532),
.B2(n_519),
.C(n_517),
.Y(n_544)
);

OAI311xp33_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_545),
.A3(n_515),
.B1(n_522),
.C1(n_536),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_546),
.A2(n_530),
.B(n_518),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_512),
.C(n_511),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_12),
.C(n_15),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_18),
.B(n_16),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g551 ( 
.A(n_550),
.B(n_18),
.CI(n_1),
.CON(n_551),
.SN(n_551)
);


endmodule