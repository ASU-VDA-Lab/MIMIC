module fake_jpeg_2685_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_79),
.Y(n_89)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_73),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_62),
.B1(n_61),
.B2(n_53),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_91),
.B1(n_92),
.B2(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_61),
.B1(n_55),
.B2(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_73),
.B1(n_55),
.B2(n_65),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_109),
.Y(n_142)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_119),
.Y(n_126)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_78),
.B(n_80),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_110),
.B(n_56),
.C(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_111),
.Y(n_137)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_74),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_79),
.B(n_68),
.C(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_67),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_83),
.B(n_88),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_56),
.C(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_77),
.B1(n_69),
.B2(n_70),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_2),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_118),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_80),
.B1(n_78),
.B2(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_90),
.B1(n_58),
.B2(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_66),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_25),
.B(n_38),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_58),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_0),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_71),
.C(n_48),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_138),
.C(n_4),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_24),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_47),
.C(n_46),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_4),
.C(n_5),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_117),
.B(n_115),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_42),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_16),
.C(n_19),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_154),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_158),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_9),
.B(n_10),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_10),
.B(n_11),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_162),
.A2(n_167),
.B1(n_142),
.B2(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_14),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_15),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_181),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_19),
.B1(n_20),
.B2(n_28),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_178),
.B(n_185),
.Y(n_193)
);

NAND2x1p5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_32),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_33),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_154),
.B1(n_160),
.B2(n_166),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_157),
.B(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_175),
.B1(n_170),
.B2(n_182),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_150),
.C(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_35),
.C(n_41),
.Y(n_194)
);

HAxp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_171),
.CON(n_195),
.SN(n_195)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_172),
.B(n_180),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_174),
.B1(n_145),
.B2(n_169),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_178),
.B(n_188),
.C(n_183),
.D(n_193),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_177),
.B1(n_202),
.B2(n_205),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_201),
.C(n_198),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_196),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_210),
.A2(n_195),
.B(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_194),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_173),
.Y(n_214)
);


endmodule