module real_jpeg_23355_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_56),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_71),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_4),
.A2(n_35),
.B1(n_58),
.B2(n_168),
.Y(n_350)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_6),
.B(n_62),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_6),
.A2(n_66),
.B(n_80),
.C(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_6),
.A2(n_63),
.B1(n_66),
.B2(n_169),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_6),
.B(n_28),
.C(n_44),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_169),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_25),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_123),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_60),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_63),
.B1(n_66),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_8),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_159),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_159),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_159),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_49),
.B1(n_63),
.B2(n_66),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_9),
.A2(n_49),
.B1(n_56),
.B2(n_59),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_63),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_59),
.B1(n_84),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_59),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_63),
.B1(n_66),
.B2(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_107),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_107),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_39),
.B1(n_63),
.B2(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_39),
.B1(n_72),
.B2(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_16),
.A2(n_26),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_16),
.Y(n_191)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_16),
.A2(n_26),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_346),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_333),
.B(n_345),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_134),
.A3(n_148),
.B(n_330),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_21),
.B(n_112),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_24),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_25),
.A2(n_176),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_25),
.A2(n_96),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_25),
.A2(n_259),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_26),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_28),
.B1(n_44),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_27),
.B(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_41),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_40),
.B(n_251),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_41),
.A2(n_81),
.B(n_169),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_42),
.A2(n_50),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_42),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_42),
.A2(n_50),
.B1(n_226),
.B2(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_47),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_87),
.B1(n_101),
.B2(n_163),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_47),
.B(n_169),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_47),
.A2(n_164),
.B(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_50),
.B(n_165),
.Y(n_227)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_68),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_61),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_58),
.B1(n_65),
.B2(n_67),
.Y(n_74)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_58),
.Y(n_181)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_109),
.B1(n_131),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_61),
.A2(n_68),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_62),
.A2(n_73),
.B1(n_106),
.B2(n_200),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_62),
.A2(n_73),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_62),
.A2(n_73),
.B1(n_341),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_66),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_63),
.A2(n_67),
.B(n_170),
.C(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_SL g180 ( 
.A(n_65),
.B(n_66),
.C(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_72),
.B(n_169),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_73),
.A2(n_111),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_78),
.A2(n_79),
.B1(n_125),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_78),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_78),
.A2(n_197),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_79),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_79),
.A2(n_103),
.B(n_185),
.Y(n_309)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_87),
.A2(n_225),
.B(n_227),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_87),
.A2(n_227),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_91),
.A2(n_92),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_104),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_93),
.A2(n_94),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_95),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_97),
.B(n_169),
.Y(n_263)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_97),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_97),
.A2(n_233),
.B(n_257),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_102),
.B(n_104),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.C(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_133),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_123),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_122),
.A2(n_123),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_123),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_127),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_127),
.B(n_141),
.C(n_145),
.Y(n_344)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_130),
.B(n_137),
.C(n_140),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_135),
.A2(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_147),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_136),
.B(n_147),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_142),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_146),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_323),
.B(n_329),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_313),
.B(n_322),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_212),
.B(n_296),
.C(n_312),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_192),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_152),
.B(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_171),
.C(n_182),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_153),
.A2(n_154),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_166),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_161),
.C(n_166),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_171),
.A2(n_172),
.B1(n_182),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_182),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_191),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_201),
.B1(n_202),
.B2(n_211),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_193),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.CI(n_198),
.CON(n_193),
.SN(n_193)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_194),
.B(n_195),
.C(n_198),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_203),
.B(n_210),
.C(n_211),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_204),
.B(n_209),
.Y(n_310)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_289),
.B(n_295),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_244),
.B(n_288),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_236),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_217),
.B(n_236),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_235),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_218),
.B(n_224),
.C(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_230),
.B(n_232),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_241),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_282),
.B(n_287),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_272),
.B(n_281),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_260),
.B(n_271),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_267),
.B(n_270),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_280),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_280),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_311),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_311),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_301),
.C(n_303),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.C(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_344),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_337),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_339),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_342),
.C(n_344),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_351),
.Y(n_352)
);


endmodule