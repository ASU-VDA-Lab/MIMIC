module fake_jpeg_29528_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_51),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_25),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_55),
.B1(n_38),
.B2(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_62),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_44),
.B1(n_24),
.B2(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_18),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_35),
.C(n_17),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_99),
.B1(n_38),
.B2(n_63),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_89),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_44),
.B1(n_22),
.B2(n_24),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_68),
.B1(n_104),
.B2(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_79),
.B1(n_23),
.B2(n_40),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_32),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_36),
.B1(n_26),
.B2(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_90),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_56),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_95),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_85),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_34),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_34),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_20),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_38),
.B1(n_17),
.B2(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_23),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.Y(n_131)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_106),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_120),
.B1(n_123),
.B2(n_108),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_67),
.B(n_51),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_112),
.A2(n_125),
.B(n_40),
.C(n_37),
.D(n_31),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_67),
.C(n_63),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_93),
.C(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_94),
.B1(n_103),
.B2(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_41),
.B(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_135),
.B1(n_40),
.B2(n_37),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_45),
.B1(n_50),
.B2(n_41),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_126),
.B1(n_122),
.B2(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_70),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_145),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_110),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_83),
.B(n_41),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_165),
.B1(n_126),
.B2(n_109),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_101),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_75),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_167),
.C(n_138),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_84),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_76),
.B1(n_69),
.B2(n_102),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_45),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_124),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_128),
.B1(n_139),
.B2(n_115),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_85),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_115),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_45),
.B1(n_97),
.B2(n_82),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_96),
.B1(n_73),
.B2(n_91),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_97),
.C(n_73),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_31),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_130),
.B(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_9),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_177),
.B1(n_184),
.B2(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_136),
.B1(n_131),
.B2(n_122),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_131),
.B(n_109),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_197),
.B1(n_0),
.B2(n_16),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_113),
.B(n_138),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_165),
.B1(n_145),
.B2(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_9),
.C(n_2),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_191),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_140),
.A2(n_128),
.B1(n_139),
.B2(n_134),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_17),
.B1(n_134),
.B2(n_86),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_206),
.C(n_218),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_211),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_167),
.B1(n_141),
.B2(n_169),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_217),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_159),
.B1(n_154),
.B2(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_172),
.A2(n_106),
.B1(n_31),
.B2(n_33),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_215),
.A2(n_171),
.B1(n_170),
.B2(n_190),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_190),
.B(n_177),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_15),
.C(n_2),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_196),
.C(n_179),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_228),
.B1(n_238),
.B2(n_232),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_196),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_234),
.B1(n_200),
.B2(n_3),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_181),
.B1(n_178),
.B2(n_189),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_195),
.B(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_193),
.B1(n_195),
.B2(n_192),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_0),
.B(n_2),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_214),
.B(n_215),
.C(n_4),
.D(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_198),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_248),
.B1(n_255),
.B2(n_222),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_206),
.C(n_198),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_220),
.C(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_200),
.B1(n_213),
.B2(n_192),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_226),
.C(n_239),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_226),
.B1(n_221),
.B2(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_228),
.C(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_234),
.C(n_225),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_246),
.C(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_221),
.B1(n_250),
.B2(n_229),
.Y(n_268)
);

BUFx12f_ASAP7_75t_SL g266 ( 
.A(n_244),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_231),
.B1(n_254),
.B2(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_273),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_242),
.C(n_231),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_263),
.C(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_8),
.C(n_3),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_279),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_266),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_280),
.B(n_5),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_259),
.B(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_11),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_10),
.C(n_4),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_278),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_286),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_283),
.B(n_6),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_287),
.B(n_288),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g293 ( 
.A1(n_292),
.A2(n_12),
.B(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_0),
.B1(n_14),
.B2(n_291),
.Y(n_295)
);


endmodule