module fake_jpeg_11937_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_1),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_16),
.B(n_18),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AOI22x1_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_8),
.B1(n_12),
.B2(n_6),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_27),
.B(n_18),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_14),
.C(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.C(n_34),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_18),
.B(n_12),
.C(n_8),
.Y(n_41)
);

NAND4xp25_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_20),
.C(n_22),
.D(n_12),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_20),
.B(n_22),
.Y(n_43)
);


endmodule