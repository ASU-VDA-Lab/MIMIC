module fake_jpeg_22436_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2x1_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx2_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_55),
.Y(n_76)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_69),
.Y(n_100)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_85),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_77),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_33),
.B(n_35),
.C(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_81),
.Y(n_109)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_83),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_98),
.B1(n_31),
.B2(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_39),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AOI22x1_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_71),
.B1(n_73),
.B2(n_72),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_64),
.B1(n_53),
.B2(n_52),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_108),
.B1(n_114),
.B2(n_126),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_43),
.B1(n_45),
.B2(n_38),
.Y(n_108)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_64),
.B1(n_71),
.B2(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_89),
.B1(n_96),
.B2(n_82),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_119),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_43),
.B1(n_48),
.B2(n_37),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_28),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_124),
.Y(n_140)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_132),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_80),
.B(n_66),
.C(n_40),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_137),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_31),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_149),
.B(n_150),
.Y(n_161)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_133),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_75),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_87),
.C(n_42),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_114),
.C(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_0),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_156),
.Y(n_174)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_154),
.Y(n_185)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_116),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_129),
.B1(n_122),
.B2(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_169),
.B1(n_186),
.B2(n_139),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_115),
.B1(n_129),
.B2(n_102),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_183),
.B(n_187),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_171),
.C(n_178),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_165),
.A2(n_176),
.B1(n_23),
.B2(n_1),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_170),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_128),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_147),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_109),
.B1(n_128),
.B2(n_116),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.C(n_145),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_128),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_23),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_109),
.B1(n_122),
.B2(n_99),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_88),
.B1(n_123),
.B2(n_101),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_101),
.B1(n_121),
.B2(n_103),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_135),
.B1(n_138),
.B2(n_152),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_121),
.C(n_40),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_117),
.A3(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_42),
.C(n_84),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_19),
.C(n_18),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_84),
.B1(n_22),
.B2(n_20),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_146),
.B1(n_150),
.B2(n_156),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_117),
.B(n_22),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_191),
.B(n_203),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_210),
.B1(n_221),
.B2(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_208),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_138),
.B1(n_152),
.B2(n_148),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_158),
.B1(n_173),
.B2(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_19),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_21),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_21),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_209),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_19),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_164),
.C(n_178),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_18),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_171),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_232),
.C(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_210),
.B1(n_221),
.B2(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_161),
.B1(n_172),
.B2(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_202),
.B1(n_195),
.B2(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_187),
.C(n_1),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_10),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_238),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_16),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_0),
.C(n_2),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_246),
.C(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_2),
.C(n_4),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_258),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_191),
.C(n_215),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_211),
.B(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_201),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_200),
.C(n_205),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_268),
.C(n_224),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_234),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_196),
.B1(n_213),
.B2(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_194),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_233),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_206),
.C(n_222),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_230),
.A2(n_209),
.B1(n_5),
.B2(n_8),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_274),
.C(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_240),
.C(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_248),
.B1(n_227),
.B2(n_243),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_249),
.B1(n_267),
.B2(n_250),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_257),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_227),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_232),
.C(n_236),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_296),
.C(n_300),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_264),
.B1(n_251),
.B2(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_287),
.B1(n_279),
.B2(n_277),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_254),
.B(n_258),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_302),
.B(n_275),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_272),
.B(n_262),
.Y(n_296)
);

BUFx12_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_263),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_271),
.A2(n_209),
.B(n_255),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_285),
.B(n_270),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_310),
.B(n_289),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_275),
.C(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_286),
.B(n_255),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_209),
.C(n_256),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_256),
.C(n_5),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_5),
.C(n_6),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_298),
.C(n_299),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_6),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_6),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_316),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_321),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_297),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_322),
.A2(n_292),
.B1(n_312),
.B2(n_12),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_297),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_8),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_309),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_326),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_317),
.B(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_11),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_333),
.B(n_327),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.C(n_331),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_11),
.B(n_12),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_11),
.C(n_13),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_14),
.B(n_16),
.C(n_324),
.D(n_335),
.Y(n_341)
);


endmodule