module fake_aes_1804_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
HB1xp67_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_14), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_6), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_3), .Y(n_21) );
NOR2xp33_ASAP7_75t_SL g22 ( .A(n_10), .B(n_1), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_13), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_16), .B(n_0), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_23), .B(n_0), .Y(n_26) );
BUFx6f_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
NAND3xp33_ASAP7_75t_L g28 ( .A(n_25), .B(n_19), .C(n_18), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_24), .B(n_21), .Y(n_29) );
OAI21x1_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_17), .B(n_20), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_18), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_32), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_30), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI32xp33_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_31), .A3(n_30), .B1(n_22), .B2(n_32), .Y(n_36) );
NAND2xp5_ASAP7_75t_SL g37 ( .A(n_33), .B(n_28), .Y(n_37) );
INVxp67_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
NAND4xp25_ASAP7_75t_L g39 ( .A(n_36), .B(n_34), .C(n_29), .D(n_4), .Y(n_39) );
OAI22xp5_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_33), .B1(n_29), .B2(n_19), .Y(n_40) );
NAND4xp75_ASAP7_75t_L g41 ( .A(n_39), .B(n_33), .C(n_2), .D(n_5), .Y(n_41) );
BUFx12f_ASAP7_75t_L g42 ( .A(n_38), .Y(n_42) );
NAND4xp75_ASAP7_75t_L g43 ( .A(n_40), .B(n_1), .C(n_2), .D(n_6), .Y(n_43) );
NOR4xp25_ASAP7_75t_L g44 ( .A(n_42), .B(n_23), .C(n_27), .D(n_15), .Y(n_44) );
NAND3xp33_ASAP7_75t_L g45 ( .A(n_41), .B(n_23), .C(n_27), .Y(n_45) );
OR2x2_ASAP7_75t_SL g46 ( .A(n_45), .B(n_43), .Y(n_46) );
AOI22xp5_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_44), .B1(n_7), .B2(n_12), .Y(n_47) );
endmodule