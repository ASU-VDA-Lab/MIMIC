module real_aes_15450_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_13;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g44 ( .A(n_0), .Y(n_44) );
INVx2_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
HB1xp67_ASAP7_75t_L g45 ( .A(n_2), .Y(n_45) );
CKINVDCx20_ASAP7_75t_R g46 ( .A(n_3), .Y(n_46) );
INVx1_ASAP7_75t_L g27 ( .A(n_4), .Y(n_27) );
INVx2_ASAP7_75t_L g23 ( .A(n_5), .Y(n_23) );
BUFx3_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g39 ( .A(n_7), .Y(n_39) );
AOI32xp33_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_17), .A3(n_24), .B1(n_28), .B2(n_31), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
BUFx8_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_13), .B(n_15), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
BUFx6f_ASAP7_75t_L g30 ( .A(n_16), .Y(n_30) );
OAI21xp33_ASAP7_75t_SL g31 ( .A1(n_17), .A2(n_25), .B(n_32), .Y(n_31) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_20), .B(n_22), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
INVx1_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g40 ( .A(n_24), .B(n_41), .Y(n_40) );
INVx1_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_25), .B(n_34), .Y(n_33) );
BUFx2_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
INVx3_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_33), .B(n_40), .Y(n_32) );
INVx2_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_39), .Y(n_38) );
NOR3xp33_ASAP7_75t_L g41 ( .A(n_42), .B(n_45), .C(n_46), .Y(n_41) );
INVx2_ASAP7_75t_SL g42 ( .A(n_43), .Y(n_42) );
INVx2_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
endmodule