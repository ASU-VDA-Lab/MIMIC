module real_jpeg_12349_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_297, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_297;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_213;
wire n_128;
wire n_244;
wire n_216;
wire n_133;
wire n_179;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_28),
.B1(n_33),
.B2(n_68),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_58),
.B1(n_60),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_4),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_4),
.B(n_33),
.C(n_63),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_81),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_93),
.B(n_153),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_42),
.B(n_80),
.C(n_180),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_38),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_58),
.B1(n_60),
.B2(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_5),
.A2(n_28),
.B1(n_33),
.B2(n_83),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_57),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_28),
.B1(n_33),
.B2(n_40),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_40),
.B1(n_58),
.B2(n_60),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_58),
.B1(n_60),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_10),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_28),
.B1(n_33),
.B2(n_149),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_149),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_149),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_28),
.B1(n_33),
.B2(n_102),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_102),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_102),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_13),
.B(n_43),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_34),
.B1(n_58),
.B2(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_51),
.B1(n_58),
.B2(n_60),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_15),
.A2(n_28),
.B1(n_33),
.B2(n_51),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_51),
.Y(n_187)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_124),
.B1(n_294),
.B2(n_295),
.Y(n_18)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_19),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_105),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_21),
.B(n_105),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_87),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_70),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_36),
.B2(n_52),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_36),
.B(n_70),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_26),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_30),
.B(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_27),
.A2(n_30),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_154),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_27),
.A2(n_30),
.B1(n_92),
.B2(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx5_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_28),
.B(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_30),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_32),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_39),
.A2(n_47),
.B(n_137),
.C(n_224),
.Y(n_223)
);

AOI32xp33_ASAP7_75t_L g237 ( 
.A1(n_39),
.A2(n_42),
.A3(n_44),
.B1(n_225),
.B2(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_41),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_41),
.A2(n_45),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_41),
.A2(n_47),
.B1(n_101),
.B2(n_252),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_61),
.B1(n_69),
.B2(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_60),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_58),
.B(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_60),
.A2(n_79),
.B(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_69),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_61),
.B(n_139),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_61),
.A2(n_69),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_61),
.A2(n_69),
.B1(n_97),
.B2(n_231),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_65),
.B(n_137),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_65),
.A2(n_150),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_71),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_86),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_75),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_73),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_73),
.A2(n_138),
.B(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_76),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_76),
.A2(n_84),
.B1(n_200),
.B2(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_76),
.A2(n_186),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_81),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_77),
.B(n_187),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_81),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_84),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_84),
.A2(n_99),
.B(n_201),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_87),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.C(n_100),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_88),
.A2(n_89),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_93),
.A2(n_94),
.B1(n_182),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_93),
.A2(n_94),
.B1(n_208),
.B2(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_94),
.A2(n_159),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_137),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_94),
.A2(n_167),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_98),
.B(n_100),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_104),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_121),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_124),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_288),
.B(n_293),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_276),
.B(n_287),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_244),
.A3(n_269),
.B1(n_274),
.B2(n_275),
.C(n_297),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_217),
.B(n_243),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_194),
.B(n_216),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_175),
.B(n_193),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_155),
.B(n_174),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_151),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_147),
.C(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_163),
.B(n_173),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_161),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_172),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_188),
.C(n_192),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_181),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_209),
.B2(n_210),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_212),
.C(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_203),
.C(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_234),
.C(n_235),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_232),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_227),
.C(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_259),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_255),
.C(n_258),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_247),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_253),
.C(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_268),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_263),
.C(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_286),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);


endmodule