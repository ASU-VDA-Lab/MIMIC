module fake_aes_5000_n_17 (n_1, n_2, n_4, n_3, n_0, n_17);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_1), .B(n_2), .Y(n_6) );
BUFx6f_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI21x1_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_6), .B(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
INVxp67_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_12), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_14), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
endmodule