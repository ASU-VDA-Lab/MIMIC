module fake_jpeg_2323_n_105 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_40),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_38),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_33),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_50),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_48),
.B1(n_45),
.B2(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_54),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_1),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_82),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_28),
.B(n_3),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_10),
.B(n_11),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_81),
.B1(n_76),
.B2(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_19),
.C2(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_24),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_89),
.C(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_94),
.C(n_93),
.Y(n_103)
);

INVxp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_91),
.Y(n_105)
);


endmodule