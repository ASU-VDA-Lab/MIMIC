module fake_jpeg_21039_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_23),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_26),
.B1(n_15),
.B2(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_15),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_52),
.B1(n_40),
.B2(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_15),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_30),
.B1(n_22),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_79),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_19),
.B1(n_25),
.B2(n_22),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_66),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_40),
.B1(n_39),
.B2(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_67),
.B1(n_80),
.B2(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_37),
.B1(n_33),
.B2(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_78),
.B1(n_49),
.B2(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_35),
.B(n_2),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_35),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_16),
.B1(n_20),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_24),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_24),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_66),
.B1(n_74),
.B2(n_76),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_51),
.B(n_50),
.C(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_31),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_41),
.C(n_33),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_60),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_113),
.B1(n_71),
.B2(n_41),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_74),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_123),
.B(n_128),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_80),
.B1(n_58),
.B2(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_72),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_94),
.C(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_65),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_67),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_88),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_35),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_129),
.B(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_13),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_140),
.B(n_111),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_136),
.C(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_98),
.C(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_104),
.B(n_35),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_104),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_97),
.C(n_62),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_61),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_101),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_1),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_127),
.C(n_113),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_126),
.B1(n_116),
.B2(n_109),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_165),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_116),
.B1(n_106),
.B2(n_119),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_81),
.B1(n_105),
.B2(n_50),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_114),
.B1(n_127),
.B2(n_117),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_137),
.B1(n_140),
.B2(n_151),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_152),
.B1(n_120),
.B2(n_107),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_147),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_150),
.Y(n_175)
);

XOR2x1_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_138),
.C(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_181),
.C(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_97),
.C(n_81),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_70),
.B1(n_3),
.B2(n_4),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_174),
.B1(n_162),
.B2(n_180),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_35),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_167),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_156),
.C(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_196),
.B1(n_197),
.B2(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_8),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_155),
.B(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_195),
.B1(n_176),
.B2(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_168),
.C(n_165),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_175),
.C(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_177),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_5),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_179),
.C(n_165),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_70),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_206),
.B1(n_198),
.B2(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_6),
.C(n_8),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_216),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_198),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_204),
.B(n_209),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_210),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_227),
.A3(n_215),
.B1(n_225),
.B2(n_199),
.C1(n_223),
.C2(n_202),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_229),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_10),
.B(n_11),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_11),
.Y(n_232)
);


endmodule