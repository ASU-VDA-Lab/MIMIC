module fake_netlist_5_992_n_1821 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1821);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1821;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_60),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_56),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_99),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_110),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_18),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_64),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_40),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_93),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_100),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_34),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_45),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_126),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_15),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_71),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_53),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_53),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_116),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_34),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_70),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_58),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_167),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_112),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_58),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_105),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_83),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_63),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_43),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_6),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_37),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_109),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_123),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_52),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_12),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_38),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_139),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_48),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_85),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_69),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_46),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_90),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_134),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_66),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_7),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_124),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_30),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_113),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_23),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_152),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_75),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_42),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_114),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_87),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_102),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_140),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_157),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_136),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_104),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_65),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_117),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_23),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_59),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_47),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_35),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_84),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_129),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_22),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_148),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_106),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_20),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_47),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_44),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_151),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_103),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_165),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_56),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_150),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_171),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_121),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_173),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_33),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_67),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_60),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_144),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_50),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_74),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_31),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_62),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_32),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_79),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_95),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_0),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_33),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_156),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_159),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_17),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_89),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_25),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_119),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_13),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_20),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_4),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_16),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_128),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_52),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_168),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_51),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_5),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_41),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_204),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_183),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_331),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_174),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_179),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_254),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_183),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_196),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_204),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_204),
.Y(n_365)
);

BUFx2_ASAP7_75t_SL g366 ( 
.A(n_227),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_204),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_204),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_204),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_220),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_231),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_220),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_232),
.Y(n_375)
);

BUFx2_ASAP7_75t_SL g376 ( 
.A(n_257),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_220),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_243),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_220),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_220),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_332),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_263),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_198),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_211),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_219),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_184),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_258),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_252),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_282),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_184),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_222),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_225),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_280),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_226),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_334),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_250),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_250),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_251),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_175),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_251),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_253),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_253),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_256),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_256),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_266),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_229),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_294),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_266),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_192),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_234),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_192),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_194),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_186),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_235),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_199),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_206),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_207),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_238),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_255),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_260),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_195),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_252),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_278),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_339),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_291),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_351),
.B(n_175),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_358),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_356),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_409),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_180),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_374),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_388),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_390),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_361),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_372),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_400),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_373),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_351),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_188),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_188),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_378),
.B(n_180),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_401),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_353),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_380),
.B(n_314),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_403),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_357),
.B(n_214),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_181),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_383),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_362),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_359),
.A2(n_350),
.B1(n_212),
.B2(n_305),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_364),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_384),
.B(n_314),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_387),
.B(n_389),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_315),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_363),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_363),
.B(n_315),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_419),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_393),
.B(n_317),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_364),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_365),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_317),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_365),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_382),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_421),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_360),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_367),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_367),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_369),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_398),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_369),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_368),
.A2(n_289),
.B1(n_262),
.B2(n_346),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_370),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_404),
.B(n_181),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_416),
.Y(n_516)
);

AND3x2_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_297),
.C(n_435),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_443),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_493),
.B(n_385),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_493),
.B(n_395),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_451),
.B(n_487),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_467),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_489),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_467),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_422),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_448),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_516),
.B(n_402),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_472),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_491),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_512),
.B(n_475),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_452),
.B(n_427),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_487),
.B(n_370),
.C(n_426),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_449),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_497),
.B(n_176),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_491),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_468),
.B(n_218),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_492),
.A2(n_237),
.B1(n_324),
.B2(n_190),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_468),
.B(n_239),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_424),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_479),
.A2(n_236),
.B1(n_242),
.B2(n_210),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_478),
.B(n_288),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_458),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_454),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_458),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_465),
.A2(n_425),
.B(n_182),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_478),
.B(n_312),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_464),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_439),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_479),
.A2(n_304),
.B1(n_268),
.B2(n_259),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_455),
.B(n_352),
.Y(n_573)
);

AND3x2_ASAP7_75t_L g574 ( 
.A(n_439),
.B(n_423),
.C(n_420),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_492),
.B(n_497),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_482),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_478),
.B(n_248),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_476),
.B(n_185),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_449),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_461),
.B(n_391),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_471),
.B(n_399),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_482),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_SL g585 ( 
.A(n_513),
.B(n_247),
.C(n_354),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_486),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_474),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_495),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_501),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_476),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_513),
.A2(n_318),
.B1(n_195),
.B2(n_261),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_486),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_498),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_475),
.B(n_434),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_502),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_497),
.B(n_177),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_486),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_515),
.B(n_237),
.C(n_190),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_486),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_515),
.B(n_214),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_500),
.B(n_366),
.Y(n_607)
);

AND2x2_ASAP7_75t_SL g608 ( 
.A(n_441),
.B(n_193),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_500),
.B(n_366),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_445),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_456),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

BUFx8_ASAP7_75t_SL g614 ( 
.A(n_460),
.Y(n_614)
);

CKINVDCx6p67_ASAP7_75t_R g615 ( 
.A(n_470),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_499),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_506),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_450),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_507),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_450),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_465),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_450),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_500),
.A2(n_241),
.B1(n_228),
.B2(n_224),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_465),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_447),
.B(n_376),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_447),
.B(n_376),
.Y(n_632)
);

AND3x2_ASAP7_75t_L g633 ( 
.A(n_465),
.B(n_208),
.C(n_205),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_465),
.B(n_424),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_466),
.A2(n_324),
.B1(n_292),
.B2(n_295),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_514),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_514),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_514),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_440),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_466),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_464),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_R g645 ( 
.A(n_466),
.B(n_185),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_440),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_447),
.B(n_405),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_496),
.B(n_446),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_457),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_466),
.B(n_473),
.Y(n_650)
);

AOI21x1_ASAP7_75t_L g651 ( 
.A1(n_483),
.A2(n_425),
.B(n_217),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_473),
.B(n_406),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_457),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_459),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_442),
.B(n_187),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_459),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_463),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_463),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_469),
.Y(n_659)
);

OAI22x1_ASAP7_75t_L g660 ( 
.A1(n_473),
.A2(n_261),
.B1(n_318),
.B2(n_322),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_473),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_473),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_446),
.B(n_264),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_521),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_538),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_638),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_593),
.B(n_189),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_593),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_599),
.B(n_447),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_538),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_662),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_551),
.A2(n_437),
.B1(n_298),
.B2(n_287),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_579),
.A2(n_320),
.B(n_348),
.C(n_336),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_592),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_554),
.B(n_189),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_576),
.B(n_464),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_521),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_534),
.B(n_191),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_607),
.B(n_191),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_464),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_629),
.B(n_464),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_608),
.B(n_462),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_592),
.B(n_426),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_609),
.B(n_540),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_197),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_540),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_559),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_608),
.B(n_441),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_558),
.B(n_569),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_608),
.B(n_462),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_625),
.B(n_462),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_625),
.B(n_462),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_650),
.B(n_446),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_662),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_550),
.B(n_283),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_572),
.B(n_606),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_586),
.A2(n_299),
.B1(n_274),
.B2(n_213),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_652),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_550),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_586),
.A2(n_483),
.B(n_442),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_585),
.B(n_233),
.C(n_221),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_604),
.B(n_209),
.C(n_201),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_663),
.B(n_441),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_197),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_547),
.A2(n_349),
.B1(n_306),
.B2(n_442),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_522),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_536),
.B(n_214),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_519),
.B(n_200),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_595),
.B(n_441),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_614),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_595),
.B(n_441),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_600),
.B(n_494),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_600),
.B(n_494),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_535),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_519),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_603),
.B(n_494),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_603),
.B(n_605),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_647),
.B(n_200),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_605),
.Y(n_723)
);

OAI221xp5_ASAP7_75t_L g724 ( 
.A1(n_553),
.A2(n_547),
.B1(n_594),
.B2(n_556),
.C(n_543),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_566),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_283),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_530),
.B(n_319),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_530),
.B(n_319),
.Y(n_728)
);

OAI221xp5_ASAP7_75t_L g729 ( 
.A1(n_594),
.A2(n_249),
.B1(n_246),
.B2(n_244),
.C(n_311),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_635),
.B(n_494),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_578),
.B(n_194),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_635),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_530),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_649),
.B(n_494),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_649),
.B(n_442),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_656),
.B(n_442),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_637),
.A2(n_442),
.B1(n_240),
.B2(n_194),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_656),
.B(n_442),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_630),
.B(n_321),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_645),
.A2(n_276),
.B1(n_265),
.B2(n_267),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_643),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_657),
.B(n_442),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_632),
.B(n_321),
.Y(n_744)
);

BUFx5_ASAP7_75t_L g745 ( 
.A(n_524),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_658),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_658),
.B(n_477),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_659),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_661),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_628),
.B(n_323),
.Y(n_750)
);

INVxp67_ASAP7_75t_SL g751 ( 
.A(n_575),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_559),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_661),
.B(n_480),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_559),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_549),
.B(n_480),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_637),
.A2(n_240),
.B1(n_194),
.B2(n_347),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_549),
.A2(n_273),
.B1(n_345),
.B2(n_337),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_642),
.Y(n_758)
);

HB1xp67_ASAP7_75t_SL g759 ( 
.A(n_612),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_587),
.B(n_215),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_642),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_549),
.B(n_484),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_549),
.B(n_484),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_646),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_602),
.A2(n_335),
.B(n_329),
.C(n_508),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_602),
.B(n_485),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_544),
.B(n_323),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_646),
.Y(n_768)
);

AO221x1_ASAP7_75t_L g769 ( 
.A1(n_557),
.A2(n_660),
.B1(n_637),
.B2(n_520),
.C(n_541),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_602),
.B(n_655),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_653),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_602),
.B(n_485),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_637),
.A2(n_194),
.B1(n_240),
.B2(n_322),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_560),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_612),
.B(n_428),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_573),
.A2(n_333),
.B1(n_330),
.B2(n_327),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_653),
.B(n_488),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_560),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_571),
.B(n_428),
.Y(n_779)
);

AND2x6_ASAP7_75t_L g780 ( 
.A(n_575),
.B(n_450),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_660),
.A2(n_194),
.B1(n_240),
.B2(n_325),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_587),
.B(n_429),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_654),
.B(n_488),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_581),
.A2(n_582),
.B1(n_610),
.B2(n_623),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_587),
.B(n_326),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_567),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_524),
.A2(n_511),
.B(n_510),
.C(n_508),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_664),
.B(n_490),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_567),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_527),
.B(n_504),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_532),
.B(n_505),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_634),
.A2(n_240),
.B1(n_327),
.B2(n_325),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_567),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_537),
.B(n_326),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_575),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_539),
.B(n_510),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_634),
.B(n_240),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_523),
.B(n_328),
.C(n_438),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_539),
.A2(n_328),
.B1(n_286),
.B2(n_310),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_SL g801 ( 
.A(n_587),
.B(n_215),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_525),
.B(n_269),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_518),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_517),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_546),
.B(n_555),
.Y(n_805)
);

BUFx6f_ASAP7_75t_SL g806 ( 
.A(n_615),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_618),
.B(n_429),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_618),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_546),
.B(n_216),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_555),
.A2(n_511),
.B(n_430),
.C(n_438),
.Y(n_810)
);

XOR2xp5_ASAP7_75t_L g811 ( 
.A(n_615),
.B(n_275),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_520),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_574),
.B(n_430),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_SL g814 ( 
.A(n_633),
.B(n_215),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_561),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_561),
.Y(n_816)
);

BUFx6f_ASAP7_75t_SL g817 ( 
.A(n_565),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_565),
.B(n_223),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_583),
.A2(n_279),
.B1(n_281),
.B2(n_284),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_583),
.B(n_450),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_584),
.B(n_431),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_636),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_584),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_588),
.A2(n_302),
.B1(n_307),
.B2(n_301),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_588),
.B(n_450),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_723),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_718),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_699),
.B(n_518),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_769),
.A2(n_617),
.B1(n_596),
.B2(n_597),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_773),
.A2(n_617),
.B1(n_596),
.B2(n_597),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_SL g831 ( 
.A(n_729),
.B(n_333),
.C(n_330),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_702),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_681),
.B(n_589),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_725),
.B(n_651),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_780),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_681),
.B(n_589),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_669),
.B(n_590),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_742),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_758),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_759),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_699),
.B(n_518),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_739),
.B(n_746),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_770),
.B(n_518),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_713),
.B(n_245),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_748),
.B(n_590),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_761),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_676),
.B(n_431),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_764),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_732),
.A2(n_598),
.B1(n_616),
.B2(n_611),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_770),
.B(n_518),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_749),
.B(n_598),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_670),
.B(n_601),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_768),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_771),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_685),
.B(n_518),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_787),
.B(n_601),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_671),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_672),
.B(n_697),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_693),
.B(n_564),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_721),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_667),
.B(n_432),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_812),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_815),
.B(n_611),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_619),
.B1(n_616),
.B2(n_631),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_684),
.A2(n_683),
.B(n_678),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_815),
.B(n_619),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_823),
.B(n_701),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_812),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_806),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_665),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_745),
.B(n_564),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_745),
.B(n_564),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_671),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_816),
.Y(n_874)
);

AND2x4_ASAP7_75t_SL g875 ( 
.A(n_702),
.B(n_230),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_631),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_719),
.A2(n_639),
.B1(n_640),
.B2(n_626),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_808),
.B(n_760),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_775),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_SL g880 ( 
.A(n_704),
.B(n_277),
.C(n_270),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_696),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_R g882 ( 
.A(n_807),
.B(n_271),
.Y(n_882)
);

AND2x6_ASAP7_75t_SL g883 ( 
.A(n_775),
.B(n_432),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_673),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_822),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_821),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_733),
.B(n_639),
.Y(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_780),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_775),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_715),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_679),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_782),
.A2(n_640),
.B1(n_644),
.B2(n_570),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_716),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_720),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_L g895 ( 
.A(n_686),
.B(n_272),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_676),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_724),
.B(n_562),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_801),
.A2(n_230),
.B1(n_343),
.B2(n_342),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_773),
.A2(n_240),
.B1(n_641),
.B2(n_577),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_718),
.B(n_689),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_718),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_751),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_690),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_688),
.B(n_641),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_688),
.B(n_577),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_718),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_755),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_752),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_809),
.B(n_577),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_754),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_809),
.B(n_591),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_742),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_709),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_781),
.A2(n_240),
.B1(n_622),
.B2(n_621),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_767),
.A2(n_562),
.B1(n_644),
.B2(n_570),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_671),
.B(n_564),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_671),
.Y(n_917)
);

AO22x1_ASAP7_75t_L g918 ( 
.A1(n_704),
.A2(n_341),
.B1(n_340),
.B2(n_290),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_762),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_742),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_806),
.B(n_651),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_818),
.B(n_591),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_774),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_726),
.B(n_433),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_818),
.B(n_591),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_SL g926 ( 
.A(n_668),
.B(n_303),
.C(n_309),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_680),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_698),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_778),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_763),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_786),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_780),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_766),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_680),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_779),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_817),
.B(n_564),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_687),
.B(n_562),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_680),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_666),
.B(n_613),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_804),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_691),
.A2(n_520),
.B1(n_627),
.B2(n_541),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_811),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_745),
.B(n_691),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_813),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_796),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_790),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_772),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_666),
.B(n_613),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_730),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_777),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_784),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_794),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_745),
.B(n_620),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_783),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_780),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_784),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_745),
.B(n_620),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_803),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_709),
.B(n_562),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_781),
.A2(n_621),
.B1(n_622),
.B2(n_230),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_710),
.B(n_285),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_805),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_734),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_747),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_707),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_799),
.B(n_433),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_784),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_820),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_706),
.A2(n_644),
.B(n_626),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_799),
.B(n_436),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_756),
.A2(n_622),
.B1(n_542),
.B2(n_533),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_753),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_788),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_767),
.A2(n_644),
.B1(n_570),
.B2(n_626),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_802),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_677),
.Y(n_976)
);

AO22x1_ASAP7_75t_L g977 ( 
.A1(n_795),
.A2(n_717),
.B1(n_727),
.B2(n_728),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_791),
.Y(n_978)
);

AND2x6_ASAP7_75t_L g979 ( 
.A(n_735),
.B(n_520),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_825),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_717),
.B(n_436),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_711),
.B(n_541),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_736),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_750),
.B(n_570),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_738),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_792),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_817),
.B(n_568),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_797),
.Y(n_988)
);

NOR2x2_ASAP7_75t_L g989 ( 
.A(n_776),
.B(n_529),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_743),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_798),
.Y(n_991)
);

NOR2x1p5_ASAP7_75t_L g992 ( 
.A(n_705),
.B(n_293),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_795),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_712),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_727),
.B(n_406),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_728),
.B(n_627),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_714),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_789),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_675),
.B(n_407),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_694),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_803),
.B(n_563),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_785),
.B(n_407),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_810),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_977),
.B(n_722),
.C(n_682),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_SL g1005 ( 
.A(n_878),
.B(n_814),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_917),
.B(n_626),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_865),
.A2(n_695),
.B(n_703),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_913),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_828),
.A2(n_744),
.B(n_740),
.C(n_700),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_965),
.B(n_674),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_965),
.B(n_741),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_928),
.A2(n_757),
.B1(n_824),
.B2(n_819),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_944),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_998),
.B(n_793),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_912),
.B(n_765),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_832),
.B(n_800),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_827),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_945),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_993),
.B(n_793),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_902),
.A2(n_756),
.B1(n_708),
.B2(n_737),
.Y(n_1020)
);

NOR2x1_ASAP7_75t_L g1021 ( 
.A(n_912),
.B(n_731),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_964),
.B(n_708),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_896),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_874),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_847),
.B(n_737),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_993),
.B(n_928),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_839),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_897),
.A2(n_541),
.B(n_627),
.C(n_624),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_945),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_880),
.A2(n_956),
.B(n_967),
.C(n_951),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_848),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_838),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_838),
.B(n_920),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_853),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_827),
.Y(n_1035)
);

AO32x2_ASAP7_75t_L g1036 ( 
.A1(n_941),
.A2(n_780),
.A3(n_568),
.B1(n_2),
.B2(n_3),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_900),
.B(n_408),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_916),
.A2(n_620),
.B(n_563),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_SL g1039 ( 
.A(n_926),
.B(n_296),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_SL g1040 ( 
.A(n_835),
.B(n_531),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_852),
.A2(n_624),
.B(n_580),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_854),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_978),
.B(n_548),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_832),
.B(n_300),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_897),
.A2(n_907),
.B(n_930),
.C(n_919),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_969),
.A2(n_580),
.B(n_552),
.Y(n_1046)
);

OAI22x1_ASAP7_75t_L g1047 ( 
.A1(n_879),
.A2(n_308),
.B1(n_313),
.B2(n_408),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_826),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_838),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_841),
.A2(n_531),
.B(n_533),
.C(n_545),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_840),
.Y(n_1051)
);

OAI21xp33_ASAP7_75t_SL g1052 ( 
.A1(n_841),
.A2(n_580),
.B(n_552),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_829),
.A2(n_418),
.B(n_415),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_962),
.A2(n_418),
.B1(n_415),
.B2(n_414),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_935),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_827),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_986),
.B(n_414),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_984),
.A2(n_413),
.B(n_412),
.C(n_411),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_867),
.A2(n_413),
.B(n_412),
.C(n_411),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_860),
.A2(n_410),
.B1(n_1),
.B2(n_2),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_896),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_949),
.A2(n_410),
.B1(n_8),
.B2(n_10),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_944),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_870),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_939),
.A2(n_162),
.B(n_161),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_842),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_976),
.A2(n_153),
.B1(n_149),
.B2(n_146),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_845),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_858),
.B(n_145),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_851),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_933),
.A2(n_0),
.B(n_8),
.C(n_10),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_858),
.B(n_924),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_948),
.A2(n_143),
.B(n_135),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_947),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_920),
.B(n_131),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_988),
.B(n_14),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_884),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_830),
.A2(n_963),
.B1(n_899),
.B2(n_890),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_889),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_975),
.A2(n_130),
.B1(n_125),
.B2(n_120),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_891),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_903),
.Y(n_1082)
);

BUFx8_ASAP7_75t_SL g1083 ( 
.A(n_869),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_972),
.B(n_97),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_901),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_981),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_829),
.A2(n_96),
.B(n_91),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_901),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_835),
.A2(n_78),
.B(n_77),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_924),
.A2(n_995),
.B1(n_895),
.B2(n_894),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_901),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_972),
.B(n_17),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_950),
.B(n_19),
.Y(n_1093)
);

INVx8_ASAP7_75t_L g1094 ( 
.A(n_940),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_846),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_954),
.B(n_22),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_995),
.B(n_76),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_861),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_861),
.B(n_24),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_830),
.A2(n_899),
.B1(n_893),
.B2(n_837),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_885),
.B(n_25),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_886),
.B(n_26),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_843),
.A2(n_26),
.B(n_27),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_837),
.B(n_28),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_883),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_835),
.A2(n_61),
.B(n_31),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_875),
.B(n_29),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_908),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_942),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_910),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_875),
.B(n_29),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_992),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_882),
.B(n_36),
.C(n_37),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_923),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_843),
.A2(n_36),
.B(n_41),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_929),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_959),
.B(n_43),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_881),
.A2(n_45),
.B(n_49),
.C(n_54),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_834),
.B(n_54),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_833),
.A2(n_836),
.B1(n_997),
.B2(n_994),
.Y(n_1120)
);

AO32x2_ASAP7_75t_L g1121 ( 
.A1(n_989),
.A2(n_55),
.A3(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_989),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_959),
.B(n_55),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_937),
.A2(n_57),
.B(n_831),
.C(n_990),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_994),
.B(n_1000),
.Y(n_1125)
);

AND2x6_ASAP7_75t_L g1126 ( 
.A(n_955),
.B(n_985),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_906),
.Y(n_1127)
);

AO32x2_ASAP7_75t_L g1128 ( 
.A1(n_855),
.A2(n_859),
.A3(n_850),
.B1(n_914),
.B2(n_960),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_961),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_L g1130 ( 
.A(n_966),
.B(n_970),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_863),
.B(n_866),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_876),
.B(n_904),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_966),
.B(n_970),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1002),
.B(n_898),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_834),
.B(n_898),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_857),
.B(n_873),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_942),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1002),
.B(n_918),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_931),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_882),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_850),
.A2(n_855),
.B(n_859),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_946),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_987),
.B(n_926),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_936),
.B(n_927),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1002),
.A2(n_960),
.B1(n_973),
.B2(n_999),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1134),
.B(n_831),
.C(n_937),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1046),
.A2(n_953),
.B(n_957),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1045),
.A2(n_905),
.B(n_922),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1100),
.A2(n_914),
.B1(n_971),
.B2(n_856),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1027),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1008),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_L g1152 ( 
.A(n_1032),
.B(n_921),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1007),
.A2(n_888),
.B(n_932),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1086),
.B(n_983),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1140),
.B(n_862),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1120),
.A2(n_1100),
.B(n_1132),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1120),
.A2(n_911),
.B(n_909),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1031),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1034),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1042),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1087),
.A2(n_971),
.B1(n_925),
.B2(n_892),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1117),
.A2(n_982),
.B(n_996),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1061),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_906),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_SL g1165 ( 
.A(n_1005),
.B(n_961),
.C(n_921),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1050),
.A2(n_872),
.B(n_871),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1068),
.B(n_980),
.Y(n_1167)
);

NOR2xp67_ASAP7_75t_SL g1168 ( 
.A(n_1032),
.B(n_1051),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1141),
.A2(n_864),
.B(n_887),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1072),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_L g1171 ( 
.A1(n_1123),
.A2(n_936),
.B(n_871),
.C(n_953),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1024),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1141),
.A2(n_915),
.B(n_974),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1131),
.A2(n_958),
.B(n_1001),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1070),
.B(n_968),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1032),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1066),
.B(n_985),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1029),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1125),
.B(n_1025),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1078),
.B(n_868),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1028),
.A2(n_1003),
.A3(n_991),
.B(n_952),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1078),
.B(n_927),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1104),
.A2(n_1004),
.B(n_1135),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1035),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1124),
.A2(n_979),
.A3(n_877),
.B(n_999),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1087),
.A2(n_849),
.B1(n_906),
.B2(n_934),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1020),
.A2(n_979),
.A3(n_999),
.B(n_987),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1072),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1048),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1086),
.B(n_844),
.Y(n_1190)
);

AO32x2_ASAP7_75t_L g1191 ( 
.A1(n_1145),
.A2(n_979),
.A3(n_906),
.B1(n_934),
.B2(n_938),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1095),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1005),
.B(n_934),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1022),
.B(n_934),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1075),
.B(n_958),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1136),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1009),
.A2(n_979),
.B(n_1052),
.Y(n_1197)
);

NAND3xp33_ASAP7_75t_L g1198 ( 
.A(n_1010),
.B(n_1113),
.C(n_1004),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1110),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1139),
.Y(n_1200)
);

BUFx12f_ASAP7_75t_L g1201 ( 
.A(n_1129),
.Y(n_1201)
);

AOI221x1_ASAP7_75t_L g1202 ( 
.A1(n_1062),
.A2(n_1060),
.B1(n_1039),
.B2(n_1071),
.C(n_1074),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1040),
.A2(n_1118),
.A3(n_1062),
.B(n_1060),
.Y(n_1203)
);

AOI221x1_ASAP7_75t_L g1204 ( 
.A1(n_1047),
.A2(n_1106),
.B1(n_1092),
.B2(n_1011),
.C(n_1076),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1057),
.B(n_1133),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1130),
.B(n_1049),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1065),
.A2(n_1073),
.B(n_1038),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1084),
.A2(n_1097),
.B(n_1006),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1064),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1023),
.B(n_1122),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1043),
.A2(n_1016),
.A3(n_1101),
.B(n_1128),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1023),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1094),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1019),
.B(n_1077),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1081),
.B(n_1116),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1017),
.B(n_1056),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1082),
.B(n_1142),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1055),
.B(n_1119),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_SL g1220 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_1053),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1021),
.A2(n_1015),
.B(n_1053),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1128),
.A2(n_1054),
.A3(n_1089),
.B(n_1036),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1108),
.B(n_1114),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1012),
.A2(n_1090),
.B(n_1138),
.C(n_1143),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1079),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1058),
.A2(n_1059),
.B(n_1126),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1013),
.Y(n_1227)
);

NAND3x1_ASAP7_75t_L g1228 ( 
.A(n_1107),
.B(n_1111),
.C(n_1102),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1083),
.Y(n_1229)
);

AOI31xp67_ASAP7_75t_L g1230 ( 
.A1(n_1080),
.A2(n_1067),
.A3(n_1026),
.B(n_1036),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1033),
.B(n_1098),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_1017),
.B(n_1091),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1128),
.A2(n_1037),
.B(n_1036),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1037),
.A2(n_1112),
.B(n_1063),
.Y(n_1235)
);

AO32x2_ASAP7_75t_L g1236 ( 
.A1(n_1121),
.A2(n_1091),
.A3(n_1056),
.B1(n_1144),
.B2(n_1126),
.Y(n_1236)
);

AO32x2_ASAP7_75t_L g1237 ( 
.A1(n_1121),
.A2(n_1126),
.A3(n_1044),
.B1(n_1099),
.B2(n_1088),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1121),
.A2(n_1069),
.B(n_1099),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1069),
.B(n_1137),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1035),
.A2(n_1085),
.B(n_1088),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_SL g1241 ( 
.A1(n_1035),
.A2(n_1085),
.B(n_1088),
.C(n_1127),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1094),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1085),
.B(n_1127),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1033),
.A2(n_1127),
.B1(n_1105),
.B2(n_1109),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1094),
.A2(n_1046),
.B(n_865),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1045),
.A2(n_1028),
.A3(n_897),
.B(n_1100),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1072),
.B(n_1130),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1008),
.Y(n_1248)
);

O2A1O1Ixp5_ASAP7_75t_L g1249 ( 
.A1(n_1117),
.A2(n_977),
.B(n_1123),
.C(n_722),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1086),
.B(n_782),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1032),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_1109),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1068),
.B(n_998),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_1087),
.A2(n_1123),
.B(n_1117),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1045),
.A2(n_897),
.B(n_865),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1046),
.A2(n_865),
.B(n_1041),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1068),
.B(n_998),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1068),
.B(n_998),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1068),
.B(n_998),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_SL g1260 ( 
.A1(n_1045),
.A2(n_1087),
.B(n_1124),
.C(n_1014),
.Y(n_1260)
);

BUFx2_ASAP7_75t_R g1261 ( 
.A(n_1083),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1068),
.B(n_998),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1100),
.A2(n_1087),
.B1(n_998),
.B2(n_1066),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1027),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1061),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1007),
.A2(n_943),
.B(n_865),
.Y(n_1266)
);

NAND2x1_ASAP7_75t_L g1267 ( 
.A(n_1126),
.B(n_917),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1136),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1007),
.A2(n_943),
.B(n_865),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1141),
.A2(n_1045),
.B(n_1007),
.Y(n_1270)
);

O2A1O1Ixp5_ASAP7_75t_L g1271 ( 
.A1(n_1117),
.A2(n_977),
.B(n_1123),
.C(n_722),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1008),
.Y(n_1272)
);

O2A1O1Ixp5_ASAP7_75t_L g1273 ( 
.A1(n_1117),
.A2(n_977),
.B(n_1123),
.C(n_722),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1032),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1061),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1007),
.A2(n_841),
.B(n_828),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1087),
.A2(n_1124),
.B1(n_1123),
.B2(n_1117),
.C(n_1134),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1008),
.Y(n_1278)
);

NAND3x1_ASAP7_75t_L g1279 ( 
.A(n_1134),
.B(n_594),
.C(n_599),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1086),
.B(n_782),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1086),
.B(n_782),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1018),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1007),
.A2(n_841),
.B(n_828),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1045),
.A2(n_897),
.B(n_865),
.Y(n_1284)
);

NOR2x1_ASAP7_75t_SL g1285 ( 
.A(n_1100),
.B(n_835),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1068),
.B(n_998),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1086),
.B(n_782),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1045),
.A2(n_897),
.B(n_865),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1150),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1277),
.A2(n_1271),
.B(n_1249),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1255),
.A2(n_1288),
.B(n_1284),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1198),
.B(n_1254),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1255),
.A2(n_1288),
.B(n_1284),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1153),
.A2(n_1269),
.B(n_1266),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1197),
.A2(n_1157),
.B(n_1148),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1211),
.B(n_1154),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1279),
.A2(n_1262),
.B1(n_1286),
.B2(n_1253),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1160),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_L g1301 ( 
.A(n_1273),
.B(n_1204),
.C(n_1146),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1247),
.B(n_1206),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1250),
.B(n_1280),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1242),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1147),
.A2(n_1283),
.B(n_1276),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1176),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1183),
.A2(n_1166),
.B(n_1182),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1151),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1182),
.A2(n_1171),
.B(n_1220),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1264),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1179),
.B(n_1263),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1226),
.A2(n_1221),
.B(n_1180),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1263),
.A2(n_1161),
.B(n_1162),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1213),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1176),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1260),
.A2(n_1224),
.B(n_1208),
.C(n_1205),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1241),
.A2(n_1226),
.B(n_1174),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1180),
.A2(n_1202),
.B(n_1162),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1214),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1165),
.A2(n_1228),
.B1(n_1190),
.B2(n_1239),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1176),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1195),
.A2(n_1149),
.B(n_1286),
.C(n_1257),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1189),
.Y(n_1323)
);

INVx3_ASAP7_75t_SL g1324 ( 
.A(n_1229),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1178),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1253),
.A2(n_1262),
.B1(n_1259),
.B2(n_1258),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1248),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1194),
.A2(n_1186),
.B(n_1267),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1282),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1278),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1205),
.B(n_1219),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1208),
.A2(n_1215),
.B(n_1238),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1257),
.A2(n_1258),
.B1(n_1259),
.B2(n_1281),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1167),
.A2(n_1175),
.B1(n_1179),
.B2(n_1177),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1209),
.B(n_1164),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1177),
.B(n_1175),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1192),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1235),
.A2(n_1193),
.B1(n_1275),
.B2(n_1265),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1287),
.B(n_1188),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1201),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1230),
.A2(n_1215),
.B(n_1169),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1233),
.A2(n_1240),
.B(n_1172),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1247),
.A2(n_1244),
.B1(n_1252),
.B2(n_1170),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1167),
.A2(n_1155),
.B1(n_1244),
.B2(n_1163),
.C(n_1225),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1199),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1200),
.A2(n_1173),
.B1(n_1234),
.B2(n_1270),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1261),
.Y(n_1347)
);

AO32x2_ASAP7_75t_L g1348 ( 
.A1(n_1237),
.A2(n_1236),
.A3(n_1191),
.B1(n_1234),
.B2(n_1212),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1216),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1272),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1285),
.A2(n_1237),
.B1(n_1236),
.B2(n_1232),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1218),
.A2(n_1223),
.B(n_1232),
.Y(n_1352)
);

AOI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1227),
.A2(n_1231),
.B1(n_1218),
.B2(n_1223),
.C(n_1206),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1232),
.B(n_1168),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1152),
.B(n_1268),
.C(n_1196),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1243),
.B(n_1231),
.Y(n_1356)
);

CKINVDCx6p67_ASAP7_75t_R g1357 ( 
.A(n_1251),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1217),
.A2(n_1203),
.B(n_1246),
.C(n_1185),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1203),
.A2(n_1246),
.B(n_1185),
.C(n_1187),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1251),
.B(n_1274),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1181),
.A2(n_1185),
.B(n_1187),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1251),
.B(n_1274),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1237),
.A2(n_1236),
.B(n_1191),
.C(n_1222),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1222),
.A2(n_1191),
.B(n_1184),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1213),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1210),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1254),
.A2(n_1249),
.B(n_1273),
.C(n_1271),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1150),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1150),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1254),
.A2(n_1285),
.A3(n_1277),
.B(n_1263),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1249),
.A2(n_1273),
.B(n_1271),
.C(n_1254),
.Y(n_1371)
);

NAND2xp33_ASAP7_75t_L g1372 ( 
.A(n_1279),
.B(n_725),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1229),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1150),
.Y(n_1374)
);

BUFx2_ASAP7_75t_R g1375 ( 
.A(n_1229),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1150),
.Y(n_1376)
);

AO32x2_ASAP7_75t_L g1377 ( 
.A1(n_1263),
.A2(n_956),
.A3(n_967),
.B1(n_951),
.B2(n_1062),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1195),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1210),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1279),
.A2(n_1087),
.B1(n_1257),
.B2(n_1253),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1245),
.A2(n_1207),
.B(n_1256),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1245),
.A2(n_1207),
.B(n_1256),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1250),
.B(n_1280),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1151),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1179),
.B(n_1156),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1151),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1156),
.A2(n_1277),
.B(n_1271),
.Y(n_1387)
);

AO21x1_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_1123),
.B(n_1117),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1151),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1210),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1179),
.B(n_1156),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1255),
.A2(n_1288),
.B(n_1284),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1164),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1254),
.A2(n_1285),
.A3(n_1277),
.B(n_1263),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1179),
.B(n_1156),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1179),
.B(n_1156),
.Y(n_1396)
);

INVx8_ASAP7_75t_L g1397 ( 
.A(n_1164),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1247),
.B(n_1206),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1213),
.Y(n_1399)
);

BUFx8_ASAP7_75t_L g1400 ( 
.A(n_1151),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1210),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1254),
.A2(n_1030),
.B(n_1087),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1249),
.A2(n_1273),
.B(n_1271),
.C(n_1254),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1247),
.B(n_1206),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1150),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1176),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1254),
.A2(n_1285),
.A3(n_1277),
.B(n_1263),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1179),
.B(n_1156),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1209),
.B(n_1087),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1255),
.A2(n_1288),
.B(n_1284),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1303),
.B(n_1383),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1347),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1339),
.B(n_1331),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1331),
.B(n_1356),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1335),
.B(n_1393),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1289),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1333),
.B(n_1298),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1320),
.A2(n_1409),
.B1(n_1343),
.B2(n_1333),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1388),
.A2(n_1313),
.B(n_1387),
.C(n_1290),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1296),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1314),
.B(n_1365),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1336),
.B(n_1326),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1364),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1336),
.B(n_1326),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1290),
.A2(n_1367),
.B(n_1387),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1380),
.A2(n_1292),
.B(n_1299),
.C(n_1316),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1299),
.B(n_1316),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1300),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1314),
.B(n_1365),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1344),
.A2(n_1378),
.B1(n_1327),
.B2(n_1330),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1366),
.B(n_1379),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1390),
.B(n_1401),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1334),
.B(n_1349),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1334),
.B(n_1399),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1344),
.A2(n_1378),
.B1(n_1389),
.B2(n_1353),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1402),
.A2(n_1403),
.B(n_1371),
.C(n_1372),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1301),
.A2(n_1371),
.B1(n_1403),
.B2(n_1322),
.C(n_1311),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1375),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1341),
.A2(n_1317),
.B(n_1361),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1373),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1442)
);

AOI21x1_ASAP7_75t_SL g1443 ( 
.A1(n_1385),
.A2(n_1396),
.B(n_1408),
.Y(n_1443)
);

O2A1O1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1322),
.A2(n_1399),
.B(n_1408),
.C(n_1395),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1353),
.A2(n_1355),
.B1(n_1386),
.B2(n_1384),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1352),
.B(n_1391),
.C(n_1396),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1335),
.A2(n_1354),
.B(n_1410),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1385),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1308),
.A2(n_1350),
.B1(n_1351),
.B2(n_1311),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1391),
.B(n_1395),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1310),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1400),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1364),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1340),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1354),
.A2(n_1410),
.B(n_1392),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1332),
.B(n_1323),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1309),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1341),
.A2(n_1295),
.B(n_1305),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1352),
.A2(n_1358),
.B(n_1337),
.C(n_1345),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1291),
.A2(n_1293),
.B(n_1338),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1332),
.B(n_1368),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1302),
.A2(n_1404),
.B(n_1398),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1369),
.B(n_1374),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1376),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1306),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1360),
.A2(n_1362),
.B(n_1297),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1321),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1405),
.B(n_1318),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1397),
.A2(n_1357),
.B1(n_1304),
.B2(n_1321),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1315),
.B(n_1406),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1397),
.A2(n_1346),
.B1(n_1375),
.B2(n_1406),
.Y(n_1471)
);

CKINVDCx12_ASAP7_75t_R g1472 ( 
.A(n_1324),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1315),
.B(n_1407),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1315),
.B(n_1407),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1370),
.B(n_1394),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1370),
.B(n_1394),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1358),
.A2(n_1359),
.B(n_1324),
.C(n_1363),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1370),
.B(n_1407),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1400),
.B(n_1407),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1342),
.B(n_1328),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1307),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1312),
.A2(n_1394),
.B1(n_1377),
.B2(n_1348),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1381),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1382),
.B(n_1377),
.Y(n_1484)
);

INVx4_ASAP7_75t_SL g1485 ( 
.A(n_1348),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1320),
.A2(n_1279),
.B1(n_1331),
.B2(n_898),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1393),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1364),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1316),
.A2(n_1087),
.B(n_1378),
.Y(n_1489)
);

O2A1O1Ixp5_ASAP7_75t_L g1490 ( 
.A1(n_1388),
.A2(n_1254),
.B(n_1313),
.C(n_1387),
.Y(n_1490)
);

AOI221x1_ASAP7_75t_SL g1491 ( 
.A1(n_1292),
.A2(n_557),
.B1(n_599),
.B2(n_572),
.C(n_1331),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1320),
.A2(n_1279),
.B1(n_1331),
.B2(n_898),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1303),
.B(n_1383),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1290),
.A2(n_1367),
.B(n_1387),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1335),
.B(n_1393),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1303),
.B(n_1383),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1319),
.B(n_1201),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1290),
.A2(n_1367),
.B(n_1387),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1335),
.B(n_1393),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1298),
.B(n_1314),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1289),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1298),
.B(n_1314),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1347),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1456),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1461),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1468),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1448),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1448),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1457),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1485),
.B(n_1476),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1457),
.Y(n_1514)
);

INVx5_ASAP7_75t_L g1515 ( 
.A(n_1480),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1485),
.B(n_1478),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1450),
.B(n_1434),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1420),
.A2(n_1490),
.B(n_1438),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1447),
.B(n_1455),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1484),
.B(n_1440),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1414),
.B(n_1411),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1440),
.B(n_1473),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1440),
.B(n_1474),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1424),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1460),
.B(n_1489),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1483),
.A2(n_1428),
.B(n_1479),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1416),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1418),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1435),
.B(n_1446),
.Y(n_1529)
);

INVx4_ASAP7_75t_SL g1530 ( 
.A(n_1415),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1444),
.B(n_1417),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_SL g1532 ( 
.A(n_1449),
.B(n_1436),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1421),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1422),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1427),
.B(n_1429),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1486),
.A2(n_1492),
.B1(n_1419),
.B2(n_1431),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1451),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1453),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1464),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1453),
.B(n_1488),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1463),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1430),
.B(n_1500),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1437),
.A2(n_1466),
.B(n_1471),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1426),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1494),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1502),
.B(n_1498),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1432),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1458),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1433),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1529),
.B(n_1413),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1511),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1548),
.B(n_1445),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1548),
.B(n_1493),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1496),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.B(n_1523),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1536),
.A2(n_1462),
.B(n_1499),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1540),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1499),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.B(n_1520),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1520),
.B(n_1442),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1510),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1544),
.B(n_1487),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1507),
.B(n_1487),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1467),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1507),
.B(n_1443),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1506),
.B(n_1512),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1504),
.B(n_1470),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1526),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1542),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1542),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1513),
.B(n_1472),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_SL g1579 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1515),
.B(n_1465),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1571),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1569),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1561),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1519),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1544),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1572),
.B(n_1545),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1568),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1566),
.A2(n_1536),
.B1(n_1540),
.B2(n_1545),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1580),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1566),
.A2(n_1531),
.B1(n_1513),
.B2(n_1572),
.C(n_1535),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1554),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1576),
.Y(n_1594)
);

AOI211xp5_ASAP7_75t_L g1595 ( 
.A1(n_1560),
.A2(n_1531),
.B(n_1535),
.C(n_1517),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1554),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1556),
.A2(n_1517),
.B1(n_1521),
.B2(n_1543),
.C(n_1505),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1556),
.B(n_1540),
.C(n_1518),
.Y(n_1599)
);

OAI31xp33_ASAP7_75t_L g1600 ( 
.A1(n_1556),
.A2(n_1532),
.A3(n_1509),
.B(n_1508),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1452),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1575),
.A2(n_1543),
.B1(n_1505),
.B2(n_1504),
.C(n_1549),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1576),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

AO31x2_ASAP7_75t_L g1605 ( 
.A1(n_1562),
.A2(n_1546),
.A3(n_1547),
.B(n_1550),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1607)
);

AOI21xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1560),
.A2(n_1454),
.B(n_1439),
.Y(n_1608)
);

OAI33xp33_ASAP7_75t_L g1609 ( 
.A1(n_1574),
.A2(n_1528),
.A3(n_1527),
.B1(n_1533),
.B2(n_1537),
.B3(n_1539),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1571),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1562),
.A2(n_1540),
.B1(n_1545),
.B2(n_1525),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1512),
.Y(n_1612)
);

OAI211xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1574),
.A2(n_1549),
.B(n_1551),
.C(n_1528),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1561),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1577),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1557),
.A2(n_1540),
.B(n_1525),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1562),
.A2(n_1540),
.B1(n_1525),
.B2(n_1518),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.B(n_1516),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1570),
.A2(n_1551),
.B1(n_1508),
.B2(n_1509),
.C(n_1527),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1564),
.A2(n_1525),
.B1(n_1518),
.B2(n_1519),
.C(n_1497),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1581),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1606),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1594),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1557),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1606),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1603),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1616),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1588),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_L g1633 ( 
.A(n_1599),
.B(n_1518),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1584),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1605),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1619),
.Y(n_1637)
);

INVx4_ASAP7_75t_SL g1638 ( 
.A(n_1585),
.Y(n_1638)
);

AND4x1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1579),
.C(n_1532),
.D(n_1439),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1595),
.B(n_1553),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1593),
.B(n_1567),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1607),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1553),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1581),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1585),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1615),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1625),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_R g1650 ( 
.A(n_1626),
.B(n_1412),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1644),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1633),
.B(n_1589),
.C(n_1600),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1634),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1646),
.B(n_1610),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1610),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1619),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1644),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1640),
.A2(n_1617),
.B1(n_1525),
.B2(n_1545),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1638),
.B(n_1644),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1627),
.B(n_1598),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.Y(n_1663)
);

OAI33xp33_ASAP7_75t_L g1664 ( 
.A1(n_1627),
.A2(n_1607),
.A3(n_1593),
.B1(n_1604),
.B2(n_1618),
.B3(n_1613),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1626),
.B(n_1587),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1604),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1641),
.B(n_1591),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1648),
.B(n_1596),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1625),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1644),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1634),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1640),
.A2(n_1609),
.B1(n_1608),
.B2(n_1622),
.C(n_1621),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1629),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1631),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1623),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1623),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1582),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1648),
.B(n_1642),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1612),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1631),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1644),
.B(n_1614),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1679),
.B(n_1645),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1649),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1679),
.B(n_1633),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1624),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1680),
.B(n_1633),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1661),
.B(n_1624),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1680),
.B(n_1636),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1650),
.A2(n_1601),
.B(n_1624),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1676),
.B(n_1636),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1661),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1652),
.A2(n_1611),
.B1(n_1628),
.B2(n_1647),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1669),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1628),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1656),
.B(n_1628),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1665),
.B(n_1636),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1654),
.B(n_1643),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1668),
.B(n_1642),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1656),
.B(n_1638),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1670),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1653),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1651),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1683),
.B(n_1638),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1668),
.B(n_1642),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1683),
.B(n_1638),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1682),
.B(n_1632),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1643),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1663),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1670),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1643),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1652),
.A2(n_1525),
.B1(n_1585),
.B2(n_1647),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1662),
.A2(n_1647),
.B1(n_1630),
.B2(n_1518),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1682),
.B(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1671),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1687),
.Y(n_1722)
);

NOR2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1630),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1708),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1707),
.B(n_1452),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1696),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1728)
);

BUFx2_ASAP7_75t_SL g1729 ( 
.A(n_1696),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1718),
.A2(n_1664),
.B1(n_1658),
.B2(n_1647),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1708),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1651),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1700),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1693),
.B(n_1674),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

CKINVDCx16_ASAP7_75t_R g1736 ( 
.A(n_1705),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1711),
.B(n_1651),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1687),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1704),
.B(n_1662),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1694),
.A2(n_1579),
.B(n_1441),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1666),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1710),
.B(n_1666),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1710),
.B(n_1667),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1717),
.B(n_1671),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1722),
.Y(n_1748)
);

OAI31xp33_ASAP7_75t_SL g1749 ( 
.A1(n_1723),
.A2(n_1719),
.A3(n_1705),
.B(n_1690),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1730),
.A2(n_1697),
.B1(n_1699),
.B2(n_1690),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1734),
.B(n_1713),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1726),
.B(n_1728),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1729),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1726),
.B(n_1692),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1738),
.Y(n_1756)
);

AOI221x1_ASAP7_75t_L g1757 ( 
.A1(n_1739),
.A2(n_1691),
.B1(n_1688),
.B2(n_1716),
.C(n_1706),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1733),
.B(n_1721),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1733),
.B(n_1701),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1725),
.Y(n_1760)
);

AOI221x1_ASAP7_75t_L g1761 ( 
.A1(n_1739),
.A2(n_1702),
.B1(n_1716),
.B2(n_1698),
.C(n_1706),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1728),
.A2(n_1699),
.B1(n_1630),
.B2(n_1638),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1727),
.Y(n_1764)
);

AOI321xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1746),
.A2(n_1583),
.A3(n_1639),
.B1(n_1712),
.B2(n_1720),
.C(n_1702),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1735),
.A2(n_1630),
.B1(n_1638),
.B2(n_1651),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1725),
.B(n_1659),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1749),
.B(n_1754),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1753),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1764),
.B(n_1725),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1760),
.B(n_1725),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1758),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1750),
.A2(n_1741),
.B1(n_1734),
.B2(n_1744),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1755),
.B(n_1727),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1765),
.A2(n_1740),
.B1(n_1731),
.B2(n_1724),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1763),
.B(n_1732),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1745),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1762),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_SL g1781 ( 
.A(n_1773),
.B(n_1761),
.C(n_1757),
.D(n_1766),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1768),
.A2(n_1749),
.B(n_1759),
.C(n_1752),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1773),
.A2(n_1767),
.B1(n_1745),
.B2(n_1740),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1779),
.B(n_1770),
.Y(n_1784)
);

AOI332xp33_ASAP7_75t_L g1785 ( 
.A1(n_1775),
.A2(n_1756),
.A3(n_1731),
.B1(n_1698),
.B2(n_1689),
.B3(n_1737),
.C1(n_1732),
.C2(n_1715),
.Y(n_1785)
);

AO21x1_ASAP7_75t_L g1786 ( 
.A1(n_1772),
.A2(n_1737),
.B(n_1742),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1769),
.B(n_1742),
.Y(n_1787)
);

AOI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1771),
.A2(n_1743),
.B(n_1747),
.Y(n_1788)
);

XNOR2xp5_ASAP7_75t_L g1789 ( 
.A(n_1778),
.B(n_1639),
.Y(n_1789)
);

OAI21xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1781),
.A2(n_1775),
.B(n_1776),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1782),
.A2(n_1777),
.B1(n_1774),
.B2(n_1780),
.C(n_1747),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1783),
.A2(n_1743),
.B(n_1720),
.C(n_1712),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1787),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1784),
.A2(n_1638),
.B1(n_1657),
.B2(n_1672),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1793),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1790),
.B(n_1788),
.C(n_1785),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1791),
.B(n_1786),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1794),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1792),
.B(n_1789),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1793),
.B(n_1659),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1796),
.B(n_1660),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1800),
.B(n_1657),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1795),
.B(n_1441),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1799),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1798),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1805),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1801),
.B(n_1412),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1804),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1806),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1809),
.B(n_1807),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1808),
.B(n_1802),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1810),
.Y(n_1812)
);

OAI22x1_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1812),
.B1(n_1503),
.B2(n_1714),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1811),
.A2(n_1715),
.B1(n_1714),
.B2(n_1503),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1813),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1815),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_R g1817 ( 
.A1(n_1816),
.A2(n_1811),
.B1(n_1814),
.B2(n_1663),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1817),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_SL g1819 ( 
.A1(n_1818),
.A2(n_1678),
.B(n_1684),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1672),
.B1(n_1657),
.B2(n_1673),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1820),
.A2(n_1684),
.B(n_1675),
.C(n_1677),
.Y(n_1821)
);


endmodule