module fake_jpeg_20595_n_233 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_96;

INVx2_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_23),
.Y(n_59)
);

AO22x2_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_14),
.B1(n_15),
.B2(n_21),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_53),
.A3(n_22),
.B1(n_18),
.B2(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_22),
.B(n_18),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_60),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_14),
.B1(n_28),
.B2(n_17),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_66),
.B1(n_71),
.B2(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_14),
.B1(n_22),
.B2(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_14),
.B1(n_28),
.B2(n_17),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_47),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_14),
.B1(n_16),
.B2(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_24),
.B1(n_19),
.B2(n_27),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_21),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_41),
.A3(n_43),
.B1(n_47),
.B2(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_90),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_74),
.B(n_24),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_40),
.C(n_47),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_74),
.C(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_95),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_58),
.B(n_25),
.C(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_98),
.B1(n_52),
.B2(n_17),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_58),
.B1(n_40),
.B2(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_103),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_70),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_113),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_70),
.C(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_23),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_64),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_62),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_62),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_124),
.B(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_88),
.B(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_80),
.B1(n_40),
.B2(n_28),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_95),
.B(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_89),
.B1(n_91),
.B2(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_136),
.B1(n_148),
.B2(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_140),
.B(n_146),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_94),
.B1(n_105),
.B2(n_120),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_143),
.Y(n_161)
);

AOI22x1_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_90),
.B1(n_83),
.B2(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_94),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_120),
.B1(n_109),
.B2(n_121),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_147),
.B(n_136),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_156),
.B(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_167),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_115),
.B1(n_127),
.B2(n_114),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_123),
.B(n_116),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_91),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_116),
.B1(n_84),
.B2(n_100),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_116),
.B(n_84),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_100),
.C(n_107),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.C(n_163),
.Y(n_173)
);

AOI211xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_112),
.B(n_113),
.C(n_73),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_82),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_82),
.C(n_73),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_165),
.B(n_145),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_158),
.B1(n_154),
.B2(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_149),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_128),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_152),
.C(n_149),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_139),
.C(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_182),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_159),
.B(n_131),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_128),
.Y(n_177)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_135),
.C(n_131),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_194),
.B1(n_195),
.B2(n_186),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_170),
.C(n_2),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_167),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_153),
.B1(n_150),
.B2(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_195),
.B(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_176),
.B1(n_180),
.B2(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_202),
.B1(n_192),
.B2(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_170),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_1),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_5),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_190),
.C(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_5),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_190),
.B(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_205),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_218),
.B(n_219),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_197),
.C(n_6),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_211),
.C(n_6),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_13),
.B(n_7),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_207),
.B(n_206),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_220),
.B(n_8),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_5),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_7),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_228),
.C(n_229),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_8),
.C(n_10),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_223),
.C(n_231),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_13),
.Y(n_233)
);


endmodule