module fake_jpeg_1678_n_498 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_498);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_498;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_75),
.Y(n_131)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_91),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx11_ASAP7_75t_SL g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_14),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_90),
.B(n_30),
.C(n_49),
.Y(n_136)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_14),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_96),
.Y(n_149)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_102),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_31),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_107),
.B(n_140),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_109),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_30),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_132),
.B(n_136),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_24),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_146),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_53),
.B(n_24),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_31),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_38),
.B(n_20),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_54),
.B(n_23),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_38),
.Y(n_176)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_97),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_57),
.B(n_25),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_168),
.B(n_181),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_117),
.A2(n_44),
.B1(n_49),
.B2(n_40),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_170),
.A2(n_172),
.B1(n_200),
.B2(n_210),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_171),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_63),
.B1(n_99),
.B2(n_92),
.Y(n_172)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_176),
.B(n_180),
.Y(n_237)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_102),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_198),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_185),
.Y(n_245)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_28),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_202),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_119),
.A2(n_74),
.B1(n_81),
.B2(n_79),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_72),
.B1(n_71),
.B2(n_62),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_23),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_205),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_207),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_22),
.B(n_48),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_114),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_209),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_128),
.A2(n_22),
.B1(n_18),
.B2(n_48),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_76),
.B1(n_56),
.B2(n_50),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_213),
.B1(n_215),
.B2(n_22),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_143),
.A2(n_50),
.B1(n_41),
.B2(n_20),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_120),
.A2(n_18),
.B1(n_48),
.B2(n_46),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_164),
.C(n_118),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_173),
.A2(n_163),
.B1(n_158),
.B2(n_157),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_238),
.B1(n_211),
.B2(n_213),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_155),
.B1(n_134),
.B2(n_40),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_250),
.B1(n_171),
.B2(n_201),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_163),
.B1(n_158),
.B2(n_157),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_142),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_197),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_147),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_258),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_185),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_174),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_255),
.B(n_262),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_273),
.B(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_195),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_265),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_196),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_266),
.Y(n_288)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

BUFx16f_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_202),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_197),
.B1(n_206),
.B2(n_201),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_218),
.B1(n_190),
.B2(n_193),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_197),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_276),
.Y(n_308)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_214),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_214),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_246),
.Y(n_297)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_234),
.A2(n_191),
.B1(n_177),
.B2(n_209),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_245),
.B(n_230),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_283),
.B(n_265),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_240),
.B1(n_238),
.B2(n_223),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_295),
.B1(n_303),
.B2(n_274),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_302),
.B1(n_252),
.B2(n_274),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_268),
.B(n_279),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_307),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_231),
.B(n_235),
.Y(n_292)
);

XOR2x1_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_294),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_231),
.B(n_247),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_246),
.B1(n_229),
.B2(n_227),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_227),
.C(n_244),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_307),
.C(n_290),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_266),
.A2(n_189),
.B1(n_133),
.B2(n_135),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_222),
.B1(n_169),
.B2(n_121),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g305 ( 
.A1(n_257),
.A2(n_248),
.A3(n_244),
.B1(n_225),
.B2(n_28),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_248),
.B(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_313),
.B1(n_327),
.B2(n_328),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_297),
.C(n_308),
.Y(n_350)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_261),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_314),
.B(n_320),
.Y(n_357)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_284),
.B(n_277),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_272),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_322),
.Y(n_358)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_269),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_329),
.Y(n_352)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_280),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_224),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_330),
.Y(n_346)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_304),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_332),
.A2(n_333),
.B(n_265),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_224),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_334),
.Y(n_348)
);

CKINVDCx12_ASAP7_75t_R g336 ( 
.A(n_287),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_336),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_308),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_337),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g339 ( 
.A(n_323),
.B(n_287),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_339),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_323),
.A2(n_287),
.B(n_296),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_315),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_285),
.B1(n_294),
.B2(n_286),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_351),
.B1(n_361),
.B2(n_325),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_300),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_362),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_335),
.B(n_329),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_349),
.B(n_313),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_363),
.C(n_362),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_331),
.B1(n_337),
.B2(n_322),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_282),
.B(n_295),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_356),
.A2(n_364),
.B(n_332),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_318),
.A2(n_303),
.B1(n_282),
.B2(n_302),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_275),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_264),
.C(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_382),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_320),
.B1(n_314),
.B2(n_326),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_368),
.A2(n_369),
.B1(n_370),
.B2(n_375),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_360),
.A2(n_344),
.B1(n_357),
.B2(n_346),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_317),
.B1(n_310),
.B2(n_319),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_374),
.B(n_356),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_325),
.C(n_316),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_379),
.C(n_383),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_391),
.Y(n_399)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_306),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_380),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_328),
.C(n_327),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_SL g380 ( 
.A(n_364),
.B(n_291),
.C(n_153),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_340),
.B(n_291),
.CI(n_260),
.CON(n_381),
.SN(n_381)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_343),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_260),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_184),
.C(n_205),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_384),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_178),
.C(n_267),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_386),
.C(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_186),
.C(n_188),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_388),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_339),
.B(n_142),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_354),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_194),
.C(n_179),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_153),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_351),
.B(n_365),
.Y(n_394)
);

AOI21x1_ASAP7_75t_SL g415 ( 
.A1(n_394),
.A2(n_414),
.B(n_381),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_396),
.A2(n_153),
.B(n_175),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_373),
.A2(n_363),
.B(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_345),
.C(n_341),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_401),
.C(n_412),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_352),
.C(n_361),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_127),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_383),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_359),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_408),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_359),
.C(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_420),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_409),
.A2(n_389),
.B1(n_382),
.B2(n_391),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_422),
.B1(n_433),
.B2(n_397),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_372),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_406),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_390),
.B1(n_376),
.B2(n_150),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_423),
.B(n_426),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_410),
.A2(n_156),
.B1(n_141),
.B2(n_50),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_156),
.C(n_150),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_428),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_394),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_396),
.A2(n_46),
.B(n_28),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_429),
.A2(n_46),
.B(n_26),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_411),
.B1(n_403),
.B2(n_407),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_127),
.C(n_113),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_397),
.C(n_408),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_113),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_432),
.B(n_0),
.Y(n_448)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_433),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_440),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_437),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_406),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_400),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_438),
.B(n_441),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_413),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_399),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_417),
.B1(n_416),
.B2(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_448),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_415),
.A2(n_26),
.B(n_25),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_449),
.A2(n_429),
.B(n_423),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_454),
.B1(n_450),
.B2(n_4),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_426),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_455),
.A2(n_450),
.B(n_435),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_436),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_457),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_431),
.C(n_125),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_125),
.C(n_26),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_458),
.B(n_461),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_25),
.C(n_16),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_1),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_465),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_460),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_467),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_445),
.C(n_437),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_473),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_461),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_1),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_475),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_454),
.C(n_457),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_464),
.B(n_1),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_16),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_476),
.A2(n_4),
.B(n_6),
.Y(n_485)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_459),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_455),
.C(n_458),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_482),
.Y(n_486)
);

AOI21xp33_ASAP7_75t_L g489 ( 
.A1(n_483),
.A2(n_479),
.B(n_480),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_12),
.C(n_6),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_471),
.C(n_474),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_468),
.B(n_6),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_490),
.C(n_4),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_489),
.B(n_481),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_473),
.C(n_7),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_491),
.A2(n_492),
.B(n_493),
.Y(n_494)
);

AOI32xp33_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_481),
.A3(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_7),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_10),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_496),
.B(n_10),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_10),
.Y(n_498)
);


endmodule