module fake_aes_12631_n_697 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_87), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_35), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_84), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_83), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_65), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_36), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_52), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_90), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_20), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_58), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_77), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_69), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_32), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_43), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_86), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_10), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_62), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_88), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_39), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_28), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_66), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_47), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_51), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_64), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_38), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_42), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_25), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_80), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_14), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_4), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_98), .B(n_0), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_99), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_113), .B(n_0), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_102), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_93), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_112), .B(n_1), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_102), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_105), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_94), .B(n_5), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_94), .A2(n_6), .B(n_7), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_114), .B(n_6), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_119), .B(n_7), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_142), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
NAND2xp33_ASAP7_75t_L g154 ( .A(n_132), .B(n_104), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_132), .B(n_115), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_142), .B(n_93), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_134), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_144), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_135), .B(n_115), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_142), .A2(n_129), .B1(n_128), .B2(n_93), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_135), .B(n_93), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_144), .A2(n_96), .B1(n_126), .B2(n_97), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_139), .B(n_101), .Y(n_166) );
BUFx10_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_134), .B(n_104), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_139), .B(n_103), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_133), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
BUFx6f_ASAP7_75t_SL g174 ( .A(n_134), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_130), .B(n_109), .Y(n_177) );
OAI22xp33_ASAP7_75t_SL g178 ( .A1(n_140), .A2(n_127), .B1(n_125), .B2(n_107), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_162), .B(n_107), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_158), .B(n_138), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_174), .B(n_140), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_168), .B(n_130), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_151), .A2(n_147), .B(n_145), .C(n_138), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_158), .B(n_138), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_176), .A2(n_136), .B1(n_105), .B2(n_108), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_177), .B(n_145), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_151), .B(n_145), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_174), .A2(n_147), .B1(n_136), .B2(n_108), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_151), .B(n_147), .Y(n_192) );
NOR2x2_ASAP7_75t_L g193 ( .A(n_178), .B(n_167), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_174), .A2(n_111), .B1(n_120), .B2(n_116), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
AND2x6_ASAP7_75t_SL g196 ( .A(n_157), .B(n_118), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_154), .B(n_122), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_152), .B(n_122), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_121), .B(n_124), .C(n_137), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_152), .B(n_125), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_152), .B(n_127), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_159), .B(n_100), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_159), .B(n_106), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_110), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_162), .B(n_111), .Y(n_213) );
NOR2xp67_ASAP7_75t_L g214 ( .A(n_157), .B(n_137), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_164), .B(n_110), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_178), .A2(n_137), .B1(n_148), .B2(n_146), .Y(n_216) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_164), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_182), .B(n_166), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_182), .B(n_164), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_192), .A2(n_170), .B(n_155), .C(n_161), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_217), .A2(n_160), .B(n_150), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_188), .B(n_166), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_197), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_197), .B(n_210), .Y(n_224) );
BUFx12f_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_186), .B(n_170), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_189), .B(n_155), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_187), .B(n_163), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_185), .A2(n_160), .B(n_150), .C(n_153), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_198), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_183), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_198), .A2(n_153), .B(n_169), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_165), .B(n_161), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_184), .B(n_165), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_191), .B(n_167), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_183), .A2(n_167), .B1(n_163), .B2(n_179), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_210), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_210), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_190), .B(n_163), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_209), .A2(n_163), .B(n_173), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_183), .A2(n_163), .B1(n_137), .B2(n_175), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_216), .A2(n_137), .B(n_175), .C(n_179), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_203), .B(n_8), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_215), .B(n_175), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_190), .A2(n_216), .B(n_207), .C(n_200), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_229), .A2(n_200), .B(n_180), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_222), .B(n_191), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_249), .A2(n_202), .B(n_214), .C(n_180), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_213), .B(n_208), .C(n_206), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_220), .A2(n_205), .B(n_201), .C(n_204), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_249), .A2(n_149), .A3(n_211), .B(n_148), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_225), .B(n_194), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_218), .B1(n_226), .B2(n_236), .C(n_247), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_219), .B(n_207), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_219), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_219), .A2(n_215), .B1(n_195), .B2(n_212), .Y(n_260) );
AOI21xp5_ASAP7_75t_SL g261 ( .A1(n_244), .A2(n_215), .B(n_181), .Y(n_261) );
AO22x1_ASAP7_75t_L g262 ( .A1(n_246), .A2(n_193), .B1(n_215), .B2(n_199), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_246), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_233), .A2(n_214), .B(n_212), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_239), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_228), .B(n_212), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_221), .A2(n_173), .B(n_172), .Y(n_268) );
NOR2xp67_ASAP7_75t_SL g269 ( .A(n_225), .B(n_123), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_175), .B(n_179), .C(n_149), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_259), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_232), .B1(n_243), .B2(n_246), .C(n_241), .Y(n_273) );
INVx6_ASAP7_75t_L g274 ( .A(n_259), .Y(n_274) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_270), .A2(n_234), .B(n_149), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_263), .B(n_230), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_271), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_251), .B(n_224), .Y(n_280) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_252), .A2(n_149), .B(n_242), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
CKINVDCx6p67_ASAP7_75t_R g284 ( .A(n_269), .Y(n_284) );
BUFx12f_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_260), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_254), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_255), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_253), .A2(n_245), .B(n_230), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_250), .A2(n_245), .B(n_248), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_266), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_265), .A2(n_248), .B(n_237), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_279), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
AOI21x1_ASAP7_75t_L g297 ( .A1(n_289), .A2(n_262), .B(n_260), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_289), .A2(n_261), .B(n_268), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_287), .B(n_278), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_287), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_282), .B(n_255), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_291), .A2(n_267), .B(n_146), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_282), .B(n_256), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_276), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_291), .A2(n_276), .B(n_288), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_238), .Y(n_309) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_292), .B(n_231), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_283), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_290), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_281), .A2(n_146), .B(n_148), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_273), .B(n_231), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_286), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_277), .B(n_224), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_277), .B(n_239), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_273), .B(n_123), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_296), .B(n_319), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_306), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_320), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_296), .B(n_272), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_303), .B(n_292), .Y(n_333) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_319), .B(n_284), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_319), .B(n_275), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_275), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_305), .B(n_292), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_307), .Y(n_338) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_297), .A2(n_293), .B(n_275), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
NOR2x1_ASAP7_75t_SL g341 ( .A(n_311), .B(n_285), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_295), .B(n_275), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_295), .B(n_272), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_295), .B(n_280), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_301), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_299), .B(n_275), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_311), .B(n_274), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_294), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_294), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_300), .B(n_274), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_299), .B(n_293), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_307), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_300), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_299), .B(n_9), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_302), .A2(n_284), .B(n_143), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_308), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_324), .B(n_123), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_308), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_305), .B(n_285), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_308), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_304), .B(n_117), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_309), .B(n_274), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_312), .B(n_9), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_304), .B(n_117), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_304), .B(n_274), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_304), .B(n_317), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_323), .B(n_143), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_323), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_328), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_328), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_340), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_347), .B(n_323), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_347), .B(n_316), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_372), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_326), .B(n_313), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
INVx4_ASAP7_75t_L g391 ( .A(n_338), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_348), .B(n_316), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_348), .B(n_316), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_335), .B(n_298), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_372), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_335), .B(n_298), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_327), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_327), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_298), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_326), .B(n_313), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_357), .B(n_298), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_353), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_338), .Y(n_404) );
AND2x4_ASAP7_75t_SL g405 ( .A(n_333), .B(n_325), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_358), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_333), .B(n_325), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_327), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_349), .B(n_322), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g413 ( .A(n_361), .B(n_322), .C(n_318), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_349), .B(n_318), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_360), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_367), .B(n_309), .C(n_320), .D(n_321), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_333), .B(n_297), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_345), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_361), .B(n_309), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_333), .B(n_143), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_336), .B(n_143), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_329), .B(n_321), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_354), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_371), .B(n_321), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_377), .B(n_320), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_371), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_375), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_336), .B(n_143), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_331), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_345), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_342), .B(n_143), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_342), .B(n_143), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_362), .B(n_346), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_346), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_365), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_362), .B(n_365), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_378), .B(n_10), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_373), .B(n_274), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_374), .Y(n_445) );
NOR2x1_ASAP7_75t_L g446 ( .A(n_363), .B(n_284), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_378), .B(n_11), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_330), .B(n_310), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_330), .B(n_310), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_380), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_356), .B(n_310), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_331), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_377), .B(n_11), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_370), .B(n_12), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_344), .B(n_13), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_370), .B(n_13), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_332), .B(n_14), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_332), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_401), .B(n_403), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_389), .B(n_351), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_446), .A2(n_341), .B(n_334), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_438), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_334), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_427), .B(n_334), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_401), .B(n_368), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_391), .B(n_440), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_427), .B(n_376), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_389), .B(n_351), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_400), .B(n_352), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_427), .B(n_376), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_410), .B(n_379), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_408), .B(n_368), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_410), .B(n_344), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_408), .B(n_369), .Y(n_476) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_446), .B(n_337), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_409), .B(n_369), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_391), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_454), .B(n_343), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_391), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_400), .B(n_359), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_416), .A2(n_350), .B1(n_285), .B2(n_343), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_359), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_454), .B(n_352), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_416), .A2(n_364), .B(n_341), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_391), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_415), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_431), .B(n_364), .Y(n_490) );
OAI332xp33_ASAP7_75t_L g491 ( .A1(n_419), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_339), .C1(n_364), .C2(n_156), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_431), .B(n_364), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_418), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_418), .Y(n_494) );
OR2x6_ASAP7_75t_L g495 ( .A(n_440), .B(n_339), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_440), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_433), .B(n_339), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_456), .B(n_15), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_439), .B(n_16), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_406), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_439), .Y(n_503) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_443), .B(n_17), .Y(n_504) );
INVx3_ASAP7_75t_SL g505 ( .A(n_440), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_381), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_429), .B(n_18), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_405), .B(n_19), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_381), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_433), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_382), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_413), .A2(n_156), .B(n_179), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_443), .B(n_26), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_382), .B(n_27), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_383), .Y(n_515) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_404), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_385), .B(n_29), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_425), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_385), .B(n_30), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_399), .A2(n_156), .B1(n_172), .B2(n_171), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_428), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_414), .B(n_31), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_447), .B(n_33), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_445), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_426), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_447), .B(n_34), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_430), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_441), .B(n_40), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_405), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_394), .B(n_41), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_451), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_394), .B(n_44), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_451), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_428), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_396), .B(n_45), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_442), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_414), .B(n_48), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_399), .B(n_50), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_425), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_450), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_402), .B(n_384), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_542), .B(n_412), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_481), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_462), .A2(n_457), .B(n_455), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_475), .B(n_402), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_504), .A2(n_457), .B(n_455), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_525), .B(n_450), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_468), .B(n_458), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_527), .B(n_444), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_469), .B(n_405), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_530), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_472), .B(n_421), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_473), .B(n_421), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_463), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_487), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_468), .B(n_458), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_537), .B(n_423), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_502), .B(n_384), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_466), .B(n_420), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_466), .B(n_420), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_474), .B(n_420), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_521), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_474), .B(n_407), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_480), .B(n_417), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_484), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_496), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_476), .B(n_407), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_461), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_470), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_476), .B(n_407), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_486), .B(n_490), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_486), .B(n_417), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g576 ( .A(n_483), .B(n_449), .C(n_448), .D(n_452), .Y(n_576) );
NOR2xp67_ASAP7_75t_L g577 ( .A(n_510), .B(n_395), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_488), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_478), .B(n_390), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_478), .B(n_390), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_471), .B(n_395), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_482), .B(n_388), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_485), .B(n_388), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_477), .B(n_437), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_505), .B(n_387), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_494), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_508), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_492), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_540), .B(n_387), .Y(n_592) );
NOR2xp33_ASAP7_75t_SL g593 ( .A(n_508), .B(n_437), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_541), .B(n_390), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_479), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_464), .B(n_436), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_465), .B(n_436), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_497), .B(n_432), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_518), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_528), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_532), .B(n_432), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_534), .B(n_422), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_499), .B(n_422), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_510), .A2(n_386), .B1(n_392), .B2(n_393), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_498), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_503), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_506), .B(n_453), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_509), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_511), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_582), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_547), .B(n_515), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_548), .A2(n_507), .B1(n_495), .B2(n_500), .C(n_538), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_600), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_586), .B(n_495), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_545), .A2(n_539), .B1(n_522), .B2(n_538), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_564), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_569), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_565), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_556), .B(n_501), .Y(n_619) );
OAI322xp33_ASAP7_75t_L g620 ( .A1(n_543), .A2(n_522), .A3(n_501), .B1(n_539), .B2(n_519), .C1(n_514), .C2(n_517), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_593), .A2(n_491), .B(n_513), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_588), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_548), .A2(n_523), .B(n_526), .Y(n_623) );
NOR3xp33_ASAP7_75t_SL g624 ( .A(n_576), .B(n_491), .C(n_514), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_546), .B(n_536), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_591), .B(n_567), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_577), .A2(n_529), .B(n_533), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_571), .B(n_434), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_578), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_531), .B(n_386), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_553), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_585), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_575), .A2(n_392), .B1(n_393), .B2(n_517), .C1(n_519), .C2(n_520), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_575), .A2(n_453), .B1(n_459), .B2(n_434), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_603), .B(n_459), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_552), .B(n_459), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_604), .A2(n_512), .B(n_434), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_549), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_561), .B(n_411), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_568), .B(n_411), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_574), .B(n_398), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_594), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_574), .B(n_398), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g645 ( .A1(n_590), .A2(n_397), .A3(n_54), .B1(n_55), .B2(n_56), .Y(n_645) );
AOI321xp33_ASAP7_75t_L g646 ( .A1(n_621), .A2(n_550), .A3(n_558), .B1(n_551), .B2(n_602), .C(n_598), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_623), .A2(n_560), .B1(n_559), .B2(n_544), .Y(n_647) );
OAI222xp33_ASAP7_75t_L g648 ( .A1(n_612), .A2(n_557), .B1(n_554), .B2(n_596), .C1(n_597), .C2(n_555), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_610), .B(n_609), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_623), .A2(n_602), .B1(n_595), .B2(n_572), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_631), .A2(n_601), .B1(n_584), .B2(n_583), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_615), .A2(n_589), .B(n_606), .C(n_605), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_611), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_618), .Y(n_654) );
OAI221xp5_ASAP7_75t_SL g655 ( .A1(n_630), .A2(n_581), .B1(n_562), .B2(n_563), .C(n_566), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_624), .A2(n_608), .B1(n_579), .B2(n_573), .C(n_563), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_627), .A2(n_579), .B1(n_566), .B2(n_580), .Y(n_657) );
AOI322xp5_ASAP7_75t_L g658 ( .A1(n_617), .A2(n_580), .A3(n_570), .B1(n_599), .B2(n_397), .C1(n_607), .C2(n_592), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_639), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_613), .B(n_570), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g661 ( .A(n_614), .B(n_53), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_616), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_627), .A2(n_171), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_663) );
AOI321xp33_ASAP7_75t_L g664 ( .A1(n_614), .A2(n_619), .A3(n_644), .B1(n_622), .B2(n_626), .C(n_642), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_633), .B(n_57), .Y(n_665) );
NOR2xp33_ASAP7_75t_SL g666 ( .A(n_637), .B(n_63), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_634), .B(n_67), .C(n_68), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_644), .A2(n_71), .B(n_72), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_640), .A2(n_73), .B(n_74), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_625), .A2(n_75), .B1(n_76), .B2(n_78), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_629), .A2(n_79), .B1(n_81), .B2(n_82), .C1(n_85), .C2(n_632), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_645), .A2(n_638), .B(n_641), .C(n_628), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_643), .A2(n_635), .B(n_636), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_620), .B(n_621), .C(n_612), .D(n_548), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_614), .B(n_623), .Y(n_675) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_664), .B(n_646), .C(n_656), .Y(n_676) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_674), .B(n_665), .C(n_656), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_654), .A2(n_675), .B(n_652), .C(n_658), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_672), .B(n_663), .C(n_648), .Y(n_679) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_667), .B(n_650), .Y(n_680) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_647), .B(n_659), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_681), .B(n_653), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_661), .B(n_666), .C(n_668), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_678), .Y(n_684) );
NOR2xp67_ASAP7_75t_SL g685 ( .A(n_680), .B(n_669), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_684), .B(n_676), .C(n_679), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_682), .Y(n_687) );
NOR4xp25_ASAP7_75t_L g688 ( .A(n_683), .B(n_655), .C(n_657), .D(n_649), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_687), .B(n_685), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_686), .Y(n_690) );
AOI21xp33_ASAP7_75t_SL g691 ( .A1(n_690), .A2(n_688), .B(n_683), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_689), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_692), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_693), .Y(n_694) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_694), .A2(n_691), .B(n_671), .Y(n_695) );
OA22x2_ASAP7_75t_L g696 ( .A1(n_695), .A2(n_670), .B1(n_673), .B2(n_662), .Y(n_696) );
AOI21xp33_ASAP7_75t_SL g697 ( .A1(n_696), .A2(n_651), .B(n_660), .Y(n_697) );
endmodule