module fake_jpeg_24629_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_8),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_30),
.B1(n_28),
.B2(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_67),
.B1(n_74),
.B2(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_16),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_40),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_83),
.B1(n_31),
.B2(n_29),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_88),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_16),
.B1(n_20),
.B2(n_33),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_108),
.B1(n_110),
.B2(n_54),
.Y(n_136)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_25),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

OA22x2_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_34),
.B1(n_17),
.B2(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_54),
.A2(n_40),
.B1(n_49),
.B2(n_34),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_119),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_63),
.A2(n_23),
.B1(n_33),
.B2(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_27),
.B1(n_29),
.B2(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_73),
.Y(n_143)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_66),
.B1(n_58),
.B2(n_27),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_62),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_105),
.B1(n_100),
.B2(n_96),
.Y(n_159)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_139),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_108),
.B1(n_94),
.B2(n_92),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_119),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_153),
.C(n_2),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_9),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_86),
.B(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_1),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_88),
.B(n_27),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_159),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_184),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_108),
.B1(n_100),
.B2(n_112),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_118),
.B1(n_92),
.B2(n_107),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_93),
.B1(n_99),
.B2(n_104),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_171),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_110),
.B1(n_111),
.B2(n_90),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_169),
.B1(n_185),
.B2(n_152),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_91),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_110),
.B1(n_116),
.B2(n_103),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_110),
.B(n_85),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_141),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_182),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_111),
.B(n_19),
.C(n_109),
.Y(n_175)
);

XOR2x1_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_138),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_122),
.B(n_85),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_177),
.B1(n_186),
.B2(n_150),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_138),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_123),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_149),
.B1(n_139),
.B2(n_153),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_3),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_190),
.B(n_203),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_206),
.B(n_219),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_132),
.B1(n_153),
.B2(n_130),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_218),
.B1(n_176),
.B2(n_173),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_153),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_6),
.B(n_7),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_135),
.B1(n_128),
.B2(n_126),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_196),
.A2(n_201),
.B1(n_176),
.B2(n_167),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_210),
.Y(n_235)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_135),
.B1(n_128),
.B2(n_126),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_212),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_145),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_166),
.C(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_221),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_187),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_157),
.CI(n_179),
.CON(n_226),
.SN(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_160),
.A2(n_152),
.B1(n_125),
.B2(n_6),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_4),
.B(n_5),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_5),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_185),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_157),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_225),
.B(n_241),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_181),
.B(n_160),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_232),
.B1(n_247),
.B2(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_245),
.C(n_197),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_167),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_244),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_219),
.B1(n_201),
.B2(n_195),
.Y(n_260)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_6),
.A3(n_7),
.B1(n_13),
.B2(n_14),
.C1(n_176),
.C2(n_217),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_242),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_13),
.C(n_14),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_194),
.B(n_191),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_210),
.Y(n_250)
);

OAI31xp33_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_235),
.A3(n_224),
.B(n_226),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_259),
.C(n_261),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_192),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_266),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_205),
.B1(n_203),
.B2(n_190),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_258),
.B1(n_272),
.B2(n_242),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_200),
.B1(n_207),
.B2(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_192),
.C(n_196),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_262),
.B1(n_265),
.B2(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_211),
.C(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_227),
.B1(n_230),
.B2(n_237),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_237),
.B1(n_236),
.B2(n_248),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_223),
.A2(n_225),
.B1(n_238),
.B2(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_224),
.A2(n_244),
.B1(n_231),
.B2(n_240),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_235),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_285),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_233),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_258),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_281),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_224),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_226),
.C(n_245),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_289),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_292),
.B(n_252),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_296),
.B(n_284),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_268),
.B(n_229),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_262),
.B1(n_260),
.B2(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_257),
.B1(n_229),
.B2(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_272),
.B1(n_254),
.B2(n_266),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_307),
.B1(n_241),
.B2(n_280),
.Y(n_314)
);

BUFx12_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_234),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_275),
.A2(n_268),
.B1(n_251),
.B2(n_234),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_311),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_292),
.B(n_286),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_287),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_274),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_280),
.C(n_285),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_320),
.B1(n_301),
.B2(n_300),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_274),
.C(n_276),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_255),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_318),
.B(n_294),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_327),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_326),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_315),
.C(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_301),
.C(n_312),
.Y(n_332)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_277),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_319),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_332),
.A2(n_333),
.B(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_305),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_328),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_309),
.C(n_295),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_325),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_306),
.B(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_329),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_341),
.A2(n_340),
.B(n_337),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_342),
.C(n_331),
.Y(n_345)
);

XNOR2x2_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_330),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_323),
.C(n_293),
.Y(n_347)
);


endmodule