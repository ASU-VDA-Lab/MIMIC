module fake_jpeg_3757_n_296 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_34),
.B(n_24),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_24),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_17),
.B1(n_29),
.B2(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_54),
.Y(n_77)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_62),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_23),
.B1(n_33),
.B2(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_17),
.B1(n_44),
.B2(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_32),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_33),
.B(n_23),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_94),
.C(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_55),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_103),
.B(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_59),
.B(n_45),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_109),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_93),
.C(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_53),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_117),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_36),
.B1(n_43),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_81),
.B1(n_80),
.B2(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.Y(n_150)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_28),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_62),
.C(n_66),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_23),
.C(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_96),
.B1(n_31),
.B2(n_28),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_78),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_143),
.B1(n_80),
.B2(n_74),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_88),
.B1(n_43),
.B2(n_36),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_70),
.B1(n_65),
.B2(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2x1p5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_36),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_42),
.B1(n_35),
.B2(n_43),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_69),
.B(n_79),
.C(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_120),
.B(n_100),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_104),
.B(n_98),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_96),
.B1(n_69),
.B2(n_43),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_44),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_110),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_172),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_155),
.B(n_168),
.Y(n_199)
);

NAND2x1_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_127),
.C(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_177),
.C(n_129),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_106),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_173),
.B1(n_92),
.B2(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_167),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_89),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_86),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_176),
.B(n_20),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_79),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_84),
.C(n_74),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_57),
.B(n_89),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_179),
.B1(n_136),
.B2(n_44),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_57),
.B(n_42),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_140),
.C(n_129),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_172),
.C(n_199),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_188),
.C(n_193),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_135),
.C(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_125),
.B1(n_146),
.B2(n_145),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_192),
.B1(n_200),
.B2(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_195),
.B1(n_205),
.B2(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_162),
.B1(n_163),
.B2(n_152),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_147),
.B1(n_43),
.B2(n_72),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_126),
.C(n_42),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_72),
.B1(n_44),
.B2(n_42),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_42),
.C(n_35),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_168),
.C(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_128),
.B1(n_22),
.B2(n_20),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_18),
.C(n_16),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_168),
.C(n_16),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_1),
.C(n_2),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_212),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_202),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_217),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_224),
.B1(n_227),
.B2(n_21),
.Y(n_237)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_225),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_167),
.B1(n_151),
.B2(n_166),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_180),
.A2(n_18),
.B(n_34),
.Y(n_226)
);

AOI31xp67_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_201),
.A3(n_199),
.B(n_196),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_26),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_18),
.B(n_34),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_209),
.B(n_217),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_193),
.B(n_187),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_236),
.B(n_216),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_8),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_194),
.B(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_212),
.C(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_255),
.C(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

OAI221xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_247),
.B1(n_231),
.B2(n_245),
.C(n_243),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_221),
.B1(n_210),
.B2(n_214),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_261),
.B1(n_231),
.B2(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_234),
.C(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_7),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_260),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_8),
.C(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_259),
.B1(n_266),
.B2(n_252),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_10),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_261),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_232),
.B(n_241),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_251),
.B(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.C(n_257),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_12),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_240),
.C(n_238),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_10),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_272),
.B(n_13),
.C(n_14),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_276),
.B(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_279),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_253),
.B(n_248),
.Y(n_277)
);

AOI21x1_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_13),
.B(n_14),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_12),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_12),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_284),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_286),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_14),
.C(n_285),
.Y(n_292)
);

AOI21x1_ASAP7_75t_SL g293 ( 
.A1(n_292),
.A2(n_291),
.B(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_294),
.Y(n_296)
);


endmodule