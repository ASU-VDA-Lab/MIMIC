module fake_netlist_1_4796_n_591 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_591);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_591;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_56), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_1), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_3), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_45), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_43), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_6), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_48), .Y(n_93) );
NOR2xp67_ASAP7_75t_L g94 ( .A(n_1), .B(n_39), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_40), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_74), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_73), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_80), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_63), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_54), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_9), .Y(n_106) );
BUFx8_ASAP7_75t_SL g107 ( .A(n_29), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_81), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_79), .B(n_34), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_46), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_31), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_10), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_47), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_68), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_61), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
OR2x6_ASAP7_75t_L g122 ( .A(n_112), .B(n_0), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_115), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_115), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_87), .B(n_30), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_87), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_112), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_120), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_111), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_84), .B(n_4), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_94), .B(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_121), .B(n_5), .Y(n_137) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_91), .A2(n_33), .B(n_76), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_120), .B(n_6), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_110), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_86), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_123), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_122), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_129), .B(n_108), .Y(n_149) );
INVx2_ASAP7_75t_SL g150 ( .A(n_122), .Y(n_150) );
NAND3xp33_ASAP7_75t_L g151 ( .A(n_127), .B(n_118), .C(n_117), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_133), .B(n_103), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_122), .A2(n_95), .B1(n_85), .B2(n_114), .Y(n_156) );
OR2x6_ASAP7_75t_L g157 ( .A(n_122), .B(n_95), .Y(n_157) );
XNOR2xp5_ASAP7_75t_SL g158 ( .A(n_144), .B(n_90), .Y(n_158) );
OAI22xp33_ASAP7_75t_SL g159 ( .A1(n_130), .A2(n_90), .B1(n_97), .B2(n_116), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_127), .B(n_88), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_146), .B(n_88), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_128), .B(n_93), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_134), .A2(n_106), .B1(n_102), .B2(n_113), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_128), .B(n_93), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_150), .B(n_146), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_170), .B(n_131), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_164), .B(n_131), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_171), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
NAND2xp33_ASAP7_75t_L g180 ( .A(n_150), .B(n_126), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_154), .B(n_135), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_163), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_149), .B(n_135), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_174), .B(n_146), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_160), .B(n_117), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_154), .B(n_141), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_174), .B(n_142), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_154), .B(n_143), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_153), .B(n_142), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_154), .B(n_143), .Y(n_193) );
AOI22xp33_ASAP7_75t_SL g194 ( .A1(n_148), .A2(n_126), .B1(n_99), .B2(n_113), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_156), .B(n_99), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_157), .B(n_139), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_157), .B(n_140), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_162), .A2(n_138), .B(n_118), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_157), .B(n_140), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
OAI221xp5_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_151), .B1(n_136), .B2(n_140), .C(n_124), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_159), .B(n_124), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_162), .B(n_136), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_167), .B(n_124), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_160), .A2(n_82), .B(n_100), .C(n_101), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_169), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_167), .B(n_98), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_186), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_183), .A2(n_160), .B(n_105), .C(n_104), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_179), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_210), .A2(n_172), .B1(n_167), .B2(n_158), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_186), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_180), .A2(n_167), .B(n_172), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_172), .B1(n_143), .B2(n_145), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_206), .A2(n_172), .B1(n_143), .B2(n_145), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_186), .B(n_119), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_181), .A2(n_138), .B(n_168), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_190), .B(n_145), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_181), .A2(n_138), .B(n_168), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_190), .B(n_158), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_184), .B(n_145), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_182), .B(n_145), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_187), .B(n_143), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_176), .A2(n_109), .B(n_171), .C(n_173), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_189), .A2(n_138), .B(n_152), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_189), .A2(n_152), .B(n_166), .Y(n_233) );
NOR3xp33_ASAP7_75t_L g234 ( .A(n_203), .B(n_173), .C(n_166), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_191), .A2(n_193), .B(n_211), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_182), .B(n_7), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_147), .B(n_166), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_193), .A2(n_161), .B(n_155), .Y(n_238) );
NAND3xp33_ASAP7_75t_L g239 ( .A(n_194), .B(n_173), .C(n_132), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_185), .B(n_107), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_206), .A2(n_173), .B(n_161), .C(n_155), .Y(n_241) );
BUFx8_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_192), .A2(n_161), .B(n_155), .C(n_147), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_202), .B(n_132), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_196), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_201), .A2(n_132), .B1(n_125), .B2(n_123), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g247 ( .A(n_202), .B(n_147), .Y(n_247) );
BUFx8_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
OAI21xp5_ASAP7_75t_SL g249 ( .A1(n_227), .A2(n_196), .B(n_200), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_216), .Y(n_250) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_232), .A2(n_199), .B(n_209), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_218), .A2(n_208), .B(n_176), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_241), .A2(n_198), .B(n_195), .C(n_204), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_226), .A2(n_204), .B1(n_188), .B2(n_132), .Y(n_254) );
BUFx2_ASAP7_75t_SL g255 ( .A(n_236), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_132), .B(n_125), .C(n_205), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_228), .A2(n_125), .B(n_197), .C(n_178), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_245), .B(n_11), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_240), .B(n_188), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_222), .A2(n_188), .B(n_125), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_231), .A2(n_125), .B(n_188), .C(n_13), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_224), .A2(n_188), .B(n_41), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_243), .A2(n_38), .B(n_72), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_242), .B(n_11), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_42), .B(n_71), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_220), .A2(n_12), .B(n_14), .Y(n_268) );
AOI21x1_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_37), .B(n_70), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_236), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_270) );
NOR2x1_ASAP7_75t_SL g271 ( .A(n_225), .B(n_16), .Y(n_271) );
NOR3xp33_ASAP7_75t_L g272 ( .A(n_221), .B(n_17), .C(n_18), .Y(n_272) );
AND2x6_ASAP7_75t_L g273 ( .A(n_215), .B(n_19), .Y(n_273) );
BUFx10_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
AOI21x1_ASAP7_75t_SL g275 ( .A1(n_223), .A2(n_20), .B(n_22), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_212), .B(n_77), .Y(n_277) );
AO22x2_ASAP7_75t_L g278 ( .A1(n_239), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_255), .B(n_230), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_260), .A2(n_246), .B(n_220), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_266), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g282 ( .A(n_277), .B(n_217), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_249), .B(n_248), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_251), .A2(n_244), .B(n_237), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_249), .B(n_234), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_270), .A2(n_234), .B(n_229), .C(n_219), .Y(n_287) );
BUFx12f_ASAP7_75t_L g288 ( .A(n_274), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_238), .B(n_233), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_246), .B(n_247), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_263), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_65), .B(n_27), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_64), .B(n_28), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_264), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_257), .A2(n_26), .B(n_32), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_277), .B(n_44), .Y(n_297) );
AOI21x1_ASAP7_75t_L g298 ( .A1(n_278), .A2(n_267), .B(n_252), .Y(n_298) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_268), .A2(n_49), .B(n_50), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_250), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
AO21x1_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_51), .B(n_52), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_250), .B(n_53), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_297), .Y(n_304) );
AND2x4_ASAP7_75t_SL g305 ( .A(n_297), .B(n_276), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_291), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_297), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_291), .A2(n_262), .B(n_275), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_297), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_288), .Y(n_310) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_298), .A2(n_271), .B(n_272), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_297), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_278), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_298), .A2(n_254), .B(n_259), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_286), .B(n_273), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_297), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_289), .A2(n_273), .B(n_258), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_282), .B(n_273), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_295), .A2(n_273), .B(n_58), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_282), .A2(n_265), .B1(n_59), .B2(n_60), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_295), .A2(n_57), .B(n_62), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_309), .B(n_284), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_309), .A2(n_284), .B1(n_288), .B2(n_301), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_315), .A2(n_289), .B(n_295), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_322), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_313), .B(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_316), .B(n_300), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_313), .B(n_301), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_316), .B(n_294), .Y(n_338) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_321), .B(n_301), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_304), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_320), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_316), .B(n_299), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_307), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g347 ( .A1(n_319), .A2(n_302), .B(n_287), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_307), .B(n_285), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_279), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_299), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_318), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_314), .B(n_299), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_305), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_359), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_348), .B(n_307), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_345), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_336), .B(n_338), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_359), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_336), .B(n_314), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_341), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_338), .B(n_318), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_304), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_343), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_342), .B(n_317), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_342), .B(n_317), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_331), .B(n_325), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_350), .B(n_325), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_352), .B(n_328), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_350), .B(n_328), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_356), .B(n_305), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_328), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_335), .B(n_319), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_319), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_358), .B(n_319), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_337), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_332), .B(n_310), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_348), .B(n_321), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_358), .B(n_321), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_357), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_359), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_321), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_353), .B(n_321), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_359), .B(n_323), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_359), .B(n_326), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_345), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_379), .B(n_355), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_368), .B(n_340), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
INVx3_ASAP7_75t_SL g411 ( .A(n_361), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_355), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_369), .B(n_349), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_365), .B(n_360), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_372), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_372), .B(n_353), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_367), .B(n_360), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_373), .B(n_347), .C(n_329), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_364), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_375), .B(n_357), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_379), .B(n_357), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_376), .B(n_329), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_382), .B(n_329), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_377), .B(n_329), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_382), .B(n_344), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_371), .B(n_344), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_367), .B(n_344), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_398), .B(n_344), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_371), .B(n_339), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_405), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_339), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_377), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_406), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_381), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_390), .B(n_347), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_390), .B(n_333), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_359), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_370), .B(n_339), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_397), .B(n_310), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_397), .A2(n_302), .B1(n_326), .B2(n_310), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_384), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_396), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_361), .B(n_283), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_385), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_391), .B(n_333), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_391), .B(n_383), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_397), .B(n_333), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_395), .B(n_283), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_449), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_457), .B(n_399), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_440), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_423), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_410), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_459), .A2(n_386), .B(n_389), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_414), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_416), .B(n_370), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_451), .B(n_401), .C(n_397), .D(n_363), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_416), .B(n_401), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_454), .A2(n_361), .B1(n_366), .B2(n_323), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_455), .B(n_383), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_441), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_442), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_409), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_457), .B(n_399), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_434), .B(n_378), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_437), .A2(n_402), .B(n_363), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_461), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_412), .B(n_378), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_420), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_444), .B(n_374), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_415), .B(n_363), .Y(n_493) );
NOR2xp67_ASAP7_75t_SL g494 ( .A(n_438), .B(n_283), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_444), .B(n_374), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_413), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_458), .B(n_363), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_413), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_458), .B(n_402), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_420), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_445), .B(n_404), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_408), .B(n_394), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_437), .B(n_361), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_445), .B(n_362), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_407), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_453), .Y(n_507) );
NOR2x2_ASAP7_75t_L g508 ( .A(n_421), .B(n_394), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_484), .B(n_456), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_488), .B(n_456), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_469), .A2(n_428), .B1(n_422), .B2(n_419), .C1(n_450), .C2(n_435), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_492), .B(n_426), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_489), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_475), .A2(n_428), .B(n_403), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_496), .B(n_431), .Y(n_516) );
OAI32xp33_ASAP7_75t_L g517 ( .A1(n_475), .A2(n_366), .A3(n_436), .B1(n_432), .B2(n_430), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_470), .A2(n_418), .B(n_425), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_491), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_469), .A2(n_427), .B1(n_431), .B2(n_448), .C1(n_447), .C2(n_418), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_498), .B(n_427), .Y(n_521) );
AOI321xp33_ASAP7_75t_L g522 ( .A1(n_471), .A2(n_433), .A3(n_425), .B1(n_366), .B2(n_403), .C(n_287), .Y(n_522) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_475), .B(n_403), .Y(n_523) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_487), .A2(n_392), .B(n_362), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_509), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_499), .B(n_403), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_465), .B(n_392), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_508), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_500), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_481), .A2(n_327), .B(n_279), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_501), .B(n_380), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_463), .B(n_333), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
AOI222xp33_ASAP7_75t_L g536 ( .A1(n_504), .A2(n_288), .B1(n_380), .B2(n_290), .C1(n_303), .C2(n_327), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_499), .B(n_315), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_501), .B(n_315), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_505), .B(n_315), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_505), .B(n_311), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_529), .A2(n_504), .B(n_502), .C(n_471), .Y(n_543) );
AND4x1_ASAP7_75t_L g544 ( .A(n_512), .B(n_494), .C(n_506), .D(n_508), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_518), .A2(n_467), .B1(n_495), .B2(n_483), .C(n_482), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g547 ( .A1(n_530), .A2(n_519), .B(n_514), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_529), .A2(n_502), .B1(n_497), .B2(n_474), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_516), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_515), .B(n_472), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_523), .A2(n_497), .B1(n_490), .B2(n_463), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_517), .A2(n_480), .B1(n_479), .B2(n_485), .C(n_497), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_530), .A2(n_485), .B1(n_486), .B2(n_503), .C(n_507), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_521), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_528), .A2(n_520), .B(n_531), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_526), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_522), .B(n_507), .C(n_478), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_524), .B(n_294), .Y(n_558) );
AOI221x1_ASAP7_75t_L g559 ( .A1(n_525), .A2(n_478), .B1(n_477), .B2(n_464), .C(n_493), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_534), .A2(n_539), .B1(n_528), .B2(n_510), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_534), .A2(n_486), .B1(n_477), .B2(n_464), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_511), .A2(n_524), .B(n_540), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_536), .A2(n_311), .B(n_299), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_532), .A2(n_290), .B(n_311), .C(n_294), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_541), .B(n_303), .C(n_327), .Y(n_565) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_542), .A2(n_285), .B(n_292), .C(n_311), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_535), .Y(n_567) );
A2O1A1O1Ixp25_ASAP7_75t_L g568 ( .A1(n_537), .A2(n_294), .B(n_293), .C(n_296), .D(n_308), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_538), .B(n_293), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_533), .A2(n_293), .B1(n_292), .B2(n_296), .C(n_308), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_527), .A2(n_293), .B(n_296), .C(n_308), .Y(n_571) );
AOI211xp5_ASAP7_75t_L g572 ( .A1(n_513), .A2(n_296), .B(n_308), .C(n_280), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_550), .B(n_552), .C(n_555), .Y(n_573) );
AOI211xp5_ASAP7_75t_SL g574 ( .A1(n_563), .A2(n_547), .B(n_548), .C(n_551), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_557), .B(n_546), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_543), .A2(n_545), .B(n_559), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_553), .A2(n_564), .B(n_562), .C(n_544), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_560), .A2(n_561), .B(n_566), .C(n_558), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_575), .B(n_549), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_573), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_574), .B(n_554), .Y(n_581) );
OAI22x1_ASAP7_75t_L g582 ( .A1(n_580), .A2(n_576), .B1(n_577), .B2(n_556), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_579), .B(n_578), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_583), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_582), .B(n_581), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_567), .B1(n_569), .B2(n_524), .Y(n_586) );
OAI22x1_ASAP7_75t_L g587 ( .A1(n_586), .A2(n_584), .B1(n_296), .B2(n_568), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_565), .B1(n_571), .B2(n_570), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_588), .B(n_308), .Y(n_589) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_589), .A2(n_572), .B(n_280), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_590), .A2(n_280), .B1(n_584), .B2(n_580), .Y(n_591) );
endmodule