module fake_jpeg_22539_n_288 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_28),
.B(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_48),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_34),
.B1(n_14),
.B2(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_54),
.B1(n_44),
.B2(n_49),
.Y(n_79)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_39),
.A2(n_24),
.B1(n_14),
.B2(n_16),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_68),
.B1(n_50),
.B2(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_62),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_46),
.B(n_16),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_18),
.B(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_38),
.C(n_35),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_100),
.C(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_28),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_21),
.B(n_38),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_95),
.B(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_69),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_33),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_70),
.B1(n_73),
.B2(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_117),
.C(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_65),
.B1(n_70),
.B2(n_37),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_22),
.B1(n_69),
.B2(n_26),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_65),
.B1(n_37),
.B2(n_50),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_52),
.B1(n_72),
.B2(n_73),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_80),
.B1(n_88),
.B2(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_52),
.B1(n_76),
.B2(n_71),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_24),
.B1(n_67),
.B2(n_61),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_118),
.B1(n_79),
.B2(n_96),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_36),
.C(n_17),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_90),
.B1(n_95),
.B2(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_122),
.B(n_84),
.Y(n_125)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_132),
.C(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_125),
.B(n_141),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_83),
.B(n_85),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_138),
.B(n_102),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_86),
.B(n_87),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_101),
.B(n_114),
.Y(n_156)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_135),
.B1(n_107),
.B2(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_97),
.B1(n_93),
.B2(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_142),
.B1(n_147),
.B2(n_108),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_99),
.B(n_92),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_119),
.C(n_117),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_24),
.B1(n_92),
.B2(n_27),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_137),
.B1(n_126),
.B2(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_101),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_151),
.B1(n_166),
.B2(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_121),
.B1(n_101),
.B2(n_117),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_160),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_112),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_27),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_27),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_104),
.B1(n_26),
.B2(n_25),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_26),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_132),
.C(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_13),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_170),
.A2(n_137),
.B(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_25),
.B1(n_20),
.B2(n_2),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_20),
.B1(n_13),
.B2(n_12),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_124),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_184),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_195),
.B1(n_149),
.B2(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_187),
.C(n_165),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_193),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_127),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_160),
.B1(n_157),
.B2(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_166),
.B1(n_172),
.B2(n_164),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_139),
.C(n_142),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_139),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_191),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_128),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_143),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_128),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_156),
.C(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_204),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_165),
.B1(n_153),
.B2(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_153),
.C(n_167),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_174),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_167),
.B(n_162),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_212),
.B(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_171),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_179),
.A2(n_173),
.B1(n_186),
.B2(n_194),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_208),
.B1(n_197),
.B2(n_206),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_11),
.B(n_3),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_11),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_230),
.B(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_198),
.C(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_188),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_232),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_187),
.B1(n_176),
.B2(n_189),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_224),
.B1(n_216),
.B2(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_184),
.B(n_3),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_10),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_212),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_4),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_248),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_205),
.C(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_202),
.C(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_4),
.C(n_5),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_219),
.C(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_5),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_5),
.CI(n_6),
.CON(n_248),
.SN(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_222),
.B(n_221),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_258),
.B(n_7),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_233),
.B1(n_220),
.B2(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_260),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_6),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_6),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_259),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_7),
.B(n_8),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_7),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_239),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_265),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_244),
.B1(n_240),
.B2(n_248),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_266),
.A2(n_252),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_234),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_249),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_8),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_275),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_249),
.B(n_256),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_281),
.C(n_261),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_276),
.C(n_271),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_283),
.B(n_279),
.C(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_285),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_8),
.C(n_10),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_10),
.Y(n_288)
);


endmodule