module fake_jpeg_4290_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_0),
.C(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_14),
.C(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_7),
.B1(n_11),
.B2(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_22),
.B1(n_11),
.B2(n_19),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_7),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_23),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_11),
.B1(n_24),
.B2(n_17),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_9),
.C(n_13),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_26),
.C(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_4),
.B1(n_36),
.B2(n_39),
.Y(n_41)
);


endmodule