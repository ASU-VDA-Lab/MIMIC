module fake_jpeg_16663_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_19),
.Y(n_66)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_45),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_58),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_72),
.B1(n_17),
.B2(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_17),
.B1(n_30),
.B2(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_28),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_32),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_19),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_17),
.B(n_30),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_88),
.B1(n_94),
.B2(n_105),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_45),
.B1(n_44),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_87),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_45),
.B1(n_32),
.B2(n_21),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_35),
.B1(n_21),
.B2(n_31),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_84),
.B(n_97),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_16),
.B1(n_33),
.B2(n_27),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_35),
.B1(n_21),
.B2(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_108),
.B1(n_64),
.B2(n_54),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_68),
.B1(n_48),
.B2(n_73),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_0),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_56),
.A2(n_51),
.B1(n_75),
.B2(n_70),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_23),
.B1(n_20),
.B2(n_49),
.Y(n_118)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_16),
.B(n_24),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_112),
.B(n_110),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_129),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_74),
.B(n_48),
.C(n_68),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_124),
.B(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_132),
.B1(n_139),
.B2(n_106),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_122),
.B1(n_99),
.B2(n_81),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_20),
.A3(n_23),
.B1(n_26),
.B2(n_10),
.Y(n_122)
);

AOI22x1_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_23),
.B1(n_64),
.B2(n_54),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_9),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_108),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_54),
.C(n_8),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_77),
.C(n_92),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_76),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_0),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_152),
.B(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_87),
.B1(n_95),
.B2(n_93),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_99),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_164),
.Y(n_178)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_149),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_171),
.B(n_164),
.Y(n_188)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_104),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_95),
.B1(n_96),
.B2(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_133),
.B1(n_118),
.B2(n_122),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_81),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_116),
.B(n_117),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_159),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_135),
.Y(n_186)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_80),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_174),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_84),
.B1(n_96),
.B2(n_111),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_109),
.B1(n_92),
.B2(n_79),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_175),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_120),
.A2(n_78),
.B1(n_79),
.B2(n_109),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_1),
.B(n_3),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_78),
.B1(n_10),
.B2(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_109),
.Y(n_174)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_125),
.A2(n_78),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_9),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_157),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_209),
.C(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_154),
.B1(n_185),
.B2(n_144),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_121),
.B1(n_139),
.B2(n_123),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_175),
.B1(n_145),
.B2(n_169),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_139),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_192),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_152),
.A2(n_126),
.B1(n_123),
.B2(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_170),
.B(n_175),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_138),
.C(n_126),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_138),
.C(n_11),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_150),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_212),
.A2(n_183),
.B(n_196),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_179),
.C(n_190),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_233),
.C(n_209),
.Y(n_239)
);

OR2x6_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_145),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_229),
.B(n_231),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_227),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_143),
.CI(n_148),
.CON(n_227),
.SN(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_145),
.C(n_159),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_177),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_158),
.C(n_169),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_182),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_255),
.C(n_217),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_262),
.Y(n_268)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_225),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_222),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_246),
.B(n_247),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_193),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_180),
.B1(n_199),
.B2(n_198),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_234),
.B(n_222),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_194),
.B1(n_182),
.B2(n_210),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_212),
.B(n_184),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_194),
.C(n_205),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_203),
.B1(n_201),
.B2(n_204),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_195),
.B1(n_202),
.B2(n_197),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_195),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_261),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_197),
.B1(n_191),
.B2(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_260),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_191),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_271),
.C(n_281),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_221),
.C(n_214),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_245),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_227),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_227),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_250),
.B(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_216),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_228),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_254),
.B(n_218),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_253),
.C(n_259),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_244),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_296),
.B(n_282),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_258),
.B(n_261),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_6),
.B(n_12),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_265),
.A2(n_243),
.B1(n_281),
.B2(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_297),
.B1(n_7),
.B2(n_14),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_269),
.A3(n_271),
.B1(n_280),
.B2(n_264),
.C(n_268),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_247),
.B1(n_241),
.B2(n_242),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_292),
.B1(n_272),
.B2(n_282),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_219),
.B1(n_257),
.B2(n_253),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_213),
.B(n_230),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_207),
.B1(n_169),
.B2(n_5),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_305),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_266),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_311),
.B1(n_298),
.B2(n_294),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_9),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_3),
.C(n_4),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_12),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_292),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_4),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_291),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_288),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_305),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_290),
.A3(n_300),
.B1(n_284),
.B2(n_13),
.C1(n_15),
.C2(n_12),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_308),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_307),
.B(n_297),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_328),
.B(n_329),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_322),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_318),
.C(n_317),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_330),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_314),
.B(n_313),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_332),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_318),
.B(n_5),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);


endmodule