module fake_jpeg_25530_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_20),
.Y(n_51)
);

AO22x2_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_39),
.B1(n_35),
.B2(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_55),
.B1(n_33),
.B2(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_51),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_15),
.B1(n_22),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_28),
.B1(n_15),
.B2(n_25),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_15),
.B1(n_30),
.B2(n_27),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_25),
.B(n_24),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_20),
.B1(n_30),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_33),
.B1(n_32),
.B2(n_19),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_20),
.B1(n_24),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_35),
.B1(n_32),
.B2(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_66),
.B1(n_34),
.B2(n_36),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_16),
.Y(n_106)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_82),
.Y(n_91)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_69),
.Y(n_92)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_31),
.C(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_36),
.Y(n_104)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_18),
.B1(n_16),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_72),
.B1(n_85),
.B2(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_11),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_89),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_95),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_103),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_72),
.C(n_66),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_108),
.C(n_4),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_70),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_77),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_113),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_74),
.B1(n_65),
.B2(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_109),
.B1(n_98),
.B2(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_23),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_23),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_0),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_1),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_108),
.B1(n_107),
.B2(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_2),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_130),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_3),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_116),
.B(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_90),
.B(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_130),
.B(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_141),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_102),
.A3(n_89),
.B1(n_99),
.B2(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_5),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_110),
.B1(n_111),
.B2(n_124),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_148),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_151),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_118),
.C(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_156),
.C(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_158),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_138),
.C(n_136),
.Y(n_156)
);

AO21x1_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_92),
.B(n_6),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_5),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_162),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_131),
.B1(n_139),
.B2(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_150),
.B1(n_142),
.B2(n_141),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_144),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_149),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_162),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_147),
.C(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_139),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_161),
.C(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_160),
.C(n_167),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_172),
.B1(n_169),
.B2(n_173),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_158),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_7),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_177),
.B(n_180),
.Y(n_191)
);

OAI31xp33_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_192),
.A3(n_8),
.B(n_9),
.Y(n_195)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_182),
.A3(n_174),
.B(n_175),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_179),
.B(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_187),
.B1(n_184),
.B2(n_176),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_8),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_SL g198 ( 
.A(n_196),
.B(n_8),
.C(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_196),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_197),
.Y(n_200)
);


endmodule