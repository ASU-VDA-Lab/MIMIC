module real_aes_17737_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_0), .A2(n_201), .B1(n_1134), .B2(n_1138), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_1), .A2(n_206), .B1(n_434), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_1), .A2(n_59), .B1(n_338), .B2(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g691 ( .A(n_2), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_2), .A2(n_95), .B1(n_434), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_3), .A2(n_116), .B1(n_341), .B2(n_346), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_3), .A2(n_123), .B1(n_431), .B2(n_433), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_4), .A2(n_51), .B1(n_1134), .B2(n_1138), .Y(n_1163) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_5), .A2(n_149), .B1(n_337), .B2(n_499), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g1035 ( .A(n_5), .Y(n_1035) );
XNOR2x2_ASAP7_75t_L g555 ( .A(n_6), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g789 ( .A(n_7), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_7), .A2(n_60), .B1(n_361), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_8), .A2(n_217), .B1(n_434), .B2(n_780), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_8), .A2(n_253), .B1(n_338), .B2(n_621), .Y(n_841) );
INVx1_ASAP7_75t_L g280 ( .A(n_9), .Y(n_280) );
AND2x2_ASAP7_75t_L g387 ( .A(n_9), .B(n_226), .Y(n_387) );
AND2x2_ASAP7_75t_L g413 ( .A(n_9), .B(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_9), .B(n_290), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_10), .A2(n_166), .B1(n_330), .B2(n_337), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_10), .A2(n_17), .B1(n_417), .B2(n_421), .C(n_428), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_11), .A2(n_43), .B1(n_372), .B2(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g595 ( .A(n_11), .Y(n_595) );
INVx1_ASAP7_75t_L g1049 ( .A(n_12), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_12), .A2(n_161), .B1(n_521), .B2(n_599), .C(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_13), .A2(n_68), .B1(n_434), .B2(n_721), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_13), .A2(n_135), .B1(n_338), .B2(n_499), .Y(n_1113) );
INVx2_ASAP7_75t_L g1137 ( .A(n_14), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_14), .B(n_96), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_14), .B(n_1143), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_15), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_16), .A2(n_84), .B1(n_403), .B2(n_679), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_17), .A2(n_33), .B1(n_358), .B2(n_359), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_18), .A2(n_243), .B1(n_569), .B2(n_1116), .Y(n_1348) );
INVx1_ASAP7_75t_L g1370 ( .A(n_18), .Y(n_1370) );
AOI22xp33_ASAP7_75t_SL g1351 ( .A1(n_19), .A2(n_192), .B1(n_499), .B2(n_693), .Y(n_1351) );
INVxp67_ASAP7_75t_SL g1356 ( .A(n_19), .Y(n_1356) );
INVx1_ASAP7_75t_L g315 ( .A(n_20), .Y(n_315) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_21), .A2(n_210), .B1(n_361), .B2(n_372), .Y(n_360) );
INVx1_ASAP7_75t_L g441 ( .A(n_21), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_22), .A2(n_32), .B1(n_1141), .B2(n_1144), .Y(n_1155) );
XNOR2xp5_ASAP7_75t_L g1393 ( .A(n_23), .B(n_1394), .Y(n_1393) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_24), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g636 ( .A(n_25), .Y(n_636) );
INVx1_ASAP7_75t_L g715 ( .A(n_26), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_27), .A2(n_66), .B1(n_499), .B2(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_27), .A2(n_263), .B1(n_418), .B2(n_428), .C(n_642), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_28), .A2(n_115), .B1(n_1141), .B2(n_1144), .Y(n_1172) );
INVx1_ASAP7_75t_L g714 ( .A(n_29), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_30), .A2(n_90), .B1(n_403), .B2(n_679), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_31), .A2(n_263), .B1(n_499), .B2(n_693), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_31), .A2(n_66), .B1(n_658), .B2(n_721), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_33), .A2(n_446), .B(n_450), .C(n_462), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_34), .A2(n_159), .B1(n_499), .B2(n_564), .Y(n_563) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_34), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g1057 ( .A1(n_35), .A2(n_81), .B1(n_358), .B2(n_564), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_35), .A2(n_170), .B1(n_428), .B2(n_1040), .C(n_1075), .Y(n_1074) );
XNOR2xp5_ASAP7_75t_L g813 ( .A(n_36), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_36), .A2(n_89), .B1(n_1134), .B2(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g774 ( .A(n_37), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_38), .A2(n_83), .B1(n_1134), .B2(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1380 ( .A(n_38), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_38), .A2(n_1387), .B1(n_1392), .B2(n_1396), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_39), .A2(n_55), .B1(n_393), .B2(n_403), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_39), .A2(n_408), .B(n_415), .C(n_436), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_40), .A2(n_171), .B1(n_434), .B2(n_786), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g843 ( .A1(n_40), .A2(n_118), .B1(n_375), .B2(n_490), .Y(n_843) );
INVx1_ASAP7_75t_L g939 ( .A(n_41), .Y(n_939) );
XNOR2x2_ASAP7_75t_L g296 ( .A(n_42), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g594 ( .A(n_43), .Y(n_594) );
AOI21xp33_ASAP7_75t_L g743 ( .A1(n_44), .A2(n_642), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g752 ( .A(n_44), .Y(n_752) );
INVx1_ASAP7_75t_L g322 ( .A(n_45), .Y(n_322) );
INVx1_ASAP7_75t_L g336 ( .A(n_45), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_46), .A2(n_130), .B1(n_642), .B2(n_823), .C(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_46), .A2(n_196), .B1(n_375), .B2(n_490), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_47), .A2(n_69), .B1(n_494), .B2(n_498), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_47), .A2(n_245), .B1(n_507), .B2(n_508), .C(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g677 ( .A(n_48), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_49), .A2(n_200), .B1(n_431), .B2(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g753 ( .A(n_49), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_50), .A2(n_125), .B1(n_1134), .B2(n_1149), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_52), .A2(n_224), .B1(n_1141), .B2(n_1144), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_53), .A2(n_123), .B1(n_346), .B2(n_349), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_53), .A2(n_116), .B1(n_452), .B2(n_455), .C(n_458), .Y(n_451) );
INVx1_ASAP7_75t_L g273 ( .A(n_54), .Y(n_273) );
INVx2_ASAP7_75t_L g312 ( .A(n_56), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_57), .A2(n_232), .B1(n_428), .B2(n_730), .C(n_731), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_57), .A2(n_262), .B1(n_338), .B2(n_499), .Y(n_754) );
INVx1_ASAP7_75t_L g1342 ( .A(n_58), .Y(n_1342) );
OAI222xp33_ASAP7_75t_L g1366 ( .A1(n_58), .A2(n_241), .B1(n_521), .B2(n_543), .C1(n_1367), .C2(n_1371), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_59), .A2(n_198), .B1(n_418), .B2(n_428), .C(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g788 ( .A(n_60), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_61), .A2(n_140), .B1(n_490), .B2(n_492), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_61), .A2(n_143), .B1(n_511), .B2(n_514), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_62), .A2(n_63), .B1(n_359), .B2(n_499), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_62), .A2(n_149), .B1(n_509), .B2(n_1022), .C(n_1024), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1037 ( .A(n_63), .Y(n_1037) );
AOI22xp33_ASAP7_75t_SL g1006 ( .A1(n_64), .A2(n_191), .B1(n_1007), .B2(n_1009), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_64), .A2(n_129), .B1(n_431), .B2(n_433), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_65), .A2(n_187), .B1(n_564), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_65), .A2(n_234), .B1(n_431), .B2(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g1379 ( .A(n_67), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_68), .A2(n_260), .B1(n_499), .B2(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g541 ( .A(n_69), .Y(n_541) );
INVx1_ASAP7_75t_L g965 ( .A(n_70), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_70), .A2(n_126), .B1(n_642), .B2(n_730), .C(n_979), .Y(n_978) );
AOI21xp33_ASAP7_75t_L g778 ( .A1(n_71), .A2(n_731), .B(n_744), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_71), .A2(n_179), .B1(n_490), .B2(n_802), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1013 ( .A1(n_72), .A2(n_256), .B1(n_361), .B2(n_372), .Y(n_1013) );
INVx1_ASAP7_75t_L g1029 ( .A(n_72), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_73), .A2(n_181), .B1(n_351), .B2(n_1055), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_73), .A2(n_78), .B1(n_780), .B2(n_1072), .Y(n_1071) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_74), .A2(n_598), .B(n_771), .C(n_775), .Y(n_770) );
INVx1_ASAP7_75t_L g797 ( .A(n_74), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_75), .A2(n_99), .B1(n_1134), .B2(n_1138), .Y(n_1133) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_76), .A2(n_117), .B1(n_1141), .B2(n_1144), .Y(n_1195) );
INVx1_ASAP7_75t_L g485 ( .A(n_77), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g503 ( .A1(n_77), .A2(n_504), .B(n_505), .C(n_516), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_78), .A2(n_100), .B1(n_1007), .B2(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g818 ( .A(n_79), .Y(n_818) );
INVx1_ASAP7_75t_L g1344 ( .A(n_80), .Y(n_1344) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_81), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_82), .A2(n_128), .B1(n_393), .B2(n_581), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g825 ( .A1(n_84), .A2(n_504), .B(n_826), .C(n_830), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_85), .Y(n_550) );
INVx1_ASAP7_75t_L g877 ( .A(n_86), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_86), .A2(n_218), .B1(n_759), .B2(n_905), .C(n_907), .Y(n_904) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_87), .Y(n_275) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_87), .B(n_273), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_88), .A2(n_265), .B1(n_624), .B2(n_626), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_88), .A2(n_533), .B(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g781 ( .A1(n_90), .A2(n_408), .B(n_782), .C(n_787), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_91), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_92), .A2(n_252), .B1(n_372), .B2(n_575), .Y(n_637) );
INVx1_ASAP7_75t_L g645 ( .A(n_92), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_93), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_94), .A2(n_124), .B1(n_490), .B2(n_566), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_94), .A2(n_177), .B1(n_533), .B2(n_606), .C(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g701 ( .A(n_95), .Y(n_701) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_96), .B(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1143 ( .A(n_96), .Y(n_1143) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_97), .A2(n_230), .B1(n_930), .B2(n_933), .Y(n_929) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_97), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_98), .A2(n_173), .B1(n_1141), .B2(n_1144), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_100), .A2(n_181), .B1(n_507), .B2(n_533), .C(n_590), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_101), .A2(n_174), .B1(n_372), .B2(n_575), .Y(n_1058) );
INVx1_ASAP7_75t_L g1080 ( .A(n_101), .Y(n_1080) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_102), .A2(n_196), .B1(n_721), .B2(n_734), .Y(n_1102) );
AOI22xp5_ASAP7_75t_L g1115 ( .A1(n_102), .A2(n_130), .B1(n_490), .B2(n_1116), .Y(n_1115) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_103), .A2(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g1100 ( .A(n_104), .Y(n_1100) );
INVx1_ASAP7_75t_L g1105 ( .A(n_105), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_106), .A2(n_245), .B1(n_492), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g531 ( .A(n_106), .Y(n_531) );
INVx1_ASAP7_75t_L g686 ( .A(n_107), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_107), .A2(n_533), .B(n_642), .Y(n_719) );
INVx2_ASAP7_75t_L g314 ( .A(n_108), .Y(n_314) );
INVx1_ASAP7_75t_L g356 ( .A(n_108), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_108), .B(n_312), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_109), .A2(n_157), .B1(n_347), .B2(n_910), .Y(n_969) );
INVx1_ASAP7_75t_L g980 ( .A(n_109), .Y(n_980) );
AOI21xp33_ASAP7_75t_L g821 ( .A1(n_110), .A2(n_822), .B(n_823), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_110), .A2(n_171), .B1(n_490), .B2(n_802), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_111), .Y(n_517) );
INVx1_ASAP7_75t_L g561 ( .A(n_112), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g597 ( .A1(n_112), .A2(n_193), .B1(n_598), .B2(n_599), .C(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g889 ( .A(n_113), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_114), .A2(n_150), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_114), .A2(n_205), .B1(n_490), .B2(n_909), .Y(n_908) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_118), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_119), .A2(n_228), .B1(n_581), .B2(n_679), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_119), .A2(n_504), .B(n_708), .C(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g1363 ( .A(n_120), .Y(n_1363) );
INVx1_ASAP7_75t_L g834 ( .A(n_121), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_122), .A2(n_239), .B1(n_1141), .B2(n_1144), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_124), .A2(n_180), .B1(n_586), .B2(n_587), .Y(n_585) );
XNOR2xp5_ASAP7_75t_L g940 ( .A(n_125), .B(n_941), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g958 ( .A1(n_126), .A2(n_244), .B1(n_339), .B2(n_959), .C(n_960), .Y(n_958) );
XOR2x2_ASAP7_75t_L g1043 ( .A(n_127), .B(n_1044), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_127), .A2(n_131), .B1(n_1134), .B2(n_1138), .Y(n_1194) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_128), .A2(n_408), .B(n_584), .C(n_593), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_129), .A2(n_238), .B1(n_1007), .B2(n_1009), .Y(n_1010) );
INVx1_ASAP7_75t_L g832 ( .A(n_132), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_132), .A2(n_184), .B1(n_575), .B2(n_809), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_133), .A2(n_207), .B1(n_499), .B2(n_1347), .Y(n_1346) );
INVxp67_ASAP7_75t_SL g1372 ( .A(n_133), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_134), .A2(n_163), .B1(n_568), .B2(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1369 ( .A(n_134), .Y(n_1369) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_135), .A2(n_260), .B1(n_423), .B2(n_592), .C(n_730), .Y(n_1101) );
INVx1_ASAP7_75t_L g1104 ( .A(n_136), .Y(n_1104) );
INVx1_ASAP7_75t_L g737 ( .A(n_137), .Y(n_737) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_138), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_138), .A2(n_504), .B(n_640), .C(n_644), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_139), .A2(n_248), .B1(n_624), .B2(n_626), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_139), .A2(n_265), .B1(n_434), .B2(n_512), .Y(n_643) );
INVx1_ASAP7_75t_L g526 ( .A(n_140), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g1106 ( .A1(n_141), .A2(n_679), .B(n_1107), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_142), .A2(n_146), .B1(n_1141), .B2(n_1144), .Y(n_1162) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_143), .A2(n_145), .B1(n_489), .B2(n_490), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_144), .A2(n_258), .B1(n_930), .B2(n_933), .Y(n_948) );
INVxp33_ASAP7_75t_SL g989 ( .A(n_144), .Y(n_989) );
INVx1_ASAP7_75t_L g535 ( .A(n_145), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_147), .A2(n_262), .B1(n_410), .B2(n_721), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_147), .A2(n_232), .B1(n_499), .B2(n_759), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_148), .A2(n_178), .B1(n_393), .B2(n_581), .Y(n_1017) );
OAI211xp5_ASAP7_75t_SL g1019 ( .A1(n_148), .A2(n_408), .B(n_1020), .C(n_1026), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_150), .A2(n_250), .B1(n_626), .B2(n_902), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g1375 ( .A1(n_151), .A2(n_679), .B(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g736 ( .A(n_152), .Y(n_736) );
INVx1_ASAP7_75t_L g1362 ( .A(n_153), .Y(n_1362) );
INVx1_ASAP7_75t_L g615 ( .A(n_154), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_154), .A2(n_156), .B1(n_521), .B2(n_543), .C(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g306 ( .A(n_155), .Y(n_306) );
INVx1_ASAP7_75t_L g616 ( .A(n_156), .Y(n_616) );
INVx1_ASAP7_75t_L g974 ( .A(n_157), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_158), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_159), .A2(n_237), .B1(n_589), .B2(n_590), .C(n_592), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_160), .A2(n_234), .B1(n_489), .B2(n_564), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_160), .A2(n_187), .B1(n_418), .B2(n_428), .C(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g1048 ( .A(n_161), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1150 ( .A1(n_162), .A2(n_165), .B1(n_1141), .B2(n_1144), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1359 ( .A1(n_163), .A2(n_243), .B1(n_434), .B2(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g955 ( .A(n_164), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_164), .A2(n_199), .B1(n_642), .B2(n_730), .C(n_973), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_166), .B(n_461), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_167), .A2(n_227), .B1(n_1134), .B2(n_1138), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_168), .A2(n_253), .B1(n_418), .B2(n_509), .C(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_168), .A2(n_217), .B1(n_359), .B2(n_489), .Y(n_844) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_170), .A2(n_231), .B1(n_359), .B2(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g943 ( .A(n_172), .Y(n_943) );
INVx1_ASAP7_75t_L g1079 ( .A(n_174), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_175), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g872 ( .A1(n_176), .A2(n_205), .B1(n_855), .B2(n_873), .C(n_875), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g903 ( .A1(n_176), .A2(n_211), .B1(n_499), .B2(n_564), .C(n_806), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_177), .A2(n_180), .B1(n_566), .B2(n_569), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_179), .A2(n_246), .B1(n_434), .B2(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g963 ( .A(n_182), .Y(n_963) );
INVx1_ASAP7_75t_L g1087 ( .A(n_183), .Y(n_1087) );
INVx1_ASAP7_75t_L g831 ( .A(n_184), .Y(n_831) );
XOR2xp5_ASAP7_75t_L g997 ( .A(n_185), .B(n_998), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_186), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_188), .A2(n_235), .B1(n_521), .B2(n_543), .C(n_739), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_188), .A2(n_235), .B1(n_481), .B2(n_704), .Y(n_760) );
INVx1_ASAP7_75t_L g482 ( .A(n_189), .Y(n_482) );
OAI222xp33_ASAP7_75t_L g520 ( .A1(n_189), .A2(n_259), .B1(n_521), .B2(n_522), .C1(n_534), .C2(n_542), .Y(n_520) );
INVx1_ASAP7_75t_L g551 ( .A(n_190), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_191), .A2(n_238), .B1(n_458), .B2(n_1039), .C(n_1040), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_192), .Y(n_1374) );
INVx1_ASAP7_75t_L g560 ( .A(n_193), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_194), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_195), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_197), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_198), .A2(n_206), .B1(n_359), .B2(n_800), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g968 ( .A1(n_199), .A2(n_351), .B(n_907), .Y(n_968) );
INVx1_ASAP7_75t_L g757 ( .A(n_200), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_202), .Y(n_391) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_203), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_203), .A2(n_246), .B1(n_346), .B2(n_375), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_204), .Y(n_1016) );
AOI21xp33_ASAP7_75t_L g1358 ( .A1(n_207), .A2(n_592), .B(n_822), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_208), .B(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_208), .A2(n_632), .B1(n_633), .B2(n_664), .Y(n_631) );
INVx1_ASAP7_75t_L g666 ( .A(n_208), .Y(n_666) );
OA22x2_ASAP7_75t_L g767 ( .A1(n_209), .A2(n_768), .B1(n_811), .B2(n_812), .Y(n_767) );
CKINVDCx16_ASAP7_75t_R g811 ( .A(n_209), .Y(n_811) );
INVx1_ASAP7_75t_L g437 ( .A(n_210), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_211), .A2(n_218), .B1(n_857), .B2(n_859), .C(n_861), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_212), .A2(n_229), .B1(n_393), .B2(n_581), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g1083 ( .A1(n_213), .A2(n_1084), .B1(n_1085), .B2(n_1119), .Y(n_1083) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_213), .Y(n_1119) );
INVx1_ASAP7_75t_L g301 ( .A(n_214), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_215), .A2(n_264), .B1(n_581), .B2(n_679), .Y(n_763) );
INVx1_ASAP7_75t_L g1002 ( .A(n_216), .Y(n_1002) );
OAI221xp5_ASAP7_75t_SL g1030 ( .A1(n_216), .A2(n_261), .B1(n_542), .B2(n_598), .C(n_1031), .Y(n_1030) );
INVxp67_ASAP7_75t_SL g892 ( .A(n_219), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_219), .A2(n_222), .B1(n_922), .B2(n_924), .C(n_926), .Y(n_921) );
INVx1_ASAP7_75t_L g762 ( .A(n_220), .Y(n_762) );
OAI211xp5_ASAP7_75t_SL g949 ( .A1(n_221), .A2(n_919), .B(n_926), .C(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g985 ( .A(n_221), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_222), .A2(n_233), .B1(n_864), .B2(n_869), .C(n_870), .Y(n_863) );
OAI211xp5_ASAP7_75t_L g816 ( .A1(n_223), .A2(n_598), .B(n_817), .C(n_819), .Y(n_816) );
INVx1_ASAP7_75t_L g839 ( .A(n_223), .Y(n_839) );
INVx1_ASAP7_75t_L g1092 ( .A(n_225), .Y(n_1092) );
BUFx3_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
INVx1_ASAP7_75t_L g414 ( .A(n_226), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g1069 ( .A1(n_229), .A2(n_504), .B(n_1070), .C(n_1078), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g884 ( .A(n_230), .Y(n_884) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_231), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_233), .A2(n_236), .B1(n_912), .B2(n_915), .Y(n_911) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_236), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_237), .A2(n_249), .B1(n_499), .B2(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g309 ( .A(n_240), .Y(n_309) );
INVx2_ASAP7_75t_L g328 ( .A(n_240), .Y(n_328) );
INVx1_ASAP7_75t_L g370 ( .A(n_240), .Y(n_370) );
INVx1_ASAP7_75t_L g1341 ( .A(n_241), .Y(n_1341) );
INVx1_ASAP7_75t_L g1094 ( .A(n_242), .Y(n_1094) );
INVx1_ASAP7_75t_L g975 ( .A(n_244), .Y(n_975) );
INVx1_ASAP7_75t_L g791 ( .A(n_247), .Y(n_791) );
INVx1_ASAP7_75t_L g650 ( .A(n_248), .Y(n_650) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_249), .Y(n_604) );
INVx1_ASAP7_75t_L g876 ( .A(n_250), .Y(n_876) );
OAI22xp33_ASAP7_75t_SL g703 ( .A1(n_251), .A2(n_257), .B1(n_481), .B2(n_704), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_251), .A2(n_257), .B1(n_543), .B2(n_598), .C(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g647 ( .A(n_252), .Y(n_647) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_254), .B(n_675), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_255), .Y(n_957) );
INVx1_ASAP7_75t_L g1027 ( .A(n_256), .Y(n_1027) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_258), .Y(n_946) );
INVx1_ASAP7_75t_L g479 ( .A(n_259), .Y(n_479) );
INVx1_ASAP7_75t_L g1003 ( .A(n_261), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g727 ( .A1(n_264), .A2(n_504), .B(n_728), .C(n_735), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_291), .B(n_1122), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_276), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_270), .B(n_279), .Y(n_1385) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_272), .B(n_275), .Y(n_1391) );
INVx1_ASAP7_75t_L g1398 ( .A(n_272), .Y(n_1398) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_275), .B(n_1398), .Y(n_1400) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g429 ( .A(n_280), .B(n_290), .Y(n_429) );
AND2x4_ASAP7_75t_L g459 ( .A(n_280), .B(n_289), .Y(n_459) );
AND2x4_ASAP7_75t_SL g1384 ( .A(n_281), .B(n_1385), .Y(n_1384) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
INVxp67_ASAP7_75t_L g461 ( .A(n_283), .Y(n_461) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g537 ( .A(n_284), .Y(n_537) );
BUFx4f_ASAP7_75t_L g1034 ( .A(n_284), .Y(n_1034) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g389 ( .A(n_286), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_286), .Y(n_397) );
INVx2_ASAP7_75t_L g412 ( .A(n_286), .Y(n_412) );
AND2x2_ASAP7_75t_L g420 ( .A(n_286), .B(n_287), .Y(n_420) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_427), .Y(n_426) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_286), .B(n_287), .Y(n_525) );
INVx1_ASAP7_75t_L g390 ( .A(n_287), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_287), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g427 ( .A(n_287), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_287), .B(n_412), .Y(n_449) );
BUFx2_ASAP7_75t_L g465 ( .A(n_287), .Y(n_465) );
OR2x2_ASAP7_75t_L g530 ( .A(n_287), .B(n_389), .Y(n_530) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_993), .B1(n_994), .B2(n_1121), .Y(n_291) );
INVx1_ASAP7_75t_L g1121 ( .A(n_292), .Y(n_1121) );
XNOR2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_669), .Y(n_292) );
XOR2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_474), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_378), .C(n_406), .Y(n_297) );
NOR3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_360), .C(n_376), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_323), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_315), .B2(n_316), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_301), .A2(n_315), .B1(n_463), .B2(n_467), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_302), .A2(n_316), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_307), .Y(n_302) );
NAND2x1_ASAP7_75t_L g481 ( .A(n_303), .B(n_307), .Y(n_481) );
AND2x4_ASAP7_75t_SL g796 ( .A(n_303), .B(n_307), .Y(n_796) );
AND2x6_ASAP7_75t_L g923 ( .A(n_303), .B(n_310), .Y(n_923) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g347 ( .A(n_305), .B(n_320), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_305), .B(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g333 ( .A(n_306), .Y(n_333) );
AND2x4_ASAP7_75t_L g339 ( .A(n_306), .B(n_321), .Y(n_339) );
OR2x2_ASAP7_75t_L g364 ( .A(n_306), .B(n_335), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_306), .B(n_322), .Y(n_384) );
AND2x4_ASAP7_75t_L g316 ( .A(n_307), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g377 ( .A(n_307), .B(n_338), .Y(n_377) );
AND2x4_ASAP7_75t_SL g705 ( .A(n_307), .B(n_317), .Y(n_705) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
OR2x2_ASAP7_75t_L g385 ( .A(n_308), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g882 ( .A(n_308), .Y(n_882) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_309), .B(n_413), .Y(n_887) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_310), .B(n_332), .Y(n_404) );
AND2x2_ASAP7_75t_L g925 ( .A(n_310), .B(n_319), .Y(n_925) );
INVx1_ASAP7_75t_L g928 ( .A(n_310), .Y(n_928) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
NAND3x1_ASAP7_75t_L g354 ( .A(n_311), .B(n_355), .C(n_356), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g806 ( .A(n_311), .B(n_356), .Y(n_806) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx3_ASAP7_75t_L g326 ( .A(n_312), .Y(n_326) );
NAND2xp33_ASAP7_75t_SL g684 ( .A(n_312), .B(n_314), .Y(n_684) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND3x4_ASAP7_75t_L g325 ( .A(n_314), .B(n_326), .C(n_327), .Y(n_325) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_316), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_316), .A2(n_480), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_316), .A2(n_480), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_316), .A2(n_480), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
AOI33xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_329), .A3(n_340), .B1(n_348), .B2(n_352), .B3(n_357), .Y(n_323) );
AOI33xp33_ASAP7_75t_L g487 ( .A1(n_324), .A2(n_488), .A3(n_491), .B1(n_496), .B2(n_497), .B3(n_500), .Y(n_487) );
AOI33xp33_ASAP7_75t_L g1004 ( .A1(n_324), .A2(n_1005), .A3(n_1006), .B1(n_1010), .B2(n_1011), .B3(n_1012), .Y(n_1004) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI33xp33_ASAP7_75t_L g562 ( .A1(n_325), .A2(n_352), .A3(n_563), .B1(n_565), .B2(n_571), .B3(n_572), .Y(n_562) );
AOI33xp33_ASAP7_75t_L g619 ( .A1(n_325), .A2(n_500), .A3(n_620), .B1(n_623), .B2(n_627), .B3(n_628), .Y(n_619) );
AOI33xp33_ASAP7_75t_L g798 ( .A1(n_325), .A2(n_799), .A3(n_801), .B1(n_803), .B2(n_804), .B3(n_807), .Y(n_798) );
AOI33xp33_ASAP7_75t_L g840 ( .A1(n_325), .A2(n_804), .A3(n_841), .B1(n_842), .B2(n_843), .B3(n_844), .Y(n_840) );
AOI33xp33_ASAP7_75t_L g1050 ( .A1(n_325), .A2(n_500), .A3(n_1051), .B1(n_1054), .B2(n_1056), .B3(n_1057), .Y(n_1050) );
AOI33xp33_ASAP7_75t_L g1112 ( .A1(n_325), .A2(n_804), .A3(n_1113), .B1(n_1114), .B2(n_1115), .B3(n_1117), .Y(n_1112) );
AOI33xp33_ASAP7_75t_L g1345 ( .A1(n_325), .A2(n_1346), .A3(n_1348), .B1(n_1349), .B2(n_1351), .B3(n_1352), .Y(n_1345) );
INVx1_ASAP7_75t_L g473 ( .A(n_327), .Y(n_473) );
INVx2_ASAP7_75t_SL g544 ( .A(n_327), .Y(n_544) );
OAI31xp33_ASAP7_75t_SL g947 ( .A1(n_327), .A2(n_948), .A3(n_949), .B(n_953), .Y(n_947) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g663 ( .A(n_328), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_328), .B(n_387), .Y(n_866) );
AND2x4_ASAP7_75t_L g548 ( .A(n_330), .B(n_374), .Y(n_548) );
AND2x4_ASAP7_75t_L g1377 ( .A(n_330), .B(n_374), .Y(n_1377) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g489 ( .A(n_331), .Y(n_489) );
INVx8_ASAP7_75t_L g499 ( .A(n_331), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_331), .Y(n_959) );
INVx8_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
BUFx3_ASAP7_75t_L g910 ( .A(n_332), .Y(n_910) );
AND2x2_ASAP7_75t_L g913 ( .A(n_332), .B(n_914), .Y(n_913) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x4_ASAP7_75t_L g344 ( .A(n_333), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g359 ( .A(n_339), .Y(n_359) );
INVx2_ASAP7_75t_L g495 ( .A(n_339), .Y(n_495) );
BUFx3_ASAP7_75t_L g564 ( .A(n_339), .Y(n_564) );
BUFx2_ASAP7_75t_L g573 ( .A(n_339), .Y(n_573) );
BUFx2_ASAP7_75t_L g693 ( .A(n_339), .Y(n_693) );
AND2x2_ASAP7_75t_L g916 ( .A(n_339), .B(n_914), .Y(n_916) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_343), .A2(n_686), .B1(n_687), .B2(n_691), .C(n_692), .Y(n_685) );
INVx3_ASAP7_75t_L g802 ( .A(n_343), .Y(n_802) );
INVx1_ASAP7_75t_L g902 ( .A(n_343), .Y(n_902) );
OR2x6_ASAP7_75t_SL g930 ( .A(n_343), .B(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_343), .Y(n_1008) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_344), .Y(n_351) );
BUFx8_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_344), .Y(n_568) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx12f_ASAP7_75t_L g490 ( .A(n_347), .Y(n_490) );
INVx5_ASAP7_75t_L g570 ( .A(n_347), .Y(n_570) );
BUFx2_ASAP7_75t_L g626 ( .A(n_347), .Y(n_626) );
AND2x4_ASAP7_75t_L g934 ( .A(n_347), .B(n_932), .Y(n_934) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_347), .Y(n_1055) );
INVx8_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g493 ( .A(n_350), .Y(n_493) );
INVx5_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_SL g625 ( .A(n_351), .Y(n_625) );
INVx3_ASAP7_75t_L g906 ( .A(n_351), .Y(n_906) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g500 ( .A(n_353), .Y(n_500) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g695 ( .A(n_354), .Y(n_695) );
INVx2_ASAP7_75t_SL g622 ( .A(n_358), .Y(n_622) );
BUFx3_ASAP7_75t_L g800 ( .A(n_358), .Y(n_800) );
INVx1_ASAP7_75t_L g1053 ( .A(n_358), .Y(n_1053) );
OR2x6_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
OR2x2_ASAP7_75t_L g575 ( .A(n_362), .B(n_365), .Y(n_575) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g810 ( .A(n_366), .B(n_802), .Y(n_810) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g374 ( .A(n_367), .Y(n_374) );
OR2x2_ASAP7_75t_L g381 ( .A(n_367), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g399 ( .A(n_367), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
OR2x2_ASAP7_75t_L g683 ( .A(n_368), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_SL g862 ( .A(n_368), .B(n_429), .Y(n_862) );
INVx1_ASAP7_75t_L g983 ( .A(n_368), .Y(n_983) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g914 ( .A(n_371), .Y(n_914) );
INVx1_ASAP7_75t_L g932 ( .A(n_371), .Y(n_932) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_373), .A2(n_517), .B1(n_519), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_373), .A2(n_548), .B1(n_714), .B2(n_715), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_373), .A2(n_548), .B1(n_736), .B2(n_737), .Y(n_764) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx2_ASAP7_75t_SL g751 ( .A(n_375), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_376), .B(n_681), .C(n_703), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g836 ( .A(n_376), .B(n_837), .C(n_845), .Y(n_836) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g501 ( .A(n_377), .Y(n_501) );
INVx3_ASAP7_75t_L g577 ( .A(n_377), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_377), .B(n_748), .C(n_760), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g793 ( .A(n_377), .B(n_794), .C(n_808), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g1108 ( .A1(n_377), .A2(n_1100), .B(n_1109), .C(n_1110), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_391), .B(n_392), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_379), .B(n_550), .Y(n_549) );
AOI21xp33_ASAP7_75t_SL g578 ( .A1(n_379), .A2(n_579), .B(n_580), .Y(n_578) );
NAND2xp33_ASAP7_75t_L g629 ( .A(n_379), .B(n_630), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_379), .A2(n_677), .B(n_678), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_379), .A2(n_762), .B(n_763), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_379), .A2(n_791), .B(n_792), .Y(n_790) );
AOI21xp33_ASAP7_75t_L g833 ( .A1(n_379), .A2(n_834), .B(n_835), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_379), .A2(n_1016), .B(n_1017), .Y(n_1015) );
AOI21xp33_ASAP7_75t_SL g1059 ( .A1(n_379), .A2(n_1060), .B(n_1061), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_379), .B(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_379), .B(n_1379), .Y(n_1378) );
INVx8_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_385), .Y(n_380) );
BUFx3_ASAP7_75t_L g956 ( .A(n_382), .Y(n_956) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_383), .Y(n_700) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g690 ( .A(n_384), .Y(n_690) );
INVx1_ASAP7_75t_L g883 ( .A(n_386), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_387), .B(n_396), .Y(n_395) );
AND2x6_ASAP7_75t_L g435 ( .A(n_387), .B(n_419), .Y(n_435) );
INVx1_ASAP7_75t_L g466 ( .A(n_387), .Y(n_466) );
AND2x2_ASAP7_75t_L g772 ( .A(n_387), .B(n_773), .Y(n_772) );
INVx3_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
AND2x2_ASAP7_75t_L g440 ( .A(n_388), .B(n_413), .Y(n_440) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_388), .Y(n_513) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_393), .Y(n_546) );
INVx2_ASAP7_75t_L g635 ( .A(n_393), .Y(n_635) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
AND2x4_ASAP7_75t_L g679 ( .A(n_394), .B(n_399), .Y(n_679) );
INVx2_ASAP7_75t_SL g987 ( .A(n_394), .Y(n_987) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .Y(n_394) );
OR2x2_ASAP7_75t_L g869 ( .A(n_395), .B(n_398), .Y(n_869) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g405 ( .A(n_398), .Y(n_405) );
INVx1_ASAP7_75t_L g898 ( .A(n_398), .Y(n_898) );
INVx3_ASAP7_75t_L g967 ( .A(n_400), .Y(n_967) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g927 ( .A(n_401), .Y(n_927) );
INVx5_ASAP7_75t_L g486 ( .A(n_403), .Y(n_486) );
INVx3_ASAP7_75t_L g1109 ( .A(n_403), .Y(n_1109) );
OR2x6_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g581 ( .A(n_404), .B(n_405), .Y(n_581) );
INVx2_ASAP7_75t_L g920 ( .A(n_404), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_445), .B(n_470), .Y(n_406) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g504 ( .A(n_409), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_409), .B(n_1344), .Y(n_1364) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g515 ( .A(n_410), .Y(n_515) );
BUFx2_ASAP7_75t_L g587 ( .A(n_410), .Y(n_587) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
INVx2_ASAP7_75t_L g659 ( .A(n_411), .Y(n_659) );
BUFx3_ASAP7_75t_L g734 ( .A(n_411), .Y(n_734) );
AND2x4_ASAP7_75t_L g444 ( .A(n_413), .B(n_425), .Y(n_444) );
AND2x4_ASAP7_75t_SL g469 ( .A(n_413), .B(n_419), .Y(n_469) );
AND2x2_ASAP7_75t_L g938 ( .A(n_413), .B(n_425), .Y(n_938) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_413), .B(n_888), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_430), .B(n_435), .Y(n_415) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g1023 ( .A(n_418), .Y(n_1023) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g507 ( .A(n_419), .Y(n_507) );
BUFx3_ASAP7_75t_L g589 ( .A(n_419), .Y(n_589) );
BUFx3_ASAP7_75t_L g608 ( .A(n_419), .Y(n_608) );
BUFx3_ASAP7_75t_L g730 ( .A(n_419), .Y(n_730) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g591 ( .A(n_424), .Y(n_591) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g732 ( .A(n_425), .Y(n_732) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_425), .Y(n_822) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
BUFx3_ASAP7_75t_L g642 ( .A(n_426), .Y(n_642) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g509 ( .A(n_429), .Y(n_509) );
INVx4_ASAP7_75t_L g592 ( .A(n_429), .Y(n_592) );
AND2x4_ASAP7_75t_L g981 ( .A(n_429), .B(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g586 ( .A(n_432), .Y(n_586) );
INVx2_ASAP7_75t_SL g721 ( .A(n_432), .Y(n_721) );
INVx1_ASAP7_75t_L g780 ( .A(n_432), .Y(n_780) );
INVx1_ASAP7_75t_L g1360 ( .A(n_432), .Y(n_1360) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g1073 ( .A(n_434), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_435), .A2(n_506), .B(n_510), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_435), .A2(n_585), .B(n_588), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_435), .A2(n_641), .B(n_643), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_435), .A2(n_709), .B(n_710), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_435), .A2(n_729), .B(n_733), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_435), .A2(n_783), .B(n_785), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_435), .A2(n_827), .B(n_829), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_435), .A2(n_1021), .B(n_1025), .Y(n_1020) );
AOI21xp5_ASAP7_75t_L g1070 ( .A1(n_435), .A2(n_1071), .B(n_1074), .Y(n_1070) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_435), .A2(n_1099), .B1(n_1100), .B2(n_1101), .C(n_1102), .Y(n_1098) );
INVx1_ASAP7_75t_L g1365 ( .A(n_435), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_441), .B2(n_442), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_438), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_438), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_438), .A2(n_596), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_438), .A2(n_596), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_440), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_440), .A2(n_444), .B1(n_736), .B2(n_737), .Y(n_735) );
AND2x4_ASAP7_75t_L g897 ( .A(n_440), .B(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_442), .A2(n_1027), .B1(n_1028), .B2(n_1029), .Y(n_1026) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_444), .Y(n_518) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_444), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_444), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_444), .A2(n_646), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_444), .A2(n_646), .B1(n_1104), .B2(n_1105), .Y(n_1103) );
AOI22xp5_ASAP7_75t_L g1361 ( .A1(n_444), .A2(n_646), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVx5_ASAP7_75t_L g1066 ( .A(n_446), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g540 ( .A(n_447), .Y(n_540) );
INVx2_ASAP7_75t_SL g603 ( .A(n_447), .Y(n_603) );
INVx2_ASAP7_75t_L g976 ( .A(n_447), .Y(n_976) );
INVx1_ASAP7_75t_L g1036 ( .A(n_447), .Y(n_1036) );
INVx8_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g874 ( .A(n_448), .Y(n_874) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g1039 ( .A(n_453), .Y(n_1039) );
INVx1_ASAP7_75t_L g1096 ( .A(n_453), .Y(n_1096) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g1077 ( .A(n_454), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g607 ( .A(n_456), .Y(n_607) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
INVx1_ASAP7_75t_L g744 ( .A(n_459), .Y(n_744) );
INVx3_ASAP7_75t_L g823 ( .A(n_459), .Y(n_823) );
INVx1_ASAP7_75t_L g1373 ( .A(n_461), .Y(n_1373) );
INVx2_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
INVx2_ASAP7_75t_L g599 ( .A(n_463), .Y(n_599) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g773 ( .A(n_465), .Y(n_773) );
INVx1_ASAP7_75t_L g868 ( .A(n_465), .Y(n_868) );
INVx2_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
INVx2_ASAP7_75t_L g598 ( .A(n_467), .Y(n_598) );
INVx4_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g1093 ( .A(n_469), .Y(n_1093) );
OAI21xp5_ASAP7_75t_L g1018 ( .A1(n_470), .A2(n_1019), .B(n_1030), .Y(n_1018) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g899 ( .A1(n_472), .A2(n_900), .B(n_917), .C(n_935), .Y(n_899) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g746 ( .A(n_473), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_552), .B1(n_553), .B2(n_668), .Y(n_474) );
INVx1_ASAP7_75t_L g668 ( .A(n_475), .Y(n_668) );
XOR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_551), .Y(n_475) );
NAND3x1_ASAP7_75t_SL g476 ( .A(n_477), .B(n_502), .C(n_549), .Y(n_476) );
AND4x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_484), .C(n_487), .D(n_501), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_482), .B2(n_483), .Y(n_478) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_486), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_486), .B(n_1344), .Y(n_1343) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_490), .Y(n_1009) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g759 ( .A(n_495), .Y(n_759) );
INVx2_ASAP7_75t_L g1118 ( .A(n_495), .Y(n_1118) );
INVx1_ASAP7_75t_L g1347 ( .A(n_495), .Y(n_1347) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_501), .Y(n_1014) );
O2A1O1Ixp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_520), .B(n_544), .C(n_545), .Y(n_502) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g712 ( .A(n_513), .Y(n_712) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_526), .B1(n_527), .B2(n_531), .C(n_532), .Y(n_522) );
BUFx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g742 ( .A(n_524), .Y(n_742) );
OR2x2_ASAP7_75t_L g891 ( .A(n_524), .B(n_887), .Y(n_891) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_525), .Y(n_653) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g858 ( .A(n_530), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g1367 ( .A1(n_532), .A2(n_858), .B1(n_1368), .B2(n_1369), .C(n_1370), .Y(n_1367) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_538), .B2(n_541), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_536), .A2(n_601), .B1(n_602), .B2(n_604), .C(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g855 ( .A(n_536), .Y(n_855) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_537), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
OAI22x1_ASAP7_75t_SL g979 ( .A1(n_537), .A2(n_957), .B1(n_976), .B2(n_980), .Y(n_979) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g854 ( .A(n_539), .Y(n_854) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_544), .A2(n_583), .B(n_597), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g1062 ( .A1(n_544), .A2(n_1063), .B(n_1069), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_548), .A2(n_810), .B1(n_1104), .B2(n_1105), .Y(n_1107) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_609), .B2(n_667), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_578), .C(n_582), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_574), .C(n_576), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g697 ( .A(n_568), .Y(n_697) );
INVx2_ASAP7_75t_R g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g1350 ( .A(n_570), .Y(n_1350) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND4xp25_ASAP7_75t_SL g613 ( .A(n_577), .B(n_614), .C(n_617), .D(n_619), .Y(n_613) );
AND4x1_ASAP7_75t_L g1339 ( .A(n_577), .B(n_1340), .C(n_1343), .D(n_1345), .Y(n_1339) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_596), .A2(n_646), .B1(n_831), .B2(n_832), .Y(n_830) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g667 ( .A(n_609), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_610), .B(n_631), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_629), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_SL g664 ( .A(n_613), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_629), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_638), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_637), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_648), .B(n_660), .Y(n_638) );
INVx1_ASAP7_75t_L g656 ( .A(n_642), .Y(n_656) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_642), .Y(n_784) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_642), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_646), .Y(n_1028) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_654), .C(n_657), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g718 ( .A(n_652), .Y(n_718) );
INVx2_ASAP7_75t_L g1368 ( .A(n_652), .Y(n_1368) );
INVx4_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx4f_ASAP7_75t_L g777 ( .A(n_653), .Y(n_777) );
BUFx4f_ASAP7_75t_L g860 ( .A(n_653), .Y(n_860) );
OR2x6_ASAP7_75t_L g870 ( .A(n_653), .B(n_871), .Y(n_870) );
BUFx4f_ASAP7_75t_L g1357 ( .A(n_653), .Y(n_1357) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g828 ( .A(n_656), .Y(n_828) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g888 ( .A(n_659), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_660), .A2(n_707), .B(n_716), .Y(n_706) );
OAI21xp5_ASAP7_75t_SL g769 ( .A1(n_660), .A2(n_770), .B(n_781), .Y(n_769) );
OAI21xp5_ASAP7_75t_SL g815 ( .A1(n_660), .A2(n_816), .B(n_825), .Y(n_815) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g1089 ( .A(n_661), .Y(n_1089) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x6_ASAP7_75t_L g805 ( .A(n_663), .B(n_806), .Y(n_805) );
AND2x4_ASAP7_75t_L g878 ( .A(n_663), .B(n_879), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_847), .B1(n_991), .B2(n_992), .Y(n_669) );
INVx2_ASAP7_75t_L g992 ( .A(n_670), .Y(n_992) );
AOI22x1_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_766), .B2(n_846), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AO22x2_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_723), .B1(n_724), .B2(n_765), .Y(n_673) );
INVx1_ASAP7_75t_L g765 ( .A(n_674), .Y(n_765) );
AND4x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_680), .C(n_706), .D(n_722), .Y(n_675) );
OAI22xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_685), .B1(n_694), .B2(n_696), .Y(n_681) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx8_ASAP7_75t_L g749 ( .A(n_683), .Y(n_749) );
BUFx2_ASAP7_75t_L g907 ( .A(n_684), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_687), .A2(n_751), .B1(n_752), .B2(n_753), .C(n_754), .Y(n_750) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_695), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_699), .B2(n_701), .C(n_702), .Y(n_696) );
INVx1_ASAP7_75t_L g1116 ( .A(n_697), .Y(n_1116) );
OAI211xp5_ASAP7_75t_L g717 ( .A1(n_698), .A2(n_718), .B(n_719), .C(n_720), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_699), .A2(n_740), .B1(n_751), .B2(n_757), .C(n_758), .Y(n_756) );
CKINVDCx8_ASAP7_75t_R g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_705), .A2(n_774), .B1(n_796), .B2(n_797), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_705), .A2(n_796), .B1(n_818), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_705), .A2(n_796), .B1(n_1092), .B2(n_1094), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1340 ( .A1(n_705), .A2(n_796), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g786 ( .A(n_712), .Y(n_786) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND4x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_747), .C(n_761), .D(n_764), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_738), .B(n_746), .Y(n_726) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_743), .C(n_745), .Y(n_739) );
INVx5_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
O2A1O1Ixp5_ASAP7_75t_SL g1353 ( .A1(n_746), .A2(n_1354), .B(n_1366), .C(n_1375), .Y(n_1353) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_749), .A2(n_750), .B1(n_755), .B2(n_756), .Y(n_748) );
INVx1_ASAP7_75t_L g1011 ( .A(n_755), .Y(n_1011) );
INVx1_ASAP7_75t_L g846 ( .A(n_766), .Y(n_846) );
XNOR2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_813), .Y(n_766) );
INVx1_ASAP7_75t_L g812 ( .A(n_768), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_790), .C(n_793), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_772), .B(n_818), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g1091 ( .A1(n_772), .A2(n_1092), .B1(n_1093), .B2(n_1094), .C1(n_1095), .C2(n_1097), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_778), .C(n_779), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g819 ( .A1(n_777), .A2(n_820), .B(n_821), .C(n_824), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .Y(n_794) );
INVx1_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g1352 ( .A(n_805), .Y(n_1352) );
INVx3_ASAP7_75t_L g961 ( .A(n_806), .Y(n_961) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_810), .A2(n_1362), .B1(n_1363), .B2(n_1377), .Y(n_1376) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_833), .C(n_836), .Y(n_814) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_822), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .Y(n_837) );
INVx1_ASAP7_75t_L g991 ( .A(n_847), .Y(n_991) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
XNOR2x1_ASAP7_75t_L g848 ( .A(n_849), .B(n_940), .Y(n_848) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_939), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_899), .Y(n_850) );
NAND3xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_880), .C(n_893), .Y(n_851) );
AOI211xp5_ASAP7_75t_SL g852 ( .A1(n_853), .A2(n_856), .B(n_863), .C(n_872), .Y(n_852) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_858), .A2(n_860), .B1(n_876), .B2(n_877), .C(n_878), .Y(n_875) );
INVxp67_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g986 ( .A(n_864), .Y(n_986) );
NAND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g871 ( .A(n_865), .Y(n_871) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_870), .Y(n_990) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_878), .Y(n_977) );
AOI222xp33_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_884), .B1(n_885), .B2(n_889), .C1(n_890), .C2(n_892), .Y(n_880) );
AOI21xp33_ASAP7_75t_SL g988 ( .A1(n_881), .A2(n_989), .B(n_990), .Y(n_988) );
AND2x4_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
AOI222xp33_ASAP7_75t_L g984 ( .A1(n_885), .A2(n_951), .B1(n_963), .B2(n_985), .C1(n_986), .C2(n_987), .Y(n_984) );
AND2x4_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI211xp5_ASAP7_75t_L g917 ( .A1(n_889), .A2(n_918), .B(n_921), .C(n_929), .Y(n_917) );
AOI222xp33_ASAP7_75t_L g971 ( .A1(n_890), .A2(n_952), .B1(n_972), .B2(n_977), .C1(n_978), .C2(n_981), .Y(n_971) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_897), .Y(n_942) );
AND2x4_ASAP7_75t_L g937 ( .A(n_898), .B(n_938), .Y(n_937) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_903), .B1(n_904), .B2(n_908), .C(n_911), .Y(n_900) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_906), .A2(n_955), .B1(n_956), .B2(n_957), .C(n_958), .Y(n_954) );
BUFx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_913), .A2(n_916), .B1(n_943), .B2(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx4_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_923), .A2(n_925), .B1(n_951), .B2(n_952), .Y(n_950) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OR2x6_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx3_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_937), .B(n_946), .Y(n_945) );
AOI211x1_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_943), .B(n_944), .C(n_970), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_947), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_962), .C(n_964), .Y(n_953) );
INVx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_966), .B(n_968), .C(n_969), .Y(n_964) );
INVx3_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_984), .C(n_988), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_976), .A2(n_1372), .B1(n_1373), .B2(n_1374), .Y(n_1371) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_996), .B1(n_1041), .B2(n_1042), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx2_ASAP7_75t_SL g996 ( .A(n_997), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1015), .C(n_1018), .Y(n_998) );
NOR3xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1013), .C(n_1014), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .Y(n_1000) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
NOR3xp33_ASAP7_75t_L g1045 ( .A(n_1014), .B(n_1046), .C(n_1058), .Y(n_1045) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1035), .B1(n_1036), .B2(n_1037), .C(n_1038), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1064 ( .A1(n_1032), .A2(n_1065), .B1(n_1066), .B2(n_1067), .C(n_1068), .Y(n_1064) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
BUFx6f_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1081), .B1(n_1082), .B2(n_1120), .Y(n_1042) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1043), .Y(n_1120) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1059), .C(n_1062), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1050), .Y(n_1046) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_SL g1072 ( .A(n_1073), .Y(n_1072) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .C(n_1108), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1090), .B(n_1106), .Y(n_1088) );
NAND3xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1098), .C(n_1103), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1332), .B1(n_1335), .B2(n_1381), .C(n_1386), .Y(n_1122) );
AND4x1_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1250), .C(n_1280), .D(n_1309), .Y(n_1123) );
AOI211xp5_ASAP7_75t_L g1124 ( .A1(n_1125), .A2(n_1192), .B(n_1196), .C(n_1235), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
A2O1A1Ixp33_ASAP7_75t_L g1263 ( .A1(n_1126), .A2(n_1221), .B(n_1225), .C(n_1264), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1180), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1174), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1151), .B1(n_1164), .B2(n_1167), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1129), .B(n_1175), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1129), .B(n_1153), .Y(n_1274) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1146), .Y(n_1130) );
OAI32xp33_ASAP7_75t_L g1203 ( .A1(n_1131), .A2(n_1204), .A3(n_1206), .B1(n_1211), .B2(n_1213), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1131), .B(n_1153), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1131), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1131), .Y(n_1307) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1132), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1132), .B(n_1153), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1132), .B(n_1147), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1132), .B(n_1146), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1140), .Y(n_1132) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1134), .Y(n_1334) );
AND2x6_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1135), .B(n_1139), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_1135), .B(n_1142), .Y(n_1141) );
AND2x6_ASAP7_75t_L g1144 ( .A(n_1135), .B(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1135), .B(n_1139), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1135), .B(n_1139), .Y(n_1209) );
OAI21xp5_ASAP7_75t_L g1397 ( .A1(n_1136), .A2(n_1398), .B(n_1399), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1137), .B(n_1143), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1146), .B(n_1192), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1146), .B(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1146), .B(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1146), .B(n_1193), .Y(n_1271) );
OAI32xp33_ASAP7_75t_L g1285 ( .A1(n_1146), .A2(n_1147), .A3(n_1218), .B1(n_1286), .B2(n_1288), .Y(n_1285) );
HB1xp67_ASAP7_75t_SL g1310 ( .A(n_1146), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_1147), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1147), .B(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1147), .B(n_1230), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1147), .B(n_1193), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1147), .B(n_1154), .Y(n_1319) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1150), .Y(n_1147) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1152), .B(n_1189), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1157), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1153), .B(n_1214), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1153), .B(n_1189), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1153), .B(n_1219), .Y(n_1292) );
CKINVDCx14_ASAP7_75t_R g1299 ( .A(n_1153), .Y(n_1299) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_1154), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1154), .B(n_1171), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1154), .B(n_1157), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1154), .B(n_1276), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1154), .B(n_1186), .Y(n_1284) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1154), .B(n_1177), .Y(n_1296) );
AND2x4_ASAP7_75t_SL g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1157), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1157), .B(n_1189), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1157), .B(n_1179), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1157), .B(n_1292), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1161), .Y(n_1157) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1158), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1158), .B(n_1178), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1158), .B(n_1189), .Y(n_1188) );
NOR2xp33_ASAP7_75t_L g1216 ( .A(n_1158), .B(n_1217), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1158), .B(n_1171), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1158), .B(n_1171), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1161), .Y(n_1178) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1161), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1161), .B(n_1189), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1161), .B(n_1170), .Y(n_1241) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1161), .Y(n_1273) );
NAND2x1_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1163), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1164), .B(n_1230), .Y(n_1249) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1165), .B(n_1168), .Y(n_1191) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1165), .Y(n_1294) );
OAI21xp33_ASAP7_75t_L g1181 ( .A1(n_1166), .A2(n_1182), .B(n_1185), .Y(n_1181) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1166), .Y(n_1199) );
OAI21xp5_ASAP7_75t_L g1293 ( .A1(n_1167), .A2(n_1182), .B(n_1294), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1168), .B(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1168), .B(n_1186), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1168), .B(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1168), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1168), .B(n_1306), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1168), .B(n_1297), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1170), .B(n_1184), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1171), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1171), .B(n_1186), .Y(n_1185) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1171), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1171), .B(n_1202), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1171), .B(n_1284), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1171), .B(n_1241), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1175), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1179), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1176), .B(n_1189), .Y(n_1214) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1177), .B(n_1189), .Y(n_1282) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1179), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1179), .B(n_1186), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1187), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_1182), .A2(n_1185), .B1(n_1200), .B2(n_1237), .C(n_1238), .Y(n_1236) );
NOR2xp33_ASAP7_75t_SL g1318 ( .A(n_1183), .B(n_1214), .Y(n_1318) );
OAI21xp5_ASAP7_75t_L g1187 ( .A1(n_1186), .A2(n_1188), .B(n_1190), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1186), .B(n_1259), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1186), .A2(n_1217), .B1(n_1241), .B2(n_1269), .C(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1186), .Y(n_1331) );
A2O1A1Ixp33_ASAP7_75t_L g1243 ( .A1(n_1188), .A2(n_1244), .B(n_1245), .C(n_1246), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1189), .B(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1189), .B(n_1273), .Y(n_1327) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
AOI21xp33_ASAP7_75t_L g1329 ( .A1(n_1191), .A2(n_1330), .B(n_1331), .Y(n_1329) );
OAI221xp5_ASAP7_75t_L g1322 ( .A1(n_1192), .A2(n_1228), .B1(n_1283), .B2(n_1323), .C(n_1326), .Y(n_1322) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1193), .B(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1193), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1195), .Y(n_1193) );
NAND4xp25_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1215), .C(n_1223), .D(n_1226), .Y(n_1196) );
O2A1O1Ixp33_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1200), .B(n_1201), .C(n_1203), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1199), .B(n_1230), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1199), .B(n_1266), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1199), .B(n_1287), .Y(n_1314) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1200), .Y(n_1256) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1205), .Y(n_1306) );
INVxp67_ASAP7_75t_SL g1308 ( .A(n_1206), .Y(n_1308) );
INVx3_ASAP7_75t_L g1222 ( .A(n_1207), .Y(n_1222) );
NAND3xp33_ASAP7_75t_SL g1265 ( .A(n_1207), .B(n_1225), .C(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1207), .B(n_1230), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1210), .Y(n_1207) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1212), .Y(n_1269) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OAI211xp5_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1218), .B(n_1219), .C(n_1221), .Y(n_1215) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
A2O1A1Ixp33_ASAP7_75t_L g1257 ( .A1(n_1220), .A2(n_1221), .B(n_1258), .C(n_1261), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_L g1281 ( .A1(n_1220), .A2(n_1282), .B(n_1283), .C(n_1285), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1220), .B(n_1301), .Y(n_1321) );
AOI21xp33_ASAP7_75t_L g1295 ( .A1(n_1221), .A2(n_1296), .B(n_1297), .Y(n_1295) );
CKINVDCx14_ASAP7_75t_R g1221 ( .A(n_1222), .Y(n_1221) );
AOI31xp33_ASAP7_75t_L g1235 ( .A1(n_1222), .A2(n_1236), .A3(n_1243), .B(n_1247), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1222), .B(n_1229), .Y(n_1262) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1222), .A2(n_1304), .B(n_1307), .Y(n_1303) );
A2O1A1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1222), .A2(n_1327), .B(n_1328), .C(n_1329), .Y(n_1326) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1232), .Y(n_1226) );
A2O1A1Ixp33_ASAP7_75t_L g1250 ( .A1(n_1227), .A2(n_1251), .B(n_1253), .C(n_1263), .Y(n_1250) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1231), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
NAND3xp33_ASAP7_75t_L g1239 ( .A(n_1230), .B(n_1240), .C(n_1242), .Y(n_1239) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1230), .Y(n_1266) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1231), .Y(n_1297) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_1233), .A2(n_1254), .B1(n_1255), .B2(n_1256), .C(n_1257), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1234), .B(n_1260), .Y(n_1317) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1248 ( .A(n_1241), .B(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1245), .Y(n_1330) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1246), .Y(n_1255) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1252), .B(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
CKINVDCx14_ASAP7_75t_R g1261 ( .A(n_1262), .Y(n_1261) );
A2O1A1O1Ixp25_ASAP7_75t_L g1309 ( .A1(n_1262), .A2(n_1310), .B(n_1311), .C(n_1312), .D(n_1322), .Y(n_1309) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1267), .B1(n_1268), .B2(n_1271), .C(n_1272), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1280 ( .A1(n_1266), .A2(n_1281), .B(n_1290), .Y(n_1280) );
O2A1O1Ixp33_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1274), .B(n_1275), .C(n_1277), .Y(n_1272) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1274), .Y(n_1328) );
NOR2xp33_ASAP7_75t_SL g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1288), .Y(n_1302) );
AOI331xp33_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1293), .A3(n_1295), .B1(n_1298), .B2(n_1302), .B3(n_1303), .C1(n_1308), .Y(n_1290) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1298), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1300), .Y(n_1298) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
NOR2xp33_ASAP7_75t_SL g1315 ( .A(n_1307), .B(n_1316), .Y(n_1315) );
OAI221xp5_ASAP7_75t_L g1312 ( .A1(n_1313), .A2(n_1315), .B1(n_1318), .B2(n_1319), .C(n_1320), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVxp67_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
CKINVDCx20_ASAP7_75t_R g1332 ( .A(n_1333), .Y(n_1332) );
CKINVDCx20_ASAP7_75t_R g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
XOR2xp5_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1380), .Y(n_1337) );
HB1xp67_ASAP7_75t_L g1395 ( .A(n_1338), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1353), .C(n_1378), .Y(n_1338) );
NAND4xp25_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1361), .C(n_1364), .D(n_1365), .Y(n_1354) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B(n_1358), .C(n_1359), .Y(n_1355) );
CKINVDCx20_ASAP7_75t_R g1381 ( .A(n_1382), .Y(n_1381) );
CKINVDCx20_ASAP7_75t_R g1382 ( .A(n_1383), .Y(n_1382) );
INVx3_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVxp33_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
HB1xp67_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
endmodule