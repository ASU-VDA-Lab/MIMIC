module fake_netlist_5_1112_n_1701 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1701);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1701;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_79),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_50),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_14),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_28),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_77),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_18),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_13),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_23),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_104),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_59),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_29),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_40),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_69),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_50),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_147),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_37),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_62),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_22),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_38),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_2),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_8),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_47),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_115),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_11),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_56),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_43),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_94),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_81),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_83),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_143),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_27),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_70),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_25),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_101),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_54),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_87),
.Y(n_260)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_14),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_8),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_71),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_66),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_84),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_40),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_64),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_96),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_138),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_24),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_121),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_49),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_114),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_27),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_42),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_43),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_41),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_95),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_86),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_56),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_36),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_24),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_33),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_12),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_110),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_15),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_55),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_156),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_158),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_163),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_225),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_200),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_257),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_205),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_247),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_183),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_155),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_160),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_162),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_238),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_240),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_260),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_170),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_171),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_173),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_181),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_217),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_209),
.B(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_182),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_188),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_159),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_177),
.B(n_0),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_191),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_193),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_196),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_217),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_159),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_177),
.B(n_1),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_202),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_1),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_209),
.B(n_3),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_215),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_257),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_239),
.B(n_4),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_216),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_220),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_158),
.B(n_4),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_239),
.B(n_5),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_243),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_224),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_236),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_157),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_241),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_242),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_253),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_183),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_186),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_259),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_165),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_169),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_283),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_265),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_329),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_198),
.C(n_186),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_357),
.A2(n_273),
.B(n_263),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_272),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_308),
.B(n_180),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_184),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_184),
.Y(n_406)
);

AND3x1_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_201),
.C(n_198),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

OR2x6_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_229),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_320),
.B(n_219),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_219),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_341),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_321),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_336),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_226),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_322),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_276),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_334),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_353),
.B(n_263),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_371),
.B(n_226),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_335),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_363),
.B(n_273),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_339),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_340),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_347),
.B1(n_336),
.B2(n_306),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_306),
.B1(n_294),
.B2(n_251),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_377),
.B1(n_332),
.B2(n_344),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_418),
.B1(n_424),
.B2(n_413),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_392),
.B(n_164),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_383),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_383),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_345),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_413),
.B1(n_442),
.B2(n_426),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_346),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_164),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_355),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_418),
.B(n_167),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_356),
.B1(n_315),
.B2(n_359),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_425),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_418),
.A2(n_251),
.B1(n_201),
.B2(n_210),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_364),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_404),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_367),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_427),
.B(n_368),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_440),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_404),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_L g482 ( 
.A1(n_413),
.A2(n_356),
.B1(n_315),
.B2(n_359),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_373),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_381),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_348),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_418),
.A2(n_248),
.B1(n_210),
.B2(n_211),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_413),
.A2(n_248),
.B1(n_211),
.B2(n_212),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_374),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_413),
.A2(n_442),
.B1(n_389),
.B2(n_436),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_395),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_427),
.B(n_351),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_403),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_382),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_427),
.B(n_358),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_382),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_407),
.A2(n_369),
.B1(n_365),
.B2(n_360),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_167),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_375),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_L g507 ( 
.A(n_389),
.B(n_301),
.C(n_285),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_442),
.B(n_203),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_403),
.B(n_311),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_442),
.B(n_245),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_394),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

AND3x2_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_284),
.C(n_172),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_425),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_407),
.A2(n_213),
.B1(n_307),
.B2(n_304),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_434),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_427),
.B(n_434),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_168),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_378),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_382),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_442),
.B(n_277),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_401),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_378),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_419),
.B(n_312),
.Y(n_531)
);

BUFx8_ASAP7_75t_SL g532 ( 
.A(n_433),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_387),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_430),
.B(n_230),
.C(n_223),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_387),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_413),
.A2(n_207),
.B1(n_300),
.B2(n_296),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_442),
.B(n_286),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_427),
.B(n_292),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_427),
.B(n_168),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_396),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_427),
.B(n_297),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_423),
.B(n_299),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_396),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_378),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_392),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_385),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_396),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_419),
.B(n_313),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_420),
.B(n_326),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_442),
.B(n_172),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_379),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_379),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_423),
.B(n_214),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_441),
.A2(n_195),
.B1(n_295),
.B2(n_291),
.Y(n_555)
);

BUFx4f_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_415),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_436),
.A2(n_212),
.B1(n_228),
.B2(n_303),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_396),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_396),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_379),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_400),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_400),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_436),
.A2(n_234),
.B1(n_237),
.B2(n_303),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_380),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_433),
.B(n_250),
.C(n_189),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_400),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_385),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_401),
.B(n_174),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_436),
.A2(n_228),
.B1(n_275),
.B2(n_302),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_440),
.B(n_174),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_385),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_406),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_406),
.Y(n_575)
);

BUFx8_ASAP7_75t_SL g576 ( 
.A(n_433),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_420),
.B(n_190),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_435),
.B(n_190),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_423),
.B(n_214),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_380),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_423),
.B(n_214),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_423),
.B(n_316),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_422),
.B(n_324),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_438),
.B(n_192),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_415),
.B(n_192),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_428),
.B(n_421),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_438),
.B(n_175),
.Y(n_587)
);

NOR2x1p5_ASAP7_75t_L g588 ( 
.A(n_429),
.B(n_176),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_556),
.B(n_438),
.Y(n_589)
);

INVxp33_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_451),
.A2(n_438),
.B1(n_422),
.B2(n_431),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_446),
.A2(n_438),
.B1(n_431),
.B2(n_430),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_487),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_517),
.B(n_429),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_496),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_532),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_505),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_556),
.B(n_429),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_506),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_466),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_457),
.B(n_441),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_415),
.Y(n_608)
);

AO221x1_ASAP7_75t_L g609 ( 
.A1(n_465),
.A2(n_275),
.B1(n_234),
.B2(n_237),
.C(n_244),
.Y(n_609)
);

OAI22x1_ASAP7_75t_L g610 ( 
.A1(n_509),
.A2(n_403),
.B1(n_502),
.B2(n_450),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_533),
.A2(n_390),
.B(n_244),
.C(n_289),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_545),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_536),
.B(n_429),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_574),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_556),
.B(n_421),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_575),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_552),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_443),
.B(n_421),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_474),
.A2(n_437),
.B1(n_415),
.B2(n_436),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_546),
.B(n_437),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_474),
.A2(n_437),
.B1(n_436),
.B2(n_421),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_464),
.A2(n_390),
.B1(n_197),
.B2(n_208),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_480),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_529),
.B(n_421),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_456),
.B(n_475),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_490),
.A2(n_390),
.B(n_269),
.C(n_279),
.Y(n_630)
);

AOI221xp5_ASAP7_75t_L g631 ( 
.A1(n_519),
.A2(n_252),
.B1(n_227),
.B2(n_298),
.C(n_294),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_553),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_458),
.B(n_421),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_458),
.B(n_435),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_463),
.B(n_435),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_553),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_455),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_577),
.A2(n_282),
.B(n_269),
.C(n_279),
.Y(n_638)
);

OAI221xp5_ASAP7_75t_L g639 ( 
.A1(n_468),
.A2(n_282),
.B1(n_287),
.B2(n_289),
.C(n_298),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_479),
.A2(n_287),
.B(n_302),
.C(n_246),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_483),
.A2(n_515),
.B1(n_504),
.B2(n_493),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_473),
.B(n_380),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_515),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_561),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_479),
.A2(n_486),
.B(n_578),
.C(n_572),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_503),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_546),
.B(n_428),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_524),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_458),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_453),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_565),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_472),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_583),
.B(n_409),
.Y(n_654)
);

INVxp33_ASAP7_75t_L g655 ( 
.A(n_532),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_531),
.Y(n_656)
);

NOR3xp33_ASAP7_75t_L g657 ( 
.A(n_482),
.B(n_187),
.C(n_178),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g658 ( 
.A(n_494),
.B(n_194),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_469),
.B(n_391),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_485),
.B(n_179),
.C(n_185),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_472),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_471),
.B(n_405),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_587),
.B(n_204),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_471),
.B(n_405),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_476),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_503),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_476),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_512),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_L g669 ( 
.A1(n_447),
.A2(n_206),
.B1(n_218),
.B2(n_221),
.C(n_233),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_512),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_554),
.B(n_255),
.Y(n_671)
);

NOR2x1_ASAP7_75t_L g672 ( 
.A(n_523),
.B(n_229),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_471),
.B(n_194),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_477),
.B(n_405),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_477),
.B(n_197),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_579),
.B(n_581),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_489),
.B(n_208),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_535),
.B(n_262),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_489),
.B(n_222),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_565),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_524),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_460),
.B(n_267),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_449),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_449),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_513),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_455),
.B(n_481),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_503),
.B(n_222),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_555),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_455),
.B(n_231),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_576),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_481),
.B(n_231),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_481),
.B(n_232),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_516),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_492),
.B(n_232),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_492),
.B(n_235),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_470),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_464),
.B(n_235),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_492),
.B(n_246),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_518),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_495),
.B(n_249),
.Y(n_702)
);

BUFx6f_ASAP7_75t_SL g703 ( 
.A(n_585),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_518),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_572),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_495),
.B(n_249),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_520),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_495),
.B(n_254),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_563),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_520),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_510),
.B(n_254),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_522),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_510),
.B(n_256),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_566),
.B(n_582),
.C(n_500),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_522),
.Y(n_715)
);

AOI22x1_ASAP7_75t_L g716 ( 
.A1(n_585),
.A2(n_293),
.B1(n_264),
.B2(n_266),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_464),
.A2(n_293),
.B1(n_264),
.B2(n_266),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_510),
.B(n_256),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_585),
.B(n_268),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_498),
.A2(n_261),
.B1(n_288),
.B2(n_290),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_305),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_508),
.B(n_268),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_576),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_461),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_461),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_511),
.B(n_271),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_580),
.B(n_305),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_528),
.B(n_538),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_578),
.B(n_271),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_478),
.B(n_281),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_543),
.B(n_274),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_464),
.B(n_400),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_588),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_444),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_464),
.B(n_400),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_464),
.B(n_400),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_551),
.B(n_400),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_584),
.B(n_461),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_444),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_584),
.B(n_414),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_459),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_521),
.B(n_412),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_459),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_514),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_584),
.B(n_278),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_584),
.B(n_414),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_537),
.B(n_280),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_497),
.B(n_261),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_584),
.B(n_414),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_453),
.B(n_412),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_584),
.B(n_414),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_527),
.B(n_408),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_509),
.Y(n_753)
);

BUFx8_ASAP7_75t_L g754 ( 
.A(n_703),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_628),
.B(n_448),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_605),
.B(n_521),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_539),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_650),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_650),
.B(n_542),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_650),
.A2(n_562),
.B(n_569),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_654),
.B(n_540),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_591),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_616),
.B(n_454),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_643),
.B(n_540),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_592),
.B(n_507),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_646),
.B(n_540),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_646),
.B(n_540),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_591),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_608),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_656),
.B(n_615),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_600),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_637),
.A2(n_562),
.B(n_569),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_590),
.B(n_454),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_621),
.A2(n_586),
.B1(n_540),
.B2(n_544),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_631),
.A2(n_564),
.B1(n_571),
.B2(n_558),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_590),
.B(n_498),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_596),
.B(n_562),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_637),
.A2(n_569),
.B(n_541),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_637),
.A2(n_541),
.B(n_467),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_623),
.Y(n_780)
);

AO21x1_ASAP7_75t_L g781 ( 
.A1(n_658),
.A2(n_452),
.B(n_568),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_600),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_748),
.A2(n_527),
.B(n_544),
.C(n_559),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_651),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_603),
.B(n_452),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_687),
.A2(n_541),
.B(n_491),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_738),
.A2(n_541),
.B(n_491),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_604),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_SL g789 ( 
.A1(n_610),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_594),
.B(n_540),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_604),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_640),
.A2(n_573),
.B(n_568),
.C(n_462),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_649),
.B(n_527),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_634),
.A2(n_467),
.B(n_491),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_681),
.B(n_544),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_742),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_705),
.B(n_559),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_607),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_593),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_627),
.A2(n_559),
.B(n_560),
.C(n_488),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_607),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_634),
.A2(n_467),
.B(n_548),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_747),
.B(n_669),
.C(n_682),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_676),
.B(n_560),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_750),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_592),
.B(n_410),
.Y(n_807)
);

O2A1O1Ixp5_ASAP7_75t_L g808 ( 
.A1(n_627),
.A2(n_560),
.B(n_534),
.C(n_526),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_753),
.B(n_411),
.C(n_412),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_728),
.A2(n_589),
.B(n_659),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_728),
.A2(n_491),
.B(n_548),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_625),
.A2(n_689),
.B1(n_729),
.B2(n_630),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_626),
.B(n_573),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_648),
.B(n_567),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_629),
.B(n_488),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_611),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_613),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_608),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_653),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_661),
.B(n_484),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_662),
.A2(n_567),
.B(n_563),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_660),
.B(n_408),
.Y(n_823)
);

NOR2x1p5_ASAP7_75t_SL g824 ( 
.A(n_684),
.B(n_685),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_666),
.B(n_563),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_666),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_730),
.B(n_408),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_665),
.B(n_484),
.Y(n_828)
);

AND2x6_ASAP7_75t_SL g829 ( 
.A(n_678),
.B(n_7),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_671),
.B(n_408),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_667),
.B(n_499),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_668),
.B(n_499),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_663),
.B(n_563),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_723),
.B(n_733),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_608),
.B(n_563),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_664),
.A2(n_547),
.B(n_534),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_720),
.B(n_547),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_612),
.A2(n_526),
.B(n_501),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_670),
.B(n_501),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_683),
.B(n_686),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_613),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_L g842 ( 
.A(n_714),
.B(n_462),
.C(n_402),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_694),
.B(n_402),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_725),
.B(n_402),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_612),
.A2(n_402),
.B(n_397),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_696),
.B(n_397),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_614),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_397),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_707),
.B(n_397),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_640),
.A2(n_393),
.B(n_386),
.C(n_17),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_614),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_731),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_386),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_704),
.B(n_386),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_630),
.A2(n_393),
.B1(n_386),
.B2(n_17),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_620),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_642),
.A2(n_393),
.B(n_78),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_658),
.A2(n_393),
.B(n_13),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_710),
.B(n_85),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_722),
.A2(n_10),
.B(n_23),
.C(n_28),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_674),
.A2(n_93),
.B(n_153),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_709),
.A2(n_88),
.B(n_152),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_710),
.B(n_30),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_725),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_688),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_712),
.B(n_31),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_709),
.A2(n_61),
.B(n_148),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_647),
.B(n_31),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_620),
.Y(n_870)
);

INVx11_ASAP7_75t_L g871 ( 
.A(n_655),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_632),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_636),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_709),
.A2(n_98),
.B(n_146),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_647),
.B(n_595),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_636),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_641),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_666),
.B(n_57),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_709),
.A2(n_154),
.B(n_136),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_598),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_709),
.A2(n_132),
.B(n_130),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_606),
.A2(n_127),
.B1(n_125),
.B2(n_122),
.Y(n_882)
);

BUFx4f_ASAP7_75t_L g883 ( 
.A(n_688),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_712),
.B(n_34),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_675),
.A2(n_117),
.B(n_116),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_715),
.B(n_34),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_673),
.A2(n_106),
.B(n_105),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_601),
.B(n_39),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_601),
.B(n_597),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_677),
.A2(n_99),
.B(n_45),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_624),
.B(n_606),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_722),
.A2(n_44),
.B(n_46),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_599),
.B(n_46),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_724),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_724),
.A2(n_48),
.B(n_49),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_715),
.B(n_51),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_724),
.A2(n_51),
.B(n_52),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_645),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_673),
.A2(n_52),
.B(n_54),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_598),
.B(n_55),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_679),
.A2(n_740),
.B(n_751),
.Y(n_902)
);

BUFx10_ASAP7_75t_L g903 ( 
.A(n_703),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_652),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_602),
.B(n_617),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_657),
.B(n_688),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_622),
.B(n_719),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_619),
.B(n_680),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_719),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_652),
.B(n_680),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_690),
.A2(n_706),
.B(n_713),
.C(n_711),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_684),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_719),
.B(n_702),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_679),
.A2(n_749),
.B(n_746),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_726),
.A2(n_737),
.B(n_695),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_692),
.B(n_718),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_693),
.B(n_697),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_745),
.B(n_699),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_726),
.A2(n_700),
.B(n_708),
.C(n_639),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_732),
.A2(n_736),
.B(n_735),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_618),
.A2(n_633),
.B1(n_727),
.B2(n_717),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_700),
.A2(n_708),
.B1(n_609),
.B2(n_716),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_737),
.A2(n_752),
.B(n_699),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_618),
.A2(n_633),
.B1(n_672),
.B2(n_698),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_734),
.B(n_739),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_734),
.B(n_739),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_741),
.A2(n_743),
.B(n_745),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_743),
.B(n_638),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_655),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_691),
.B(n_635),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_691),
.B(n_650),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_804),
.A2(n_889),
.B(n_919),
.C(n_852),
.Y(n_932)
);

BUFx8_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_766),
.A2(n_767),
.B(n_920),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_758),
.A2(n_917),
.B(n_916),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_755),
.A2(n_775),
.B1(n_857),
.B2(n_758),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_903),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_866),
.B(n_875),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_835),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_758),
.A2(n_911),
.B(n_759),
.Y(n_940)
);

AO32x1_ASAP7_75t_L g941 ( 
.A1(n_855),
.A2(n_887),
.A3(n_924),
.B1(n_799),
.B2(n_813),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_758),
.B(n_875),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_801),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_SL g944 ( 
.A(n_918),
.B(n_906),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_833),
.A2(n_913),
.B(n_778),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_766),
.A2(n_767),
.B(n_813),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_895),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_883),
.B(n_909),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_835),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_760),
.A2(n_811),
.B(n_772),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_796),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_756),
.B(n_763),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_871),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_895),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_773),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_902),
.A2(n_914),
.B(n_921),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_921),
.A2(n_924),
.B(n_890),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_780),
.B(n_806),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_930),
.B(n_770),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_776),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_SL g961 ( 
.A1(n_777),
.A2(n_857),
.B(n_815),
.C(n_894),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_887),
.A2(n_893),
.B(n_892),
.C(n_757),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_SL g963 ( 
.A1(n_809),
.A2(n_915),
.B(n_774),
.C(n_842),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_762),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_768),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_893),
.A2(n_755),
.B(n_861),
.C(n_775),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_907),
.A2(n_883),
.B(n_909),
.C(n_905),
.Y(n_967)
);

BUFx12f_ASAP7_75t_L g968 ( 
.A(n_903),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_SL g969 ( 
.A(n_901),
.B(n_882),
.C(n_785),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_765),
.B(n_820),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_840),
.A2(n_922),
.B1(n_908),
.B2(n_855),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_764),
.A2(n_827),
.B(n_910),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_779),
.A2(n_927),
.B(n_923),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_864),
.A2(n_886),
.B(n_884),
.C(n_867),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_771),
.B(n_788),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_915),
.A2(n_885),
.B(n_838),
.C(n_845),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_765),
.B(n_837),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_895),
.B(n_865),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_761),
.A2(n_885),
.B(n_823),
.C(n_790),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_897),
.A2(n_931),
.B(n_900),
.C(n_799),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_824),
.A2(n_860),
.B(n_830),
.C(n_800),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_860),
.A2(n_873),
.B(n_841),
.C(n_904),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_754),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_787),
.A2(n_786),
.B(n_822),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_791),
.B(n_810),
.Y(n_985)
);

INVx6_ASAP7_75t_L g986 ( 
.A(n_754),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_789),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_929),
.B(n_807),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_817),
.B(n_847),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_801),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_858),
.Y(n_991)
);

AOI33xp33_ASAP7_75t_L g992 ( 
.A1(n_850),
.A2(n_851),
.A3(n_856),
.B1(n_872),
.B2(n_876),
.B3(n_877),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_865),
.B(n_769),
.Y(n_993)
);

OAI22x1_ASAP7_75t_L g994 ( 
.A1(n_829),
.A2(n_805),
.B1(n_878),
.B2(n_797),
.Y(n_994)
);

BUFx4f_ASAP7_75t_SL g995 ( 
.A(n_880),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_782),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_926),
.A2(n_825),
.B(n_812),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_798),
.B(n_818),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_783),
.A2(n_808),
.B(n_836),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_828),
.B(n_839),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_802),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_869),
.B(n_834),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_870),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_896),
.A2(n_898),
.B(n_793),
.C(n_928),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_826),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_SL g1006 ( 
.A(n_891),
.B(n_862),
.C(n_795),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_819),
.A2(n_781),
.B1(n_826),
.B2(n_899),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_912),
.A2(n_792),
.B(n_814),
.C(n_816),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_831),
.A2(n_832),
.B(n_803),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_834),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_853),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_844),
.B(n_859),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_869),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_SL g1014 ( 
.A1(n_845),
.A2(n_838),
.B(n_846),
.C(n_843),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_853),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_794),
.A2(n_854),
.B(n_848),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_854),
.B(n_925),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_844),
.B(n_879),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_888),
.A2(n_849),
.B(n_863),
.C(n_868),
.Y(n_1019)
);

XNOR2xp5_ASAP7_75t_L g1020 ( 
.A(n_874),
.B(n_881),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_925),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_925),
.B(n_628),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_925),
.B(n_605),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_925),
.A2(n_728),
.B(n_759),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_804),
.A2(n_755),
.B1(n_451),
.B2(n_646),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_L g1028 ( 
.A(n_758),
.B(n_804),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_784),
.B(n_521),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_762),
.Y(n_1030)
);

BUFx10_ASAP7_75t_L g1031 ( 
.A(n_763),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_784),
.B(n_521),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_754),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_SL g1034 ( 
.A1(n_890),
.A2(n_650),
.B(n_857),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_782),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_796),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_766),
.A2(n_767),
.B(n_920),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_754),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_SL g1041 ( 
.A1(n_833),
.A2(n_621),
.B(n_463),
.C(n_473),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_762),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_895),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_782),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_804),
.A2(n_852),
.B1(n_621),
.B2(n_714),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_762),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_762),
.Y(n_1048)
);

OA21x2_ASAP7_75t_L g1049 ( 
.A1(n_857),
.A2(n_838),
.B(n_845),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_755),
.B(n_628),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_L g1051 ( 
.A(n_758),
.B(n_804),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_796),
.B(n_517),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_782),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_895),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_755),
.B(n_628),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_782),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_755),
.B(n_628),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_796),
.B(n_517),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_804),
.A2(n_616),
.B(n_605),
.C(n_656),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_895),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_755),
.B(n_628),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_756),
.B(n_605),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_SL g1063 ( 
.A(n_758),
.B(n_618),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_852),
.B(n_804),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_804),
.A2(n_852),
.B1(n_621),
.B2(n_714),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_852),
.B(n_804),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_758),
.A2(n_650),
.B(n_637),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_756),
.B(n_605),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_SL g1069 ( 
.A(n_986),
.B(n_937),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_954),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_962),
.A2(n_932),
.B(n_1065),
.C(n_1046),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1067),
.A2(n_945),
.B(n_940),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_954),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_958),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_954),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_952),
.B(n_1062),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_965),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1067),
.A2(n_935),
.B(n_1026),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_1043),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1027),
.A2(n_1045),
.B(n_1040),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_969),
.A2(n_987),
.B1(n_970),
.B2(n_1066),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1016),
.A2(n_997),
.B(n_999),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_957),
.A2(n_936),
.A3(n_956),
.B(n_981),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_979),
.A2(n_936),
.B(n_1025),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1030),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_986),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_961),
.A2(n_1041),
.B(n_976),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_1043),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1024),
.A2(n_1009),
.B(n_1019),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1039),
.A2(n_972),
.B(n_1034),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1064),
.A2(n_977),
.B1(n_960),
.B2(n_1068),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_959),
.A2(n_1061),
.B1(n_1057),
.B2(n_1055),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1025),
.A2(n_1014),
.B(n_946),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1000),
.A2(n_1017),
.B(n_1004),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1042),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_1043),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_1050),
.A2(n_1057),
.B(n_1061),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_1054),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_966),
.A2(n_1059),
.B(n_980),
.C(n_974),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_955),
.B(n_1052),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_982),
.A2(n_971),
.A3(n_1008),
.B(n_1017),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1058),
.B(n_1011),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_1012),
.A2(n_1063),
.B(n_971),
.C(n_944),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1047),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1022),
.A2(n_941),
.A3(n_967),
.B(n_994),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1022),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1023),
.A2(n_946),
.B(n_963),
.C(n_934),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_934),
.A2(n_1037),
.B(n_1049),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1015),
.B(n_988),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1037),
.A2(n_1049),
.B(n_1018),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_975),
.A2(n_985),
.B(n_989),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_986),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1020),
.A2(n_942),
.B(n_993),
.Y(n_1115)
);

AO21x1_ASAP7_75t_L g1116 ( 
.A1(n_1007),
.A2(n_975),
.B(n_989),
.Y(n_1116)
);

BUFx2_ASAP7_75t_R g1117 ( 
.A(n_953),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1006),
.A2(n_998),
.B(n_985),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_951),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_948),
.A2(n_941),
.B(n_978),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_941),
.A2(n_1021),
.B(n_1060),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1048),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1054),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_992),
.A2(n_939),
.B(n_949),
.C(n_1003),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1001),
.A2(n_1053),
.B(n_996),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_947),
.A2(n_939),
.B(n_949),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1035),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1044),
.A2(n_1056),
.A3(n_1005),
.B(n_943),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_943),
.A2(n_1005),
.B(n_990),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1002),
.A2(n_938),
.B1(n_1013),
.B2(n_1036),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1054),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1010),
.A2(n_938),
.B(n_990),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1013),
.A2(n_1031),
.B(n_991),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1031),
.A2(n_1038),
.B(n_1033),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_933),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_933),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_995),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1029),
.A2(n_1032),
.B(n_968),
.C(n_983),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_954),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1140)
);

AO21x2_ASAP7_75t_L g1141 ( 
.A1(n_957),
.A2(n_956),
.B(n_940),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_954),
.Y(n_1142)
);

BUFx8_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_964),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_948),
.B(n_801),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_962),
.A2(n_804),
.B(n_932),
.C(n_1046),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_962),
.A2(n_804),
.B(n_932),
.C(n_1046),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_951),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_952),
.B(n_605),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_964),
.Y(n_1152)
);

AO21x1_ASAP7_75t_L g1153 ( 
.A1(n_962),
.A2(n_957),
.B(n_1025),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_964),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1155)
);

AOI22x1_ASAP7_75t_L g1156 ( 
.A1(n_957),
.A2(n_994),
.B1(n_935),
.B2(n_656),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1157)
);

BUFx10_ASAP7_75t_L g1158 ( 
.A(n_986),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1067),
.A2(n_758),
.B(n_650),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1029),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_964),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_957),
.A2(n_979),
.B(n_936),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_954),
.Y(n_1163)
);

AOI221x1_ASAP7_75t_L g1164 ( 
.A1(n_957),
.A2(n_932),
.B1(n_936),
.B2(n_857),
.C(n_956),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_964),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_932),
.A2(n_804),
.B1(n_1049),
.B2(n_1057),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_957),
.A2(n_932),
.B1(n_936),
.B2(n_857),
.C(n_956),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_932),
.A2(n_804),
.B1(n_1049),
.B2(n_1057),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_SL g1172 ( 
.A1(n_962),
.A2(n_966),
.B1(n_631),
.B2(n_932),
.C(n_775),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1173)
);

BUFx2_ASAP7_75t_SL g1174 ( 
.A(n_991),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_932),
.A2(n_605),
.B(n_616),
.C(n_656),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_964),
.Y(n_1176)
);

BUFx2_ASAP7_75t_R g1177 ( 
.A(n_953),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_957),
.A2(n_979),
.B(n_936),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_954),
.Y(n_1179)
);

AOI211x1_ASAP7_75t_L g1180 ( 
.A1(n_1064),
.A2(n_804),
.B(n_893),
.C(n_1066),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1067),
.A2(n_758),
.B(n_650),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_933),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_957),
.A2(n_979),
.B(n_936),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1067),
.A2(n_758),
.B(n_650),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_932),
.A2(n_804),
.B1(n_1049),
.B2(n_1057),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1067),
.A2(n_758),
.B(n_650),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_964),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_962),
.A2(n_804),
.B(n_932),
.C(n_1046),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_970),
.A2(n_804),
.B1(n_952),
.B2(n_969),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_952),
.B(n_605),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_951),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_964),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_933),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_962),
.A2(n_804),
.B(n_932),
.C(n_1046),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_954),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_957),
.A2(n_936),
.A3(n_956),
.B(n_981),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_952),
.A2(n_421),
.B1(n_804),
.B2(n_586),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_950),
.A2(n_973),
.B(n_984),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_938),
.B(n_977),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1077),
.A2(n_1153),
.B1(n_1191),
.B2(n_1086),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1191),
.A2(n_1086),
.B1(n_1083),
.B2(n_1204),
.Y(n_1208)
);

AOI22x1_ASAP7_75t_SL g1209 ( 
.A1(n_1160),
.A2(n_1074),
.B1(n_1197),
.B2(n_1119),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1162),
.A2(n_1178),
.B1(n_1183),
.B2(n_1185),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1151),
.A2(n_1196),
.B1(n_1172),
.B2(n_1093),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1143),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1144),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1094),
.B(n_1075),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1094),
.A2(n_1165),
.B1(n_1189),
.B2(n_1173),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1162),
.A2(n_1178),
.B1(n_1183),
.B2(n_1170),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1119),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1117),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_1192),
.B1(n_1169),
.B2(n_1149),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1113),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1177),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1081),
.Y(n_1222)
);

INVx6_ASAP7_75t_L g1223 ( 
.A(n_1088),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1088),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1167),
.A2(n_1170),
.B1(n_1185),
.B2(n_1099),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1167),
.A2(n_1099),
.B1(n_1156),
.B2(n_1095),
.Y(n_1226)
);

BUFx4f_ASAP7_75t_SL g1227 ( 
.A(n_1136),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1114),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1155),
.B(n_1171),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1148),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1115),
.A2(n_1195),
.B1(n_1095),
.B2(n_1135),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1074),
.B2(n_1206),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1142),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1143),
.Y(n_1234)
);

INVx6_ASAP7_75t_L g1235 ( 
.A(n_1114),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1111),
.A2(n_1116),
.B1(n_1110),
.B2(n_1089),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1142),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1089),
.A2(n_1118),
.B1(n_1104),
.B2(n_1166),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1158),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1142),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1137),
.Y(n_1242)
);

BUFx2_ASAP7_75t_SL g1243 ( 
.A(n_1163),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1079),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1071),
.A2(n_1147),
.B1(n_1146),
.B2(n_1190),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1200),
.A2(n_1102),
.B1(n_1175),
.B2(n_1180),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1118),
.A2(n_1176),
.B1(n_1161),
.B2(n_1154),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1172),
.A2(n_1206),
.B1(n_1130),
.B2(n_1069),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1163),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1174),
.A2(n_1132),
.B1(n_1112),
.B2(n_1141),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1073),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1097),
.A2(n_1122),
.B1(n_1187),
.B2(n_1152),
.Y(n_1252)
);

NAND2x1_ASAP7_75t_L g1253 ( 
.A(n_1106),
.B(n_1198),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1163),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1073),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1130),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1127),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1125),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1141),
.A2(n_1108),
.B1(n_1132),
.B2(n_1120),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_SL g1260 ( 
.A(n_1073),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1134),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1131),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1128),
.Y(n_1263)
);

CKINVDCx6p67_ASAP7_75t_R g1264 ( 
.A(n_1076),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1070),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1070),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1103),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1076),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1201),
.B(n_1107),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1121),
.A2(n_1092),
.B1(n_1145),
.B2(n_1164),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1145),
.A2(n_1168),
.B1(n_1096),
.B2(n_1133),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1076),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1081),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1126),
.A2(n_1072),
.B1(n_1201),
.B2(n_1139),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1124),
.Y(n_1276)
);

CKINVDCx14_ASAP7_75t_R g1277 ( 
.A(n_1098),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1107),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_SL g1279 ( 
.A(n_1098),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1098),
.A2(n_1179),
.B1(n_1139),
.B2(n_1123),
.Y(n_1280)
);

CKINVDCx6p67_ASAP7_75t_R g1281 ( 
.A(n_1123),
.Y(n_1281)
);

INVx6_ASAP7_75t_L g1282 ( 
.A(n_1090),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1139),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1179),
.A2(n_1100),
.B1(n_1090),
.B2(n_1084),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1179),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1105),
.A2(n_1100),
.B1(n_1129),
.B2(n_1205),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1078),
.A2(n_1188),
.B1(n_1157),
.B2(n_1194),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1150),
.A2(n_1193),
.B1(n_1202),
.B2(n_1091),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1138),
.Y(n_1289)
);

INVx6_ASAP7_75t_SL g1290 ( 
.A(n_1085),
.Y(n_1290)
);

INVx8_ASAP7_75t_L g1291 ( 
.A(n_1080),
.Y(n_1291)
);

INVx8_ASAP7_75t_L g1292 ( 
.A(n_1082),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1203),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1159),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1181),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1184),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1186),
.Y(n_1297)
);

BUFx4_ASAP7_75t_R g1298 ( 
.A(n_1088),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1143),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1074),
.B(n_1104),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1077),
.A2(n_901),
.B1(n_952),
.B2(n_1191),
.Y(n_1301)
);

INVx4_ASAP7_75t_L g1302 ( 
.A(n_1142),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1088),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1148),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1113),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1113),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1077),
.A2(n_509),
.B(n_403),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1088),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1148),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1077),
.A2(n_952),
.B1(n_1083),
.B2(n_804),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1077),
.A2(n_804),
.B1(n_631),
.B2(n_952),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1113),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1087),
.Y(n_1313)
);

CKINVDCx16_ASAP7_75t_R g1314 ( 
.A(n_1136),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1087),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1077),
.A2(n_421),
.B1(n_952),
.B2(n_621),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1077),
.B(n_977),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1143),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1077),
.A2(n_804),
.B1(n_383),
.B2(n_776),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1142),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1143),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1077),
.A2(n_804),
.B1(n_631),
.B2(n_952),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1148),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1291),
.B(n_1292),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1311),
.A2(n_1322),
.B1(n_1210),
.B2(n_1216),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1233),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1290),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1311),
.A2(n_1322),
.B1(n_1210),
.B2(n_1216),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1310),
.A2(n_1245),
.B1(n_1208),
.B2(n_1207),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1294),
.A2(n_1297),
.B(n_1220),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1267),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1278),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1263),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1294),
.A2(n_1297),
.B(n_1220),
.Y(n_1334)
);

AOI222xp33_ASAP7_75t_L g1335 ( 
.A1(n_1208),
.A2(n_1307),
.B1(n_1207),
.B2(n_1270),
.C1(n_1246),
.C2(n_1317),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1305),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1306),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1258),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1312),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1219),
.B(n_1215),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1293),
.Y(n_1341)
);

BUFx2_ASAP7_75t_SL g1342 ( 
.A(n_1261),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1312),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1269),
.B(n_1225),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1290),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1316),
.A2(n_1231),
.B(n_1226),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1290),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1300),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1319),
.B(n_1301),
.Y(n_1349)
);

AO21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1226),
.A2(n_1225),
.B(n_1238),
.Y(n_1350)
);

NAND2xp33_ASAP7_75t_R g1351 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1296),
.A2(n_1259),
.B(n_1271),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1291),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1256),
.B(n_1211),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1244),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1291),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1271),
.A2(n_1236),
.B(n_1259),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1257),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1295),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1253),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1213),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1295),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1219),
.B(n_1215),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1313),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1239),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1315),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1236),
.A2(n_1238),
.B(n_1272),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1237),
.B(n_1302),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1212),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1214),
.B(n_1247),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1276),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1217),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1272),
.A2(n_1275),
.B(n_1247),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1233),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1230),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1229),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1309),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1248),
.A2(n_1288),
.B(n_1287),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1252),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1254),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1252),
.A2(n_1323),
.B1(n_1304),
.B2(n_1289),
.C(n_1250),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1265),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1262),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1286),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1243),
.B(n_1254),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1275),
.B(n_1284),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1249),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1280),
.B(n_1266),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1320),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1222),
.A2(n_1274),
.B(n_1298),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1232),
.B(n_1224),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1348),
.B(n_1277),
.Y(n_1392)
);

AO32x1_ASAP7_75t_L g1393 ( 
.A1(n_1325),
.A2(n_1285),
.A3(n_1273),
.B1(n_1268),
.B2(n_1209),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1325),
.A2(n_1241),
.B(n_1277),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1344),
.B(n_1283),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1328),
.A2(n_1222),
.B(n_1274),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1383),
.B(n_1377),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1328),
.B(n_1298),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1352),
.A2(n_1254),
.B(n_1264),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1346),
.A2(n_1241),
.B(n_1240),
.C(n_1283),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1383),
.B(n_1255),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1329),
.A2(n_1223),
.B1(n_1308),
.B2(n_1228),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1352),
.A2(n_1281),
.B(n_1279),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1344),
.B(n_1285),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1346),
.A2(n_1227),
.B(n_1299),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1356),
.B(n_1242),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1349),
.A2(n_1279),
.B(n_1260),
.C(n_1321),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1375),
.B(n_1314),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1351),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1335),
.A2(n_1318),
.B1(n_1234),
.B2(n_1227),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1354),
.A2(n_1235),
.B1(n_1303),
.B2(n_1260),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_SL g1412 ( 
.A1(n_1381),
.A2(n_1235),
.B(n_1303),
.C(n_1282),
.Y(n_1412)
);

NAND2xp33_ASAP7_75t_L g1413 ( 
.A(n_1340),
.B(n_1282),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1342),
.B(n_1382),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1381),
.A2(n_1251),
.B(n_1282),
.C(n_1340),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1342),
.B(n_1376),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1355),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1335),
.A2(n_1363),
.B1(n_1350),
.B2(n_1370),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1372),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1391),
.A2(n_1363),
.B1(n_1370),
.B2(n_1384),
.Y(n_1420)
);

NAND4xp25_ASAP7_75t_L g1421 ( 
.A(n_1388),
.B(n_1391),
.C(n_1379),
.D(n_1361),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1352),
.A2(n_1330),
.B(n_1334),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1384),
.A2(n_1372),
.B1(n_1388),
.B2(n_1379),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1327),
.B(n_1345),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1341),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1347),
.B(n_1390),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1373),
.A2(n_1386),
.B(n_1359),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1347),
.B(n_1390),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1358),
.B(n_1357),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1324),
.A2(n_1357),
.B(n_1353),
.Y(n_1430)
);

AO32x2_ASAP7_75t_L g1431 ( 
.A1(n_1380),
.A2(n_1326),
.A3(n_1341),
.B1(n_1332),
.B2(n_1331),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1357),
.B(n_1338),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1357),
.B(n_1338),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1324),
.A2(n_1357),
.B(n_1385),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1359),
.A2(n_1362),
.B(n_1380),
.C(n_1389),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1432),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1429),
.B(n_1332),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1426),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1429),
.B(n_1367),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1432),
.B(n_1333),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1434),
.B(n_1367),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1434),
.B(n_1367),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1431),
.B(n_1367),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1421),
.B(n_1387),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1410),
.A2(n_1367),
.B1(n_1378),
.B2(n_1371),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1425),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1431),
.B(n_1336),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1431),
.B(n_1336),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1426),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1428),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1409),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1417),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_L g1454 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1420),
.B(n_1387),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1431),
.B(n_1427),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1336),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1428),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1400),
.B(n_1360),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1428),
.B(n_1435),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1444),
.A2(n_1430),
.B(n_1457),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1451),
.B(n_1424),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1438),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1438),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1442),
.B(n_1399),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1447),
.B(n_1419),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1458),
.B(n_1397),
.Y(n_1467)
);

NAND2x1_ASAP7_75t_L g1468 ( 
.A(n_1454),
.B(n_1403),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

NOR2x1_ASAP7_75t_SL g1470 ( 
.A(n_1459),
.B(n_1324),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1458),
.B(n_1414),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1451),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1438),
.Y(n_1473)
);

AOI211xp5_ASAP7_75t_L g1474 ( 
.A1(n_1459),
.A2(n_1412),
.B(n_1398),
.C(n_1415),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1458),
.A2(n_1339),
.A3(n_1337),
.B(n_1343),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1439),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1448),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1454),
.A2(n_1418),
.B1(n_1398),
.B2(n_1394),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1446),
.A2(n_1418),
.B1(n_1423),
.B2(n_1412),
.C(n_1415),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1452),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1454),
.A2(n_1413),
.B(n_1407),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1446),
.A2(n_1407),
.B1(n_1409),
.B2(n_1396),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1448),
.Y(n_1484)
);

AOI33xp33_ASAP7_75t_L g1485 ( 
.A1(n_1456),
.A2(n_1395),
.A3(n_1404),
.B1(n_1392),
.B2(n_1401),
.B3(n_1416),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1439),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1449),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1441),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1449),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1437),
.B(n_1433),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1452),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1395),
.Y(n_1492)
);

INVx4_ASAP7_75t_L g1493 ( 
.A(n_1453),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1455),
.C(n_1456),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1441),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1493),
.Y(n_1496)
);

NAND2x1_ASAP7_75t_L g1497 ( 
.A(n_1493),
.B(n_1486),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1494),
.B(n_1463),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_SL g1499 ( 
.A(n_1474),
.B(n_1456),
.C(n_1408),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1473),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1463),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1476),
.B(n_1450),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1464),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1494),
.B(n_1437),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1493),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1468),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1482),
.B(n_1456),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1479),
.A2(n_1405),
.B1(n_1445),
.B2(n_1413),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1450),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1477),
.B(n_1484),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1495),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1495),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1493),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1441),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1490),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1490),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1462),
.B(n_1450),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1462),
.B(n_1460),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1462),
.B(n_1460),
.Y(n_1523)
);

INVx3_ASAP7_75t_SL g1524 ( 
.A(n_1491),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1462),
.B(n_1460),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1521),
.B(n_1470),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1512),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1498),
.B(n_1466),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1497),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1498),
.B(n_1477),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1524),
.B(n_1480),
.Y(n_1534)
);

NOR2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1468),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1521),
.B(n_1470),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1522),
.B(n_1465),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1522),
.B(n_1465),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1504),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1504),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1513),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1499),
.A2(n_1479),
.B1(n_1483),
.B2(n_1478),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1510),
.A2(n_1481),
.B(n_1483),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1519),
.B(n_1520),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1500),
.Y(n_1551)
);

NAND2xp67_ASAP7_75t_L g1552 ( 
.A(n_1524),
.B(n_1365),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1526),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1465),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1516),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1516),
.Y(n_1559)
);

AOI211xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1519),
.A2(n_1474),
.B(n_1411),
.C(n_1402),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1500),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1525),
.B(n_1487),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1487),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1503),
.B(n_1489),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1461),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1508),
.Y(n_1567)
);

INVxp33_ASAP7_75t_L g1568 ( 
.A(n_1503),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1520),
.B(n_1489),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1549),
.B(n_1485),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1535),
.B(n_1524),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1567),
.Y(n_1572)
);

AND4x1_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1481),
.C(n_1510),
.D(n_1368),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1528),
.B(n_1508),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1553),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1547),
.Y(n_1576)
);

NAND2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1551),
.Y(n_1578)
);

AOI32xp33_ASAP7_75t_L g1579 ( 
.A1(n_1560),
.A2(n_1455),
.A3(n_1444),
.B1(n_1440),
.B2(n_1443),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1551),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1552),
.B(n_1369),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1553),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1534),
.B(n_1486),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1541),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1542),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1528),
.B(n_1536),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1530),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1549),
.B(n_1518),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1530),
.B(n_1509),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1552),
.B(n_1406),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1544),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1511),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1543),
.B(n_1509),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1547),
.B(n_1471),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1467),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1537),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.B(n_1514),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1550),
.B(n_1467),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1550),
.B(n_1501),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1544),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1537),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1573),
.A2(n_1532),
.B(n_1543),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1571),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1599),
.Y(n_1607)
);

AOI32xp33_ASAP7_75t_L g1608 ( 
.A1(n_1570),
.A2(n_1532),
.A3(n_1565),
.B1(n_1555),
.B2(n_1564),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1584),
.Y(n_1609)
);

XNOR2x2_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1566),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1576),
.A2(n_1460),
.B1(n_1556),
.B2(n_1514),
.Y(n_1611)
);

OAI21xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1579),
.A2(n_1531),
.B(n_1566),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1529),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1588),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1584),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1573),
.B(n_1406),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1529),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1578),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1587),
.B(n_1538),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1529),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1579),
.A2(n_1556),
.B(n_1531),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1594),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

AOI222xp33_ASAP7_75t_L g1626 ( 
.A1(n_1577),
.A2(n_1569),
.B1(n_1545),
.B2(n_1539),
.C1(n_1540),
.C2(n_1533),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1596),
.A2(n_1569),
.B(n_1562),
.Y(n_1627)
);

AOI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1596),
.A2(n_1545),
.B1(n_1539),
.B2(n_1533),
.C1(n_1540),
.C2(n_1564),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1586),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1610),
.A2(n_1578),
.B(n_1580),
.C(n_1581),
.Y(n_1630)
);

NAND4xp25_ASAP7_75t_L g1631 ( 
.A(n_1614),
.B(n_1583),
.C(n_1592),
.D(n_1580),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1619),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1605),
.B(n_1593),
.C(n_1591),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1624),
.B(n_1574),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1606),
.A2(n_1574),
.B(n_1598),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1610),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1608),
.B(n_1599),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1619),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_1600),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1617),
.A2(n_1604),
.B1(n_1603),
.B2(n_1593),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1628),
.B(n_1604),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1609),
.Y(n_1644)
);

NAND2x1p5_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1531),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1627),
.B(n_1600),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1612),
.A2(n_1602),
.B(n_1595),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1613),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1637),
.A2(n_1623),
.B1(n_1626),
.B2(n_1625),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1632),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_L g1651 ( 
.A1(n_1637),
.A2(n_1611),
.B(n_1620),
.Y(n_1651)
);

OAI321xp33_ASAP7_75t_L g1652 ( 
.A1(n_1631),
.A2(n_1629),
.A3(n_1622),
.B1(n_1616),
.B2(n_1615),
.C(n_1595),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1635),
.B(n_1607),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1640),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1641),
.A2(n_1607),
.B1(n_1545),
.B2(n_1539),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1633),
.Y(n_1656)
);

XOR2x2_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1406),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

XOR2x2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.B(n_1590),
.Y(n_1659)
);

AOI321xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1630),
.A2(n_1590),
.A3(n_1591),
.B1(n_1603),
.B2(n_1531),
.C(n_1562),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1649),
.A2(n_1630),
.B(n_1642),
.C(n_1643),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1652),
.A2(n_1642),
.B(n_1647),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1653),
.B(n_1636),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_SL g1664 ( 
.A(n_1649),
.B(n_1641),
.C(n_1648),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1656),
.B(n_1651),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1659),
.B(n_1646),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1655),
.B(n_1645),
.Y(n_1667)
);

NAND4xp75_ASAP7_75t_L g1668 ( 
.A(n_1660),
.B(n_1650),
.C(n_1654),
.D(n_1658),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1657),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1665),
.B(n_1639),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1661),
.A2(n_1645),
.B(n_1582),
.Y(n_1671)
);

AOI21xp33_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_1582),
.B(n_1575),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1662),
.A2(n_1582),
.B(n_1575),
.C(n_1563),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1664),
.A2(n_1575),
.B1(n_1557),
.B2(n_1548),
.C(n_1559),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1671),
.A2(n_1668),
.B(n_1663),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1670),
.B(n_1667),
.C(n_1669),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1672),
.A2(n_1553),
.B1(n_1561),
.B2(n_1527),
.C(n_1558),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1674),
.Y(n_1678)
);

NAND4xp25_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1563),
.C(n_1555),
.D(n_1368),
.Y(n_1679)
);

OAI321xp33_ASAP7_75t_L g1680 ( 
.A1(n_1671),
.A2(n_1559),
.A3(n_1558),
.B1(n_1557),
.B2(n_1546),
.C(n_1548),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1546),
.C(n_1561),
.Y(n_1681)
);

NOR2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1678),
.B(n_1679),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1680),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1675),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1677),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1684),
.A2(n_1561),
.B1(n_1507),
.B2(n_1517),
.Y(n_1686)
);

AND3x1_ASAP7_75t_L g1687 ( 
.A(n_1683),
.B(n_1496),
.C(n_1507),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1681),
.B(n_1501),
.Y(n_1688)
);

XNOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1687),
.B(n_1682),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1685),
.B(n_1688),
.C(n_1686),
.Y(n_1690)
);

XNOR2xp5_ASAP7_75t_L g1691 ( 
.A(n_1690),
.B(n_1538),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1691),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1692),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1517),
.B(n_1507),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1554),
.B(n_1506),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1694),
.A2(n_1554),
.B(n_1506),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1517),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1697),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1696),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_R g1700 ( 
.A1(n_1699),
.A2(n_1496),
.B1(n_1527),
.B2(n_1514),
.C(n_1393),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1698),
.B(n_1374),
.C(n_1526),
.Y(n_1701)
);


endmodule