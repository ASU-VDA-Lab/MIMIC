module real_jpeg_26536_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_257, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_257;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_16),
.B1(n_53),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_0),
.A2(n_16),
.B1(n_43),
.B2(n_44),
.Y(n_205)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_22),
.B(n_26),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_29),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_5),
.A2(n_6),
.B(n_54),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_5),
.B(n_130),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_8),
.B(n_25),
.C(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_9),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_186)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_10),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_68),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_30),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_30),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_19),
.B1(n_27),
.B2(n_29),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_15),
.A2(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_17),
.A2(n_23),
.B(n_34),
.C(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_45),
.Y(n_46)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_61),
.C(n_62),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_31),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.C(n_48),
.Y(n_31)
);

AOI211xp5_ASAP7_75t_L g77 ( 
.A1(n_32),
.A2(n_78),
.B(n_80),
.C(n_85),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_32),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_32),
.A2(n_86),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_32),
.A2(n_86),
.B1(n_200),
.B2(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_32),
.A2(n_86),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_32),
.A2(n_200),
.B(n_220),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_32),
.A2(n_86),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_32),
.A2(n_86),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_32),
.B(n_48),
.C(n_233),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_32),
.B(n_242),
.C(n_243),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_34),
.A2(n_44),
.B(n_56),
.C(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_34),
.B(n_52),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_34),
.B(n_139),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_34),
.A2(n_43),
.B(n_45),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_36),
.A2(n_48),
.B1(n_49),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_36),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_38),
.A2(n_83),
.B1(n_130),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_48),
.A2(n_49),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_52),
.A2(n_57),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_52),
.A2(n_57),
.B1(n_60),
.B2(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_53),
.B(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_61),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_249),
.B(n_254),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_227),
.A3(n_244),
.B1(n_247),
.B2(n_248),
.C(n_257),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_211),
.B(n_226),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_192),
.B(n_210),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_117),
.B(n_174),
.C(n_191),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_107),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_74),
.B(n_107),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_96),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_87),
.B2(n_88),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_76),
.B(n_88),
.C(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_84),
.B1(n_89),
.B2(n_95),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_84),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_78),
.A2(n_84),
.B1(n_124),
.B2(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_103),
.C(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_78),
.A2(n_84),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_78),
.B(n_157),
.C(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_78),
.B(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_78),
.A2(n_84),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_78),
.B(n_183),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_86),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_84),
.B(n_151),
.C(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_82),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_81),
.B(n_86),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_103),
.C(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_82),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_82),
.B(n_217),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_85),
.A2(n_106),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_85),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_90),
.A2(n_94),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_106),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_97),
.A2(n_98),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_97),
.A2(n_98),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_104),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_104),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_104),
.B1(n_115),
.B2(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_103),
.B(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_114),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_108),
.A2(n_109),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_111),
.B1(n_147),
.B2(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_173),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_166),
.B(n_172),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_153),
.B(n_165),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_144),
.B(n_152),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_132),
.B(n_143),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_176),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_187),
.C(n_189),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_207),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_199),
.C(n_207),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_197),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_208),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_206),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_224),
.B2(n_225),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.C(n_225),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_229),
.C(n_235),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_229),
.CI(n_235),
.CON(n_246),
.SN(n_246)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);


endmodule