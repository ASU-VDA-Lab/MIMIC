module real_jpeg_26120_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_249;
wire n_166;
wire n_292;
wire n_176;
wire n_221;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_0),
.B(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_0),
.B(n_31),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_0),
.B(n_45),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_0),
.B(n_36),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_0),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_0),
.B(n_43),
.Y(n_236)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_2),
.B(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_25),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_36),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_31),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_2),
.B(n_45),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_3),
.B(n_36),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_31),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_17),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_4),
.B(n_130),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_6),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_6),
.B(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_6),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_36),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_31),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_36),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_13),
.B(n_31),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_13),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_36),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_14),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_43),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_14),
.B(n_25),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_14),
.B(n_45),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_36),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_14),
.B(n_51),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_16),
.B(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_16),
.B(n_51),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_16),
.B(n_45),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_16),
.B(n_43),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_16),
.B(n_31),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_36),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_16),
.B(n_25),
.Y(n_244)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_17),
.Y(n_131)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_17),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_150),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_52),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_31),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_38),
.B1(n_59),
.B2(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_55),
.C(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_35),
.B(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_70),
.SN(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_47),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_71),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.C(n_70),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_54),
.B(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_65),
.C(n_66),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_67),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_70),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_86),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.C(n_84),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_74),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.C(n_80),
.Y(n_74)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_77),
.CI(n_80),
.CON(n_94),
.SN(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_84),
.B1(n_90),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_88),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_105),
.C(n_109),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_105),
.CI(n_109),
.CON(n_121),
.SN(n_121)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_101),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_94),
.B(n_290),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_94),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_95),
.B(n_101),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_98),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.C(n_118),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_138),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.CI(n_116),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_297)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_121),
.Y(n_298)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_125),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.C(n_139),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_126),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.C(n_133),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_127),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_128),
.A2(n_129),
.B(n_132),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_128),
.B(n_133),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.C(n_136),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_134),
.B(n_135),
.CI(n_136),
.CON(n_256),
.SN(n_256)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_137),
.B(n_139),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.C(n_148),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_140),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_145),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_141),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_144),
.B(n_145),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_295),
.C(n_296),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_285),
.C(n_286),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_270),
.C(n_271),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_249),
.C(n_250),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_224),
.C(n_225),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_186),
.C(n_198),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_165),
.C(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_160),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_178),
.C(n_179),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_185),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_197),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_191),
.B1(n_197),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_220),
.C(n_221),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.C(n_212),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_238),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_239),
.C(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_233),
.C(n_234),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_232),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_234),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.CI(n_237),
.CON(n_234),
.SN(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_248),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.C(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_258),
.C(n_261),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_256),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_280),
.B2(n_284),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_281),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_293),
.B2(n_294),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_295)
);


endmodule