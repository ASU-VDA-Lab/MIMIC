module fake_jpeg_259_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_41),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_46),
.B(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_41),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_43),
.C(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_62),
.B1(n_50),
.B2(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_47),
.B(n_59),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_82),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_3),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_74),
.A3(n_73),
.B1(n_68),
.B2(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_69),
.B1(n_19),
.B2(n_20),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_17),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_22),
.C(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_101),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_4),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_8),
.Y(n_112)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_91),
.B1(n_93),
.B2(n_97),
.C(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_112),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_21),
.B(n_32),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_107),
.B1(n_111),
.B2(n_93),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_34),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_24),
.C(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

OA21x2_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_119),
.B(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_109),
.B1(n_114),
.B2(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_123),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_107),
.A3(n_113),
.B1(n_103),
.B2(n_104),
.C1(n_12),
.C2(n_8),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_124),
.B(n_122),
.C(n_125),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_127),
.A3(n_124),
.B1(n_117),
.B2(n_116),
.C1(n_13),
.C2(n_9),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_10),
.B(n_14),
.Y(n_132)
);


endmodule