module fake_netlist_6_2791_n_5152 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5152);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5152;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_1781;
wire n_1971;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_858;
wire n_2049;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_2016;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_1077;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_740;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_930;
wire n_2620;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_3147;
wire n_2662;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_1003;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_3289;
wire n_2733;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_4203;
wire n_3641;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_2108;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2944;
wire n_2348;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_342),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_282),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_647),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_488),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_296),
.Y(n_713)
);

INVx4_ASAP7_75t_R g714 ( 
.A(n_149),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_246),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_349),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_240),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_677),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_3),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_641),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_173),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_534),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_373),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_472),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_410),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_703),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_481),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_166),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_646),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_125),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_515),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_338),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_570),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_234),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_298),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_205),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_383),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_456),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_582),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_511),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_393),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_618),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_375),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_627),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_591),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_50),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_10),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_328),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_190),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_439),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_18),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_665),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_542),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_412),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_360),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_215),
.Y(n_756)
);

BUFx10_ASAP7_75t_L g757 ( 
.A(n_471),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_293),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_177),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_476),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_266),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_335),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_481),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_290),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_358),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_219),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_286),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_290),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_323),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_528),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_158),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_505),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_365),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_578),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_298),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_83),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_39),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_44),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_690),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_201),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_590),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_585),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_607),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_686),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_701),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_278),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_691),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_6),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_707),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_365),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_562),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_338),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_283),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_153),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_670),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_223),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_487),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_247),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_21),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_658),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_663),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_378),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_100),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_16),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_226),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_477),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_473),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_0),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_300),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_81),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_693),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_155),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_144),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_650),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_239),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_252),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_5),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_42),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_410),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_593),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_530),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_693),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_395),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_74),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_74),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_119),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_23),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_387),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_191),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_360),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_102),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_226),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_495),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_575),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_424),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_679),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_292),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_614),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_115),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_533),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_665),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_66),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_195),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_671),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_675),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_393),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_506),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_83),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_603),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_146),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_279),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_657),
.Y(n_853)
);

BUFx10_ASAP7_75t_L g854 ( 
.A(n_206),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_674),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_318),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_204),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_112),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_488),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_452),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_241),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_364),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_651),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_633),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_422),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_640),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_41),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_249),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_118),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_688),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_413),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_575),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_397),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_592),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_476),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_362),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_291),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_223),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_336),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_621),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_85),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_686),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_539),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_570),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_189),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_482),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_101),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_705),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_672),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_31),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_673),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_520),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_33),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_327),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_629),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_241),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_609),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_152),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_527),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_66),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_635),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_120),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_21),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_457),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_284),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_140),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_227),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_191),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_339),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_183),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_230),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_115),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_300),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_115),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_525),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_489),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_145),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_295),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_361),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_200),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_699),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_539),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_469),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_516),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_64),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_444),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_235),
.Y(n_927)
);

BUFx10_ASAP7_75t_L g928 ( 
.A(n_29),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_184),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_653),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_592),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_204),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_368),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_316),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_364),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_438),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_65),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_623),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_470),
.Y(n_939)
);

CKINVDCx14_ASAP7_75t_R g940 ( 
.A(n_214),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_583),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_60),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_125),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_326),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_707),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_193),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_46),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_593),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_333),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_218),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_560),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_285),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_56),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_254),
.Y(n_954)
);

CKINVDCx14_ASAP7_75t_R g955 ( 
.A(n_634),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_545),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_13),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_694),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_400),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_461),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_239),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_104),
.Y(n_962)
);

INVxp33_ASAP7_75t_L g963 ( 
.A(n_316),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_141),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_94),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_617),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_431),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_387),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_635),
.Y(n_969)
);

BUFx10_ASAP7_75t_L g970 ( 
.A(n_630),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_506),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_110),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_345),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_374),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_159),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_579),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_457),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_231),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_688),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_42),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_522),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_440),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_123),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_280),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_318),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_313),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_479),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_248),
.Y(n_988)
);

BUFx5_ASAP7_75t_L g989 ( 
.A(n_248),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_4),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_39),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_267),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_329),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_228),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_230),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_351),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_601),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_125),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_557),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_425),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_121),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_278),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_355),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_234),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_443),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_618),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_145),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_209),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_144),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_669),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_333),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_16),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_495),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_297),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_15),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_114),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_391),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_180),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_390),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_462),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_647),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_659),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_202),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_395),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_429),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_613),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_196),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_232),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_331),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_256),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_553),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_373),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_482),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_41),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_23),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_475),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_513),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_155),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_470),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_199),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_416),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_100),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_349),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_676),
.Y(n_1044)
);

CKINVDCx14_ASAP7_75t_R g1045 ( 
.A(n_754),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_950),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_989),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_989),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_777),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_989),
.Y(n_1050)
);

BUFx5_ASAP7_75t_L g1051 ( 
.A(n_710),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_989),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_989),
.Y(n_1053)
);

XOR2xp5_ASAP7_75t_L g1054 ( 
.A(n_940),
.B(n_0),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_989),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_989),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_989),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_955),
.B(n_0),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_803),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_803),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_803),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_803),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_803),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_824),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_818),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_921),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_818),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_951),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_991),
.Y(n_1069)
);

CKINVDCx16_ASAP7_75t_R g1070 ( 
.A(n_928),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_818),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_818),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_818),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_980),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_980),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_779),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_980),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_980),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_781),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_785),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_980),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_737),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_787),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_790),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_794),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_737),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_737),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_743),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_718),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_778),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_798),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_817),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_800),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_827),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_748),
.Y(n_1095)
);

BUFx10_ASAP7_75t_L g1096 ( 
.A(n_802),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_881),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_900),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_816),
.B(n_1),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_719),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_942),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_965),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_801),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_768),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_826),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_718),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_805),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_928),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_807),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_815),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_718),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_998),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1015),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_788),
.Y(n_1114)
);

BUFx10_ASAP7_75t_L g1115 ( 
.A(n_718),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_829),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_826),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_791),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_791),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_878),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_718),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_753),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_799),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_808),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_833),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_878),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_888),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_825),
.Y(n_1128)
);

BUFx5_ASAP7_75t_L g1129 ( 
.A(n_712),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_888),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_924),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_753),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_753),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_924),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_935),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_959),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_828),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_959),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_928),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1028),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_753),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_884),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_1042),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_832),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_753),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1028),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_775),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1043),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1043),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_843),
.Y(n_1151)
);

BUFx5_ASAP7_75t_L g1152 ( 
.A(n_713),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_892),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_849),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_810),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_775),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_775),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_775),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_858),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_867),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_719),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_775),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_809),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_809),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_963),
.B(n_1),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_869),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_809),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_887),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_835),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1042),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_893),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_890),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_902),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_903),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_914),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_907),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_809),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_812),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_809),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_871),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_912),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_871),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_871),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_814),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_871),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_871),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_938),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_734),
.B(n_1),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_916),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_916),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_916),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_821),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_916),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_925),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_916),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_941),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_992),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_992),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_937),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_734),
.B(n_2),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_948),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_992),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_992),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_992),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_994),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_943),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_994),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_994),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_994),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_1042),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_947),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_994),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_751),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_746),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_751),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_840),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_957),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_968),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_840),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_962),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_983),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_953),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_953),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_715),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_757),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_723),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_732),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_733),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_730),
.B(n_3),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_822),
.Y(n_1230)
);

BUFx5_ASAP7_75t_L g1231 ( 
.A(n_744),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_752),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_752),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_755),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_834),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_836),
.Y(n_1236)
);

INVxp33_ASAP7_75t_SL g1237 ( 
.A(n_746),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_837),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_765),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_986),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_771),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_987),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_780),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_782),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_783),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_789),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_793),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_839),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_844),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_847),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_848),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_792),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_757),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_792),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_795),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_757),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_806),
.Y(n_1257)
);

BUFx2_ASAP7_75t_SL g1258 ( 
.A(n_786),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_819),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_851),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_786),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_823),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1004),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_830),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_838),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_841),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_786),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_855),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_845),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_846),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_856),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_813),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_850),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_852),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_864),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_873),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_886),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_857),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_894),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_897),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_859),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_860),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_904),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_854),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_909),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_910),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_911),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_854),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_913),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_927),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_929),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_944),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_861),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_854),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_863),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_952),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_956),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_970),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_796),
.B(n_2),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_960),
.Y(n_1300)
);

BUFx5_ASAP7_75t_L g1301 ( 
.A(n_961),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_813),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_970),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_966),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_865),
.Y(n_1305)
);

CKINVDCx14_ASAP7_75t_R g1306 ( 
.A(n_970),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_967),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_804),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_866),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_868),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_870),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_872),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_988),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_875),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_820),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1006),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1013),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_876),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1018),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1007),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_877),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_880),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1014),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1019),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_820),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_882),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1030),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1037),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1017),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_883),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_885),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1039),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1044),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_831),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_895),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_896),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_831),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_862),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_862),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_891),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1029),
.Y(n_1341)
);

INVxp33_ASAP7_75t_L g1342 ( 
.A(n_891),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_923),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_898),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_899),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_923),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_933),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_901),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_933),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_977),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_905),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_977),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_906),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_984),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_796),
.B(n_2),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1031),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_908),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_747),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_915),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_984),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_917),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1020),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_918),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1020),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_811),
.Y(n_1365)
);

BUFx8_ASAP7_75t_SL g1366 ( 
.A(n_747),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_776),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_811),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_853),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_853),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_776),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_919),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_972),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1001),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_920),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_874),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_990),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_874),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_922),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_922),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_926),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_930),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_931),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_932),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_934),
.Y(n_1385)
);

CKINVDCx14_ASAP7_75t_R g1386 ( 
.A(n_1001),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_936),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_939),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_945),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1012),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_946),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_949),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_954),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_958),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_964),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_969),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_971),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_974),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_975),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_976),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1012),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_978),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_981),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1016),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_982),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_985),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_995),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_996),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1230),
.B(n_1016),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1122),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1183),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1060),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1062),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1408),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1235),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1066),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1063),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1095),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1065),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1067),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1071),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1072),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_1236),
.B(n_1238),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1248),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1095),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1249),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_L g1427 ( 
.A(n_1250),
.B(n_3),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1251),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1381),
.B(n_1034),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1260),
.Y(n_1430)
);

INVxp33_ASAP7_75t_SL g1431 ( 
.A(n_1054),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1104),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1073),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1268),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1104),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1077),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1078),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1106),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1116),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1271),
.B(n_1034),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1081),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1116),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1278),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1125),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1156),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1281),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1157),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1162),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1408),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1282),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1163),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1293),
.B(n_4),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1164),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1167),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1177),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1179),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1180),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1059),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1182),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1185),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1045),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1061),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1045),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1366),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1366),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1125),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1186),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1295),
.B(n_4),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1191),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1193),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1305),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1161),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1382),
.B(n_1035),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1195),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1309),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1310),
.Y(n_1476)
);

INVxp33_ASAP7_75t_SL g1477 ( 
.A(n_1066),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1384),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1311),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1384),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1106),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1169),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1312),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1394),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1314),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1198),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1202),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1203),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1204),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1205),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1383),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1207),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1106),
.Y(n_1493)
);

INVxp33_ASAP7_75t_SL g1494 ( 
.A(n_1068),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1209),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1169),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1385),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1176),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1212),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1059),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1074),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1074),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1389),
.B(n_5),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1392),
.B(n_5),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1395),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1176),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1187),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1402),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1187),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1196),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1075),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1196),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1075),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1403),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1240),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1158),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1158),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1258),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1339),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1082),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1373),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1405),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1240),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1406),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1407),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1377),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1086),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1046),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1046),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1087),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1242),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1068),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_R g1533 ( 
.A(n_1114),
.B(n_1035),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1394),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1123),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1124),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_L g1537 ( 
.A(n_1128),
.B(n_6),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1089),
.B(n_1041),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1356),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1138),
.Y(n_1540)
);

NOR2xp67_ASAP7_75t_L g1541 ( 
.A(n_1145),
.B(n_6),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1151),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1154),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1058),
.B(n_709),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1061),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1400),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1061),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1400),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1242),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1106),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1263),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1159),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1160),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1166),
.B(n_709),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1133),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1168),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1263),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1171),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1089),
.Y(n_1559)
);

INVxp33_ASAP7_75t_SL g1560 ( 
.A(n_1173),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1111),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1174),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1175),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1323),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1194),
.B(n_711),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1323),
.Y(n_1566)
);

NOR2xp67_ASAP7_75t_L g1567 ( 
.A(n_1199),
.B(n_7),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1206),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1111),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1121),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1387),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1211),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1217),
.B(n_711),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1220),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1121),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1132),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1132),
.Y(n_1577)
);

CKINVDCx16_ASAP7_75t_R g1578 ( 
.A(n_1064),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1146),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1388),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1329),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1146),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1221),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1386),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1148),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1386),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1076),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1148),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1189),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_L g1590 ( 
.A(n_1076),
.B(n_7),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1189),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1079),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1329),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1190),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1069),
.B(n_721),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_L g1596 ( 
.A(n_1079),
.B(n_7),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1341),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1341),
.Y(n_1598)
);

NOR2xp67_ASAP7_75t_L g1599 ( 
.A(n_1080),
.B(n_8),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1391),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1190),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_R g1602 ( 
.A(n_1080),
.B(n_716),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1197),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1049),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1393),
.B(n_716),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1083),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1197),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1049),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1083),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1115),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1084),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1100),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1133),
.Y(n_1613)
);

CKINVDCx16_ASAP7_75t_R g1614 ( 
.A(n_1306),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1084),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1115),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1115),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1358),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1085),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1117),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1214),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1085),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1396),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1224),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1226),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1091),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1091),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1093),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1093),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1103),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1397),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1103),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1227),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1107),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1228),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1398),
.B(n_717),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1358),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1234),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1107),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1239),
.Y(n_1640)
);

CKINVDCx16_ASAP7_75t_R g1641 ( 
.A(n_1306),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1399),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1109),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1109),
.B(n_8),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1241),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1178),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1243),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1178),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1147),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1367),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1184),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1244),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1184),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1192),
.B(n_717),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1245),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1367),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1192),
.Y(n_1657)
);

CKINVDCx14_ASAP7_75t_R g1658 ( 
.A(n_1371),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1371),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1147),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1246),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1247),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1255),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1401),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1257),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1401),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1133),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1318),
.Y(n_1668)
);

CKINVDCx16_ASAP7_75t_R g1669 ( 
.A(n_1070),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1374),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1259),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1262),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1264),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1265),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1318),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1266),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1105),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1269),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1321),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1322),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1326),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1326),
.B(n_720),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1270),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1105),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1273),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1274),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1330),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1404),
.Y(n_1689)
);

CKINVDCx16_ASAP7_75t_R g1690 ( 
.A(n_1108),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1330),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1275),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1276),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1201),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1277),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1279),
.Y(n_1696)
);

INVxp33_ASAP7_75t_SL g1697 ( 
.A(n_1331),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1280),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1331),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1283),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1335),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1285),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1335),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1286),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1287),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1336),
.B(n_720),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1336),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1289),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1344),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1404),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1140),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_1144),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1290),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1308),
.B(n_722),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1458),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1478),
.B(n_1133),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1620),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1493),
.Y(n_1718)
);

OA21x2_ASAP7_75t_L g1719 ( 
.A1(n_1445),
.A2(n_1048),
.B(n_1047),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1521),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1544),
.A2(n_1165),
.B1(n_1099),
.B2(n_1237),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1493),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1458),
.Y(n_1723)
);

OA21x2_ASAP7_75t_L g1724 ( 
.A1(n_1447),
.A2(n_1052),
.B(n_1050),
.Y(n_1724)
);

XNOR2xp5_ASAP7_75t_L g1725 ( 
.A(n_1418),
.B(n_1218),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1559),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1526),
.B(n_1252),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1561),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1624),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1625),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1633),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1569),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1614),
.B(n_1344),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1480),
.B(n_1484),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1570),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1571),
.A2(n_1237),
.B1(n_1143),
.B2(n_1110),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1534),
.B(n_1252),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1546),
.B(n_1342),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1635),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1462),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1641),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1638),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1493),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1548),
.B(n_1142),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1575),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1462),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1493),
.Y(n_1747)
);

AND2x2_ASAP7_75t_SL g1748 ( 
.A(n_1646),
.B(n_1299),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1576),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1516),
.B(n_1232),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1577),
.Y(n_1751)
);

AND2x6_ASAP7_75t_L g1752 ( 
.A(n_1545),
.B(n_1053),
.Y(n_1752)
);

CKINVDCx11_ASAP7_75t_R g1753 ( 
.A(n_1604),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1580),
.B(n_1142),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1640),
.Y(n_1755)
);

INVx5_ASAP7_75t_L g1756 ( 
.A(n_1438),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1645),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1579),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1595),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1600),
.B(n_1142),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1438),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1647),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1582),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1652),
.Y(n_1764)
);

CKINVDCx16_ASAP7_75t_R g1765 ( 
.A(n_1578),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1655),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1538),
.B(n_1342),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1623),
.B(n_1142),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1585),
.Y(n_1769)
);

INVx6_ASAP7_75t_L g1770 ( 
.A(n_1538),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1538),
.B(n_1232),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1631),
.B(n_1208),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1588),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1661),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1517),
.B(n_1233),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1642),
.A2(n_1153),
.B1(n_1088),
.B2(n_1345),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1602),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1429),
.A2(n_1345),
.B1(n_1351),
.B2(n_1348),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1589),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1662),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1410),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1438),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1694),
.B(n_1155),
.Y(n_1783)
);

BUFx8_ASAP7_75t_L g1784 ( 
.A(n_1547),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1663),
.Y(n_1785)
);

AOI22x1_ASAP7_75t_SL g1786 ( 
.A1(n_1604),
.A2(n_722),
.B1(n_725),
.B2(n_724),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1481),
.Y(n_1787)
);

AND2x2_ASAP7_75t_SL g1788 ( 
.A(n_1676),
.B(n_1229),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1649),
.B(n_1233),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1660),
.B(n_1272),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1591),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1473),
.A2(n_1351),
.B1(n_1353),
.B2(n_1348),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1594),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1481),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1520),
.B(n_1272),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1481),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1678),
.B(n_1325),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1448),
.A2(n_1056),
.B(n_1055),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1685),
.B(n_1325),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1411),
.B(n_1353),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1665),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1550),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1533),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1601),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1414),
.A2(n_1359),
.B1(n_1361),
.B2(n_1357),
.Y(n_1805)
);

CKINVDCx8_ASAP7_75t_R g1806 ( 
.A(n_1689),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1550),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1449),
.A2(n_1359),
.B1(n_1361),
.B2(n_1357),
.Y(n_1808)
);

OAI22x1_ASAP7_75t_L g1809 ( 
.A1(n_1612),
.A2(n_1172),
.B1(n_1181),
.B2(n_1170),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1555),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1671),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1672),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1605),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1636),
.A2(n_1057),
.B(n_1360),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1451),
.A2(n_1360),
.B(n_1119),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1519),
.B(n_1610),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1409),
.B(n_1363),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1673),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1616),
.B(n_1208),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1603),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1621),
.A2(n_1372),
.B1(n_1375),
.B2(n_1363),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1527),
.B(n_1291),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1555),
.Y(n_1823)
);

INVx4_ASAP7_75t_L g1824 ( 
.A(n_1613),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1607),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1500),
.Y(n_1826)
);

OA21x2_ASAP7_75t_L g1827 ( 
.A1(n_1453),
.A2(n_1120),
.B(n_1118),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1501),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1670),
.A2(n_1375),
.B1(n_1372),
.B2(n_1200),
.Y(n_1829)
);

AOI22x1_ASAP7_75t_SL g1830 ( 
.A1(n_1608),
.A2(n_724),
.B1(n_726),
.B2(n_725),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1674),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1677),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1613),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1667),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1679),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1684),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1686),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1454),
.A2(n_1127),
.B(n_1126),
.Y(n_1838)
);

AOI22x1_ASAP7_75t_SL g1839 ( 
.A1(n_1608),
.A2(n_726),
.B1(n_728),
.B2(n_727),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1687),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1617),
.B(n_1208),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1667),
.A2(n_1315),
.B(n_1365),
.Y(n_1842)
);

AOI22x1_ASAP7_75t_SL g1843 ( 
.A1(n_1464),
.A2(n_727),
.B1(n_729),
.B2(n_728),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1455),
.Y(n_1844)
);

NOR2x1_ASAP7_75t_L g1845 ( 
.A(n_1423),
.B(n_1225),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1412),
.B(n_1208),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1692),
.Y(n_1847)
);

AND2x6_ASAP7_75t_L g1848 ( 
.A(n_1530),
.B(n_1355),
.Y(n_1848)
);

INVx4_ASAP7_75t_L g1849 ( 
.A(n_1456),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1461),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1693),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1427),
.B(n_1452),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1468),
.B(n_1210),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1695),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1457),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1696),
.B(n_1698),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1459),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1700),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1461),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1502),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1440),
.A2(n_1390),
.B1(n_1303),
.B2(n_1284),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1460),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1467),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1702),
.B(n_1292),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1463),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1704),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1705),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1714),
.A2(n_1188),
.B1(n_1303),
.B2(n_1288),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1511),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1708),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1713),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1513),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1413),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1417),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1419),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1503),
.B(n_1296),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1504),
.B(n_1297),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1420),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1421),
.B(n_1379),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1422),
.B(n_1051),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1433),
.B(n_1379),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1436),
.B(n_1379),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1437),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1441),
.B(n_1051),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1469),
.B(n_1379),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1654),
.A2(n_1294),
.B1(n_1298),
.B2(n_1253),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1560),
.B(n_1320),
.Y(n_1887)
);

CKINVDCx16_ASAP7_75t_R g1888 ( 
.A(n_1669),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1711),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1683),
.A2(n_797),
.B1(n_842),
.B2(n_784),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1706),
.A2(n_1518),
.B1(n_1565),
.B2(n_1554),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1470),
.Y(n_1892)
);

INVx5_ASAP7_75t_L g1893 ( 
.A(n_1474),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1573),
.A2(n_889),
.B1(n_973),
.B2(n_879),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1486),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1487),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1488),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1489),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1490),
.B(n_1051),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1492),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1495),
.B(n_1130),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1499),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1574),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1535),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1584),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1590),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1596),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1599),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1586),
.Y(n_1909)
);

CKINVDCx8_ASAP7_75t_R g1910 ( 
.A(n_1539),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1592),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1627),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1415),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1651),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1644),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1560),
.B(n_1225),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1536),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1675),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1537),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1472),
.B(n_1131),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1541),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1567),
.B(n_1134),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1691),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1707),
.B(n_1135),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1424),
.B(n_1136),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1416),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1426),
.B(n_1051),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1532),
.A2(n_1315),
.B(n_1365),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1463),
.B(n_1300),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1697),
.A2(n_1315),
.B(n_1368),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1587),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1606),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1609),
.Y(n_1933)
);

BUFx12f_ASAP7_75t_L g1934 ( 
.A(n_1464),
.Y(n_1934)
);

CKINVDCx16_ASAP7_75t_R g1935 ( 
.A(n_1690),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1611),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1615),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1428),
.B(n_1304),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1430),
.B(n_1051),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1434),
.B(n_1307),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1443),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1446),
.B(n_1137),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1697),
.A2(n_993),
.B1(n_1002),
.B2(n_979),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1619),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1450),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1475),
.B(n_1051),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1476),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1479),
.B(n_1139),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1483),
.B(n_1051),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1485),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1711),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1491),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1497),
.Y(n_1953)
);

XNOR2x2_ASAP7_75t_L g1954 ( 
.A(n_1431),
.B(n_1369),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1505),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1508),
.B(n_1129),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1514),
.A2(n_729),
.B1(n_735),
.B2(n_731),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1522),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1668),
.Y(n_1959)
);

BUFx8_ASAP7_75t_L g1960 ( 
.A(n_1658),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1540),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1524),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1680),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1542),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1525),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1543),
.A2(n_731),
.B1(n_736),
.B2(n_735),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1681),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1552),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1682),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1553),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1556),
.Y(n_1971)
);

AO22x2_ASAP7_75t_L g1972 ( 
.A1(n_1622),
.A2(n_1370),
.B1(n_1380),
.B2(n_1376),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1562),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1477),
.A2(n_736),
.B1(n_739),
.B2(n_738),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1688),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1558),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1563),
.Y(n_1977)
);

OAI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1477),
.A2(n_1378),
.B(n_1368),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1568),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1572),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1583),
.Y(n_1981)
);

BUFx12f_ASAP7_75t_L g1982 ( 
.A(n_1465),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1471),
.Y(n_1983)
);

INVx5_ASAP7_75t_L g1984 ( 
.A(n_1471),
.Y(n_1984)
);

CKINVDCx11_ASAP7_75t_R g1985 ( 
.A(n_1418),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1699),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1562),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1701),
.Y(n_1988)
);

OAI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1494),
.A2(n_1378),
.B(n_1149),
.Y(n_1989)
);

OAI22x1_ASAP7_75t_L g1990 ( 
.A1(n_1622),
.A2(n_738),
.B1(n_740),
.B2(n_739),
.Y(n_1990)
);

AND2x6_ASAP7_75t_L g1991 ( 
.A(n_1494),
.B(n_1256),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1626),
.B(n_1256),
.Y(n_1992)
);

INVxp33_ASAP7_75t_SL g1993 ( 
.A(n_1626),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1709),
.B(n_1129),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1628),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1628),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1431),
.A2(n_740),
.B1(n_742),
.B2(n_741),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1629),
.B(n_1141),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1629),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1630),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1712),
.A2(n_741),
.B1(n_745),
.B2(n_742),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1630),
.B(n_1129),
.Y(n_2002)
);

AOI22x1_ASAP7_75t_SL g2003 ( 
.A1(n_1465),
.A2(n_745),
.B1(n_750),
.B2(n_749),
.Y(n_2003)
);

AO22x2_ASAP7_75t_L g2004 ( 
.A1(n_1721),
.A2(n_1261),
.B1(n_1267),
.B2(n_714),
.Y(n_2004)
);

BUFx10_ASAP7_75t_L g2005 ( 
.A(n_1817),
.Y(n_2005)
);

OAI22xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1770),
.A2(n_1813),
.B1(n_1907),
.B2(n_1906),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1813),
.A2(n_1634),
.B1(n_1639),
.B2(n_1632),
.Y(n_2007)
);

OAI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1770),
.A2(n_1632),
.B1(n_1639),
.B2(n_1634),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1727),
.B(n_1643),
.Y(n_2009)
);

OAI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1770),
.A2(n_1643),
.B1(n_1653),
.B2(n_1648),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1715),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1715),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1842),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1788),
.A2(n_1653),
.B1(n_1657),
.B2(n_1648),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1842),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1788),
.A2(n_1703),
.B1(n_1657),
.B2(n_1529),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1890),
.A2(n_1703),
.B1(n_1528),
.B2(n_1267),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_SL g2018 ( 
.A1(n_1908),
.A2(n_750),
.B1(n_756),
.B2(n_749),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1789),
.B(n_1090),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1750),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1723),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1748),
.A2(n_1528),
.B1(n_1152),
.B2(n_1231),
.Y(n_2022)
);

AO22x2_ASAP7_75t_L g2023 ( 
.A1(n_1736),
.A2(n_1261),
.B1(n_1150),
.B2(n_1313),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1734),
.B(n_1129),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1723),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1734),
.A2(n_1152),
.B1(n_1231),
.B2(n_1129),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1748),
.A2(n_1152),
.B1(n_1231),
.B2(n_1129),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_SL g2028 ( 
.A1(n_1725),
.A2(n_1637),
.B1(n_1650),
.B2(n_1618),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1815),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_SL g2030 ( 
.A1(n_2001),
.A2(n_1637),
.B1(n_1650),
.B2(n_1618),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1815),
.Y(n_2031)
);

OR2x6_ASAP7_75t_L g2032 ( 
.A(n_1720),
.B(n_1092),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1727),
.B(n_1096),
.Y(n_2033)
);

OAI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1894),
.A2(n_758),
.B1(n_759),
.B2(n_756),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1815),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1737),
.B(n_1096),
.Y(n_2036)
);

AOI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1848),
.A2(n_1152),
.B1(n_1231),
.B2(n_1129),
.Y(n_2037)
);

OA22x2_ASAP7_75t_L g2038 ( 
.A1(n_1943),
.A2(n_772),
.B1(n_1008),
.B2(n_761),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1726),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1783),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1767),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1777),
.B(n_1096),
.Y(n_2042)
);

OAI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1759),
.A2(n_759),
.B1(n_760),
.B2(n_758),
.Y(n_2043)
);

OAI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_2002),
.A2(n_761),
.B1(n_762),
.B2(n_760),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_SL g2045 ( 
.A1(n_1997),
.A2(n_1659),
.B1(n_1664),
.B2(n_1656),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1817),
.B(n_1712),
.Y(n_2046)
);

OAI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1915),
.A2(n_763),
.B1(n_764),
.B2(n_762),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_SL g2048 ( 
.A1(n_1993),
.A2(n_1659),
.B1(n_1664),
.B2(n_1656),
.Y(n_2048)
);

OR2x6_ASAP7_75t_L g2049 ( 
.A(n_1913),
.B(n_1094),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1737),
.B(n_1097),
.Y(n_2050)
);

AND2x2_ASAP7_75t_SL g2051 ( 
.A(n_1887),
.B(n_1098),
.Y(n_2051)
);

OAI22xp33_ASAP7_75t_SL g2052 ( 
.A1(n_1921),
.A2(n_764),
.B1(n_766),
.B2(n_763),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1738),
.B(n_1101),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1738),
.B(n_1102),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1848),
.B(n_1152),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1726),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1848),
.A2(n_1231),
.B1(n_1301),
.B2(n_1152),
.Y(n_2057)
);

OAI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1994),
.A2(n_767),
.B1(n_769),
.B2(n_766),
.Y(n_2058)
);

OAI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1852),
.A2(n_769),
.B1(n_770),
.B2(n_767),
.Y(n_2059)
);

OAI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1816),
.A2(n_772),
.B1(n_773),
.B2(n_770),
.Y(n_2060)
);

OAI22xp33_ASAP7_75t_SL g2061 ( 
.A1(n_1852),
.A2(n_774),
.B1(n_997),
.B2(n_773),
.Y(n_2061)
);

OAI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1781),
.A2(n_997),
.B1(n_999),
.B2(n_774),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1767),
.B(n_1112),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1728),
.Y(n_2064)
);

AND2x4_ASAP7_75t_SL g2065 ( 
.A(n_1913),
.B(n_1425),
.Y(n_2065)
);

OAI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1781),
.A2(n_1000),
.B1(n_1003),
.B2(n_999),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1930),
.Y(n_2067)
);

AO22x2_ASAP7_75t_L g2068 ( 
.A1(n_1776),
.A2(n_1316),
.B1(n_1319),
.B2(n_1317),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1728),
.Y(n_2069)
);

OAI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1861),
.A2(n_1003),
.B1(n_1005),
.B2(n_1000),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1920),
.B(n_1113),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1732),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1750),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1920),
.B(n_1338),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1732),
.Y(n_2075)
);

AOI22x1_ASAP7_75t_L g2076 ( 
.A1(n_1990),
.A2(n_1008),
.B1(n_1009),
.B2(n_1005),
.Y(n_2076)
);

NAND2xp33_ASAP7_75t_SL g2077 ( 
.A(n_1996),
.B(n_1009),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_1966),
.B(n_1324),
.Y(n_2078)
);

OA22x2_ASAP7_75t_L g2079 ( 
.A1(n_1990),
.A2(n_1886),
.B1(n_1974),
.B2(n_1957),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1891),
.B(n_1800),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1848),
.A2(n_1231),
.B1(n_1301),
.B2(n_1152),
.Y(n_2081)
);

BUFx10_ASAP7_75t_L g2082 ( 
.A(n_1916),
.Y(n_2082)
);

OAI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1927),
.A2(n_1011),
.B1(n_1021),
.B2(n_1010),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1930),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1848),
.A2(n_1301),
.B1(n_1231),
.B2(n_1011),
.Y(n_2085)
);

OAI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_1939),
.A2(n_1021),
.B1(n_1022),
.B2(n_1010),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1946),
.A2(n_1023),
.B1(n_1024),
.B2(n_1022),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_SL g2088 ( 
.A(n_1996),
.B(n_1919),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1848),
.A2(n_1301),
.B1(n_1328),
.B2(n_1327),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1800),
.A2(n_1301),
.B1(n_1333),
.B2(n_1332),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_1924),
.B(n_1023),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1771),
.B(n_1922),
.Y(n_2092)
);

OAI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1853),
.A2(n_1025),
.B1(n_1026),
.B2(n_1024),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1771),
.B(n_1338),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1922),
.B(n_1213),
.Y(n_2095)
);

OAI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1949),
.A2(n_1026),
.B1(n_1027),
.B2(n_1025),
.Y(n_2096)
);

BUFx10_ASAP7_75t_L g2097 ( 
.A(n_1916),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1735),
.Y(n_2098)
);

AO22x2_ASAP7_75t_L g2099 ( 
.A1(n_1868),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1998),
.B(n_1924),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1998),
.B(n_1215),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_SL g2102 ( 
.A1(n_1853),
.A2(n_1032),
.B1(n_1033),
.B2(n_1027),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1803),
.B(n_1216),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1778),
.A2(n_1301),
.B1(n_1302),
.B2(n_1254),
.Y(n_2104)
);

INVx11_ASAP7_75t_L g2105 ( 
.A(n_1960),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1789),
.B(n_1219),
.Y(n_2106)
);

OAI22xp33_ASAP7_75t_SL g2107 ( 
.A1(n_1729),
.A2(n_1033),
.B1(n_1036),
.B2(n_1032),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1938),
.B(n_1222),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_1789),
.B(n_1223),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1956),
.A2(n_1038),
.B1(n_1040),
.B2(n_1036),
.Y(n_2110)
);

OR2x6_ASAP7_75t_L g2111 ( 
.A(n_1913),
.B(n_1334),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1792),
.A2(n_1301),
.B1(n_1302),
.B2(n_1254),
.Y(n_2112)
);

AND2x2_ASAP7_75t_SL g2113 ( 
.A(n_1996),
.B(n_1425),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1911),
.A2(n_1040),
.B1(n_1038),
.B2(n_1254),
.Y(n_2114)
);

AO22x2_ASAP7_75t_L g2115 ( 
.A1(n_1829),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_SL g2116 ( 
.A1(n_1993),
.A2(n_1710),
.B1(n_1666),
.B2(n_1435),
.Y(n_2116)
);

OAI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_1911),
.A2(n_1302),
.B1(n_1364),
.B2(n_1254),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_1925),
.A2(n_1364),
.B1(n_1302),
.B2(n_1340),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1790),
.B(n_1337),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1938),
.B(n_1343),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_SL g2121 ( 
.A1(n_1765),
.A2(n_1710),
.B1(n_1666),
.B2(n_1435),
.Y(n_2121)
);

OAI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1912),
.A2(n_1364),
.B1(n_1347),
.B2(n_1349),
.Y(n_2122)
);

OA22x2_ASAP7_75t_L g2123 ( 
.A1(n_1809),
.A2(n_1350),
.B1(n_1352),
.B2(n_1346),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1925),
.A2(n_1364),
.B1(n_1362),
.B2(n_1354),
.Y(n_2124)
);

INVx8_ASAP7_75t_L g2125 ( 
.A(n_1991),
.Y(n_2125)
);

BUFx10_ASAP7_75t_L g2126 ( 
.A(n_1850),
.Y(n_2126)
);

OAI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1912),
.A2(n_1439),
.B1(n_1442),
.B2(n_1432),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1735),
.Y(n_2128)
);

OAI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1914),
.A2(n_1918),
.B1(n_1731),
.B2(n_1739),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_SL g2130 ( 
.A1(n_1973),
.A2(n_1439),
.B1(n_1442),
.B2(n_1432),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1938),
.B(n_1549),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_1942),
.A2(n_1466),
.B1(n_1482),
.B2(n_1444),
.Y(n_2132)
);

AO22x2_ASAP7_75t_L g2133 ( 
.A1(n_1821),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_2133)
);

OAI22xp33_ASAP7_75t_SL g2134 ( 
.A1(n_1730),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2134)
);

OAI22xp33_ASAP7_75t_SL g2135 ( 
.A1(n_1742),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1942),
.A2(n_1466),
.B1(n_1482),
.B2(n_1444),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1940),
.B(n_1597),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1948),
.A2(n_1940),
.B1(n_1856),
.B2(n_1797),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_1948),
.A2(n_1498),
.B1(n_1506),
.B2(n_1496),
.Y(n_2139)
);

AO22x2_ASAP7_75t_L g2140 ( 
.A1(n_1786),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1940),
.B(n_1598),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1790),
.B(n_14),
.Y(n_2142)
);

NAND3x1_ASAP7_75t_L g2143 ( 
.A(n_1999),
.B(n_1498),
.C(n_1496),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_SL g2144 ( 
.A1(n_1973),
.A2(n_1507),
.B1(n_1509),
.B2(n_1506),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1856),
.A2(n_1509),
.B1(n_1510),
.B2(n_1507),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1914),
.B(n_1523),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1745),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1745),
.Y(n_2148)
);

BUFx10_ASAP7_75t_L g2149 ( 
.A(n_1850),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1918),
.A2(n_1512),
.B1(n_1515),
.B2(n_1510),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_SL g2151 ( 
.A1(n_1888),
.A2(n_1515),
.B1(n_1523),
.B2(n_1512),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1856),
.A2(n_1549),
.B1(n_1551),
.B2(n_1531),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1903),
.B(n_1564),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_1876),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_SL g2155 ( 
.A1(n_1935),
.A2(n_1551),
.B1(n_1557),
.B2(n_1531),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_1790),
.A2(n_1564),
.B1(n_1566),
.B2(n_1557),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1984),
.B(n_1597),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1797),
.B(n_15),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1749),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1749),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_1992),
.B(n_17),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1751),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_R g2163 ( 
.A(n_1910),
.B(n_1566),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_1755),
.A2(n_1593),
.B1(n_1598),
.B2(n_1581),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1750),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_1797),
.A2(n_1799),
.B1(n_1972),
.B2(n_1864),
.Y(n_2166)
);

INVx5_ASAP7_75t_L g2167 ( 
.A(n_1991),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1903),
.B(n_1581),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1984),
.B(n_1593),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1751),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1758),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1758),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1763),
.Y(n_2173)
);

AO22x2_ASAP7_75t_L g2174 ( 
.A1(n_1830),
.A2(n_1839),
.B1(n_2000),
.B2(n_1808),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1763),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1769),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1983),
.B(n_696),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_1805),
.B(n_17),
.Y(n_2178)
);

NAND2xp33_ASAP7_75t_SL g2179 ( 
.A(n_1996),
.B(n_1986),
.Y(n_2179)
);

AO22x2_ASAP7_75t_L g2180 ( 
.A1(n_1983),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1905),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2181)
);

OAI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_1757),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1987),
.B(n_700),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1775),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1769),
.Y(n_2185)
);

AOI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_1799),
.A2(n_134),
.B1(n_135),
.B2(n_133),
.Y(n_2186)
);

AOI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_1799),
.A2(n_134),
.B1(n_135),
.B2(n_133),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_1762),
.A2(n_137),
.B1(n_138),
.B2(n_136),
.Y(n_2188)
);

NAND3x1_ASAP7_75t_L g2189 ( 
.A(n_1917),
.B(n_20),
.C(n_22),
.Y(n_2189)
);

OAI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_1764),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1773),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1871),
.B(n_22),
.Y(n_2192)
);

OAI22xp33_ASAP7_75t_SL g2193 ( 
.A1(n_1766),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_1775),
.Y(n_2194)
);

AOI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_1774),
.A2(n_137),
.B1(n_138),
.B2(n_136),
.Y(n_2195)
);

OAI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_1780),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1754),
.B(n_25),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1987),
.B(n_695),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_1871),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_1898),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1905),
.B(n_26),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1876),
.B(n_696),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_1785),
.A2(n_140),
.B1(n_141),
.B2(n_139),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1801),
.A2(n_142),
.B1(n_143),
.B2(n_139),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1876),
.B(n_700),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1773),
.Y(n_2206)
);

OA22x2_ASAP7_75t_L g2207 ( 
.A1(n_1809),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2207)
);

OR2x6_ASAP7_75t_L g2208 ( 
.A(n_1913),
.B(n_27),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1972),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1779),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1877),
.B(n_703),
.Y(n_2211)
);

OAI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_1811),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1779),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1984),
.B(n_30),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1984),
.B(n_30),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1791),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1877),
.B(n_706),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1791),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1793),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1793),
.Y(n_2220)
);

AOI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_1812),
.A2(n_143),
.B1(n_146),
.B2(n_142),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_1818),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2222)
);

OAI22xp33_ASAP7_75t_SL g2223 ( 
.A1(n_1831),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_1832),
.A2(n_148),
.B1(n_149),
.B2(n_147),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1835),
.A2(n_148),
.B1(n_150),
.B2(n_147),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1804),
.Y(n_2226)
);

AO22x2_ASAP7_75t_L g2227 ( 
.A1(n_1843),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_1909),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1804),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1820),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_1972),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1984),
.B(n_36),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_1836),
.A2(n_151),
.B1(n_152),
.B2(n_150),
.Y(n_2233)
);

OA22x2_ASAP7_75t_L g2234 ( 
.A1(n_1923),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1909),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1877),
.B(n_706),
.Y(n_2236)
);

OAI22xp33_ASAP7_75t_SL g2237 ( 
.A1(n_1837),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1840),
.A2(n_153),
.B1(n_154),
.B2(n_151),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1820),
.Y(n_2239)
);

AO22x2_ASAP7_75t_L g2240 ( 
.A1(n_2003),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1847),
.A2(n_156),
.B1(n_157),
.B2(n_154),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1760),
.B(n_43),
.Y(n_2242)
);

OAI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1851),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1825),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_1854),
.A2(n_1858),
.B1(n_1867),
.B2(n_1866),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1849),
.B(n_44),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_1926),
.B(n_45),
.Y(n_2247)
);

OAI22xp33_ASAP7_75t_L g2248 ( 
.A1(n_1870),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1825),
.Y(n_2249)
);

AOI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_1991),
.A2(n_157),
.B1(n_158),
.B2(n_156),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1775),
.Y(n_2251)
);

OA22x2_ASAP7_75t_L g2252 ( 
.A1(n_1929),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1826),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1824),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1988),
.B(n_704),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_1824),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1988),
.B(n_704),
.Y(n_2257)
);

AO22x2_ASAP7_75t_L g2258 ( 
.A1(n_1931),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1826),
.Y(n_2259)
);

OAI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_1717),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1986),
.B(n_159),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_1991),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1828),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1986),
.B(n_685),
.Y(n_2264)
);

OAI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_1768),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1828),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1849),
.B(n_51),
.Y(n_2267)
);

AO22x2_ASAP7_75t_L g2268 ( 
.A1(n_1932),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_1941),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1860),
.Y(n_2270)
);

AO22x2_ASAP7_75t_L g2271 ( 
.A1(n_1933),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1860),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1986),
.B(n_692),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1917),
.B(n_692),
.Y(n_2274)
);

BUFx10_ASAP7_75t_L g2275 ( 
.A(n_1859),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_SL g2276 ( 
.A1(n_1889),
.A2(n_62),
.B1(n_70),
.B2(n_54),
.Y(n_2276)
);

AND2x2_ASAP7_75t_SL g2277 ( 
.A(n_1741),
.B(n_55),
.Y(n_2277)
);

INVx3_ASAP7_75t_L g2278 ( 
.A(n_1824),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1869),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_1941),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2280)
);

AO22x2_ASAP7_75t_L g2281 ( 
.A1(n_1936),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2281)
);

OAI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_1945),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2282)
);

OAI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_1945),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1869),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_1991),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_2285)
);

OAI22xp33_ASAP7_75t_SL g2286 ( 
.A1(n_1733),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_1917),
.B(n_684),
.Y(n_2287)
);

OAI22xp33_ASAP7_75t_SL g2288 ( 
.A1(n_1733),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1928),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_1953),
.Y(n_2290)
);

OR2x6_ASAP7_75t_L g2291 ( 
.A(n_1953),
.B(n_61),
.Y(n_2291)
);

AND2x2_ASAP7_75t_SL g2292 ( 
.A(n_1953),
.B(n_1955),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_1961),
.B(n_684),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1873),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_1849),
.B(n_61),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_1991),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1928),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1961),
.B(n_687),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1772),
.B(n_62),
.Y(n_2299)
);

OAI22xp33_ASAP7_75t_SL g2300 ( 
.A1(n_1937),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1961),
.B(n_689),
.Y(n_2301)
);

AO22x2_ASAP7_75t_L g2302 ( 
.A1(n_1944),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2302)
);

OAI22xp33_ASAP7_75t_SL g2303 ( 
.A1(n_1959),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1872),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_1716),
.B(n_67),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1976),
.B(n_695),
.Y(n_2306)
);

OAI22xp33_ASAP7_75t_SL g2307 ( 
.A1(n_1963),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1873),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1875),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_1898),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_1864),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_1976),
.B(n_699),
.Y(n_2312)
);

AO22x2_ASAP7_75t_L g2313 ( 
.A1(n_1967),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2313)
);

AO22x2_ASAP7_75t_L g2314 ( 
.A1(n_1975),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_1752),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_1807),
.Y(n_2316)
);

OR2x6_ASAP7_75t_L g2317 ( 
.A(n_1953),
.B(n_71),
.Y(n_2317)
);

OAI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_1947),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_1752),
.A2(n_167),
.B1(n_168),
.B2(n_166),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_1929),
.Y(n_2320)
);

AOI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_1752),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1744),
.B(n_72),
.Y(n_2322)
);

OAI22xp33_ASAP7_75t_SL g2323 ( 
.A1(n_1819),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1864),
.B(n_1822),
.Y(n_2324)
);

AO22x2_ASAP7_75t_L g2325 ( 
.A1(n_1954),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_2325)
);

INVx4_ASAP7_75t_L g2326 ( 
.A(n_2125),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2167),
.B(n_1955),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2316),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2080),
.A2(n_2178),
.B1(n_2041),
.B2(n_2092),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2029),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2254),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2290),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_2316),
.Y(n_2333)
);

INVx2_ASAP7_75t_SL g2334 ( 
.A(n_2074),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2029),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2031),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2040),
.B(n_1995),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2050),
.B(n_1976),
.Y(n_2338)
);

OR2x6_ASAP7_75t_SL g2339 ( 
.A(n_2150),
.B(n_1859),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2031),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2035),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2005),
.B(n_1947),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2053),
.B(n_1989),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2304),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_2254),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2142),
.A2(n_2158),
.B1(n_2267),
.B2(n_2246),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2035),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2142),
.A2(n_1752),
.B1(n_1978),
.B2(n_1989),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2013),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2054),
.B(n_1978),
.Y(n_2350)
);

NOR3xp33_ASAP7_75t_L g2351 ( 
.A(n_2164),
.B(n_1951),
.C(n_1969),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2100),
.B(n_1955),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2167),
.B(n_1955),
.Y(n_2353)
);

INVx4_ASAP7_75t_L g2354 ( 
.A(n_2125),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2304),
.Y(n_2355)
);

INVx4_ASAP7_75t_L g2356 ( 
.A(n_2167),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2024),
.B(n_1874),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2013),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2005),
.B(n_1950),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2015),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2020),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2020),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_2094),
.Y(n_2363)
);

INVx4_ASAP7_75t_L g2364 ( 
.A(n_2316),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2073),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2256),
.Y(n_2366)
);

BUFx10_ASAP7_75t_L g2367 ( 
.A(n_2042),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2158),
.A2(n_1752),
.B1(n_1895),
.B2(n_1883),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2073),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2036),
.B(n_1962),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_2165),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2015),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2098),
.Y(n_2373)
);

CKINVDCx20_ASAP7_75t_R g2374 ( 
.A(n_2121),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2098),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2256),
.Y(n_2376)
);

AOI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2009),
.A2(n_1752),
.B1(n_1952),
.B2(n_1950),
.Y(n_2377)
);

BUFx10_ASAP7_75t_L g2378 ( 
.A(n_2065),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2165),
.Y(n_2379)
);

INVx5_ASAP7_75t_L g2380 ( 
.A(n_2278),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2278),
.B(n_2095),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2184),
.Y(n_2382)
);

BUFx3_ASAP7_75t_L g2383 ( 
.A(n_2199),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2128),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2153),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2184),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2194),
.Y(n_2387)
);

XNOR2xp5_ASAP7_75t_L g2388 ( 
.A(n_2151),
.B(n_1865),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2128),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_2324),
.B(n_1740),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2194),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2295),
.A2(n_1897),
.B1(n_1878),
.B2(n_1896),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2163),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2063),
.B(n_1952),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2101),
.B(n_1958),
.Y(n_2395)
);

AND2x6_ASAP7_75t_L g2396 ( 
.A(n_2067),
.B(n_1962),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2251),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2292),
.B(n_1962),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2168),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2138),
.B(n_2022),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2251),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2067),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2159),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2159),
.Y(n_2404)
);

AO22x2_ASAP7_75t_L g2405 ( 
.A1(n_2265),
.A2(n_1965),
.B1(n_1968),
.B2(n_1958),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2162),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2162),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2172),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2172),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2173),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2084),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2173),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2091),
.B(n_1965),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2084),
.Y(n_2414)
);

INVx2_ASAP7_75t_SL g2415 ( 
.A(n_2019),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2175),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2071),
.B(n_1968),
.Y(n_2417)
);

INVx2_ASAP7_75t_SL g2418 ( 
.A(n_2019),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2006),
.B(n_1962),
.Y(n_2419)
);

INVx2_ASAP7_75t_SL g2420 ( 
.A(n_2120),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2289),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2289),
.Y(n_2422)
);

OAI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2166),
.A2(n_1971),
.B1(n_1977),
.B2(n_1970),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2146),
.B(n_1970),
.Y(n_2424)
);

NOR2x1p5_ASAP7_75t_L g2425 ( 
.A(n_2199),
.B(n_1904),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2119),
.B(n_1977),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2175),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2055),
.B(n_1971),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2033),
.B(n_1971),
.Y(n_2429)
);

INVx4_ASAP7_75t_L g2430 ( 
.A(n_2199),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2185),
.Y(n_2431)
);

AO22x2_ASAP7_75t_L g2432 ( 
.A1(n_2181),
.A2(n_1980),
.B1(n_1981),
.B2(n_1979),
.Y(n_2432)
);

OR2x2_ASAP7_75t_L g2433 ( 
.A(n_2161),
.B(n_1979),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2026),
.B(n_1971),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_2026),
.B(n_2200),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2119),
.B(n_1980),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2106),
.B(n_1981),
.Y(n_2437)
);

AND2x6_ASAP7_75t_L g2438 ( 
.A(n_2297),
.B(n_1845),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2108),
.B(n_1901),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2106),
.B(n_1901),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2200),
.B(n_2310),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2185),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2320),
.A2(n_1929),
.B1(n_1794),
.B2(n_1855),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2200),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2109),
.B(n_1964),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2216),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2310),
.B(n_1904),
.Y(n_2447)
);

INVx4_ASAP7_75t_L g2448 ( 
.A(n_2310),
.Y(n_2448)
);

AND2x6_ASAP7_75t_L g2449 ( 
.A(n_2297),
.B(n_1964),
.Y(n_2449)
);

INVx3_ASAP7_75t_L g2450 ( 
.A(n_2011),
.Y(n_2450)
);

OAI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2089),
.A2(n_1746),
.B1(n_1740),
.B2(n_1865),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2216),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2219),
.Y(n_2453)
);

BUFx2_ASAP7_75t_L g2454 ( 
.A(n_2131),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2324),
.Y(n_2455)
);

BUFx10_ASAP7_75t_L g2456 ( 
.A(n_2046),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2012),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2109),
.B(n_1875),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2082),
.B(n_1806),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2274),
.B(n_1806),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2287),
.B(n_1844),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2219),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2226),
.Y(n_2463)
);

OR2x2_ASAP7_75t_L g2464 ( 
.A(n_2156),
.B(n_2078),
.Y(n_2464)
);

INVx5_ASAP7_75t_L g2465 ( 
.A(n_2111),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2226),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2284),
.Y(n_2467)
);

INVx5_ASAP7_75t_L g2468 ( 
.A(n_2111),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2284),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2214),
.A2(n_1896),
.B1(n_1878),
.B2(n_1827),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_2103),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2021),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2215),
.A2(n_1827),
.B1(n_1838),
.B2(n_1872),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2154),
.A2(n_2293),
.B1(n_2301),
.B2(n_2298),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2082),
.B(n_1910),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2039),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2025),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2294),
.B(n_2308),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2032),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2056),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2064),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2069),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2309),
.B(n_1879),
.Y(n_2483)
);

INVx4_ASAP7_75t_L g2484 ( 
.A(n_2072),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2126),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2075),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2147),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2306),
.A2(n_1855),
.B1(n_1857),
.B2(n_1844),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2148),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2051),
.B(n_1746),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2160),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2097),
.B(n_1954),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2170),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2312),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2171),
.B(n_1879),
.Y(n_2495)
);

INVx2_ASAP7_75t_SL g2496 ( 
.A(n_2032),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2126),
.Y(n_2497)
);

INVx3_ASAP7_75t_L g2498 ( 
.A(n_2176),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2097),
.B(n_1753),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2191),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2027),
.B(n_1844),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2232),
.A2(n_1827),
.B1(n_1838),
.B2(n_1872),
.Y(n_2502)
);

INVx4_ASAP7_75t_L g2503 ( 
.A(n_2206),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2007),
.B(n_2014),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2210),
.B(n_1881),
.Y(n_2505)
);

AOI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_2079),
.A2(n_1838),
.B1(n_1855),
.B2(n_1844),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2049),
.B(n_1822),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2027),
.B(n_1855),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2008),
.B(n_1753),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2213),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2049),
.B(n_1822),
.Y(n_2511)
);

XNOR2xp5_ASAP7_75t_L g2512 ( 
.A(n_2155),
.B(n_1985),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2218),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2220),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2088),
.A2(n_1857),
.B1(n_1863),
.B2(n_1862),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2229),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_2230),
.Y(n_2517)
);

INVxp67_ASAP7_75t_SL g2518 ( 
.A(n_2239),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2244),
.B(n_1881),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2202),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2105),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2085),
.B(n_1857),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2249),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2179),
.A2(n_2166),
.B1(n_2257),
.B2(n_2255),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2085),
.B(n_1857),
.Y(n_2525)
);

BUFx4f_ASAP7_75t_L g2526 ( 
.A(n_2261),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2253),
.Y(n_2527)
);

AND2x6_ASAP7_75t_L g2528 ( 
.A(n_2250),
.B(n_1882),
.Y(n_2528)
);

OAI22xp33_ASAP7_75t_L g2529 ( 
.A1(n_2262),
.A2(n_1841),
.B1(n_1863),
.B2(n_1862),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2259),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2205),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2263),
.Y(n_2532)
);

INVxp33_ASAP7_75t_L g2533 ( 
.A(n_2130),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2010),
.B(n_2037),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2266),
.B(n_1882),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2211),
.A2(n_1863),
.B1(n_1892),
.B2(n_1862),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2270),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2272),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2279),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2016),
.B(n_1985),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2217),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2305),
.Y(n_2542)
);

NOR2x1p5_ASAP7_75t_L g2543 ( 
.A(n_2247),
.B(n_1934),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2017),
.B(n_1960),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_2127),
.B(n_1960),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2245),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2322),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2236),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2149),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2197),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2177),
.B(n_1885),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2057),
.B(n_1862),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2242),
.Y(n_2553)
);

OAI22xp33_ASAP7_75t_L g2554 ( 
.A1(n_2285),
.A2(n_1892),
.B1(n_1900),
.B2(n_1863),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2264),
.B(n_2273),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2299),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2123),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2252),
.Y(n_2558)
);

AND3x2_ASAP7_75t_L g2559 ( 
.A(n_2137),
.B(n_1885),
.C(n_1795),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2180),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2124),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2070),
.B(n_1934),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2129),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2183),
.B(n_1892),
.Y(n_2564)
);

NOR2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2141),
.B(n_1982),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2081),
.B(n_1892),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2198),
.A2(n_1902),
.B1(n_1900),
.B2(n_1719),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2180),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2058),
.B(n_1982),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2118),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2068),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2157),
.B(n_1795),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2093),
.B(n_1900),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2068),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2090),
.B(n_1900),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2149),
.Y(n_2576)
);

OR2x6_ASAP7_75t_L g2577 ( 
.A(n_2208),
.B(n_1814),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2044),
.B(n_1902),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2234),
.Y(n_2579)
);

NAND3xp33_ASAP7_75t_L g2580 ( 
.A(n_2201),
.B(n_1784),
.C(n_1902),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2104),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2083),
.B(n_1902),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2112),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2086),
.B(n_2087),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2189),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2192),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2122),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2258),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2023),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2275),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2023),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2258),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2096),
.B(n_2110),
.Y(n_2593)
);

INVxp67_ASAP7_75t_L g2594 ( 
.A(n_2114),
.Y(n_2594)
);

BUFx4f_ASAP7_75t_L g2595 ( 
.A(n_2113),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2296),
.Y(n_2596)
);

CKINVDCx20_ASAP7_75t_R g2597 ( 
.A(n_2028),
.Y(n_2597)
);

AND3x2_ASAP7_75t_L g2598 ( 
.A(n_2325),
.B(n_1784),
.C(n_75),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2275),
.B(n_2208),
.Y(n_2599)
);

INVx4_ASAP7_75t_L g2600 ( 
.A(n_2291),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2102),
.B(n_1807),
.Y(n_2601)
);

INVx5_ASAP7_75t_L g2602 ( 
.A(n_2291),
.Y(n_2602)
);

AND2x2_ASAP7_75t_SL g2603 ( 
.A(n_2311),
.B(n_1719),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2317),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2169),
.B(n_2059),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2268),
.Y(n_2606)
);

INVx2_ASAP7_75t_SL g2607 ( 
.A(n_2317),
.Y(n_2607)
);

AOI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2077),
.A2(n_1880),
.B1(n_1899),
.B2(n_1884),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2132),
.B(n_1719),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2186),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2187),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2268),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2061),
.B(n_1784),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2144),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2060),
.B(n_1787),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2228),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2271),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_L g2618 ( 
.A(n_2136),
.B(n_2139),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_2004),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2038),
.Y(n_2620)
);

BUFx10_ASAP7_75t_L g2621 ( 
.A(n_2277),
.Y(n_2621)
);

INVx4_ASAP7_75t_L g2622 ( 
.A(n_2271),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2281),
.Y(n_2623)
);

INVx5_ASAP7_75t_L g2624 ( 
.A(n_2315),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2004),
.B(n_1787),
.Y(n_2625)
);

NAND3xp33_ASAP7_75t_L g2626 ( 
.A(n_2076),
.B(n_1798),
.C(n_1724),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2207),
.B(n_1814),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2311),
.B(n_1724),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2286),
.B(n_1787),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2288),
.B(n_1807),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2281),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2302),
.Y(n_2632)
);

AND2x6_ASAP7_75t_L g2633 ( 
.A(n_2209),
.B(n_2231),
.Y(n_2633)
);

BUFx4f_ASAP7_75t_L g2634 ( 
.A(n_2323),
.Y(n_2634)
);

CKINVDCx16_ASAP7_75t_R g2635 ( 
.A(n_2116),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2319),
.B(n_1807),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2235),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2145),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_L g2639 ( 
.A(n_2321),
.B(n_1810),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2117),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2302),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2313),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2188),
.B(n_1802),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_2048),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2313),
.Y(n_2645)
);

NAND2xp33_ASAP7_75t_R g2646 ( 
.A(n_2143),
.B(n_1724),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2314),
.Y(n_2647)
);

INVx1_ASAP7_75t_SL g2648 ( 
.A(n_2152),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2174),
.B(n_1798),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2314),
.Y(n_2650)
);

NAND2x1_ASAP7_75t_L g2651 ( 
.A(n_2209),
.B(n_1802),
.Y(n_2651)
);

OR2x6_ASAP7_75t_L g2652 ( 
.A(n_2174),
.B(n_2325),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2062),
.B(n_1798),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2195),
.B(n_1802),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2115),
.Y(n_2655)
);

INVx5_ASAP7_75t_L g2656 ( 
.A(n_2134),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_2135),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2043),
.B(n_1810),
.Y(n_2658)
);

AO22x2_ASAP7_75t_L g2659 ( 
.A1(n_2133),
.A2(n_2231),
.B1(n_2115),
.B2(n_2099),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2066),
.B(n_1810),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2099),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2034),
.A2(n_1782),
.B1(n_1796),
.B2(n_1761),
.Y(n_2662)
);

INVx3_ASAP7_75t_L g2663 ( 
.A(n_2133),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2076),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2047),
.B(n_1810),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2193),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2269),
.B(n_1823),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2280),
.A2(n_1834),
.B1(n_1823),
.B2(n_1782),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2203),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_L g2670 ( 
.A(n_2018),
.B(n_1823),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2204),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2221),
.B(n_1833),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2224),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2225),
.Y(n_2674)
);

NAND2xp33_ASAP7_75t_L g2675 ( 
.A(n_2233),
.B(n_1834),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2238),
.B(n_1833),
.Y(n_2676)
);

AND3x2_ASAP7_75t_L g2677 ( 
.A(n_2276),
.B(n_76),
.C(n_77),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2241),
.Y(n_2678)
);

AOI22xp33_ASAP7_75t_L g2679 ( 
.A1(n_2282),
.A2(n_2318),
.B1(n_2283),
.B2(n_2190),
.Y(n_2679)
);

BUFx6f_ASAP7_75t_L g2680 ( 
.A(n_2223),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2237),
.Y(n_2681)
);

INVx4_ASAP7_75t_L g2682 ( 
.A(n_2140),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2140),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2464),
.B(n_2045),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2373),
.Y(n_2685)
);

AO22x2_ASAP7_75t_L g2686 ( 
.A1(n_2622),
.A2(n_2645),
.B1(n_2585),
.B2(n_2632),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2542),
.B(n_2182),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2373),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2375),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2375),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2384),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2384),
.Y(n_2692)
);

CKINVDCx20_ASAP7_75t_R g2693 ( 
.A(n_2393),
.Y(n_2693)
);

BUFx4_ASAP7_75t_L g2694 ( 
.A(n_2681),
.Y(n_2694)
);

AND2x6_ASAP7_75t_L g2695 ( 
.A(n_2627),
.B(n_1823),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2542),
.B(n_2196),
.Y(n_2696)
);

OAI221xp5_ASAP7_75t_L g2697 ( 
.A1(n_2618),
.A2(n_2052),
.B1(n_2107),
.B2(n_2030),
.C(n_2300),
.Y(n_2697)
);

BUFx4f_ASAP7_75t_L g2698 ( 
.A(n_2555),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2389),
.Y(n_2699)
);

CKINVDCx20_ASAP7_75t_R g2700 ( 
.A(n_2393),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2389),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2338),
.B(n_2227),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_SL g2703 ( 
.A(n_2352),
.B(n_2303),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2403),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2403),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2338),
.B(n_2227),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2407),
.Y(n_2707)
);

INVx3_ASAP7_75t_L g2708 ( 
.A(n_2364),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2364),
.Y(n_2709)
);

INVx5_ASAP7_75t_L g2710 ( 
.A(n_2396),
.Y(n_2710)
);

INVxp67_ASAP7_75t_L g2711 ( 
.A(n_2385),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2329),
.B(n_2222),
.C(n_2212),
.Y(n_2712)
);

HB1xp67_ASAP7_75t_L g2713 ( 
.A(n_2399),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2521),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2407),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2410),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2547),
.B(n_2243),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2370),
.B(n_2240),
.Y(n_2718)
);

NAND3xp33_ASAP7_75t_L g2719 ( 
.A(n_2504),
.B(n_2260),
.C(n_2248),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2410),
.Y(n_2720)
);

NOR2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2585),
.B(n_2240),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2416),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2417),
.B(n_2307),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2416),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2328),
.Y(n_2725)
);

INVxp67_ASAP7_75t_SL g2726 ( 
.A(n_2331),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2394),
.B(n_2395),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2442),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2442),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2452),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2452),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2390),
.B(n_1761),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2547),
.B(n_1833),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2463),
.Y(n_2734)
);

BUFx6f_ASAP7_75t_L g2735 ( 
.A(n_2328),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2352),
.B(n_1834),
.Y(n_2736)
);

AND2x6_ASAP7_75t_L g2737 ( 
.A(n_2627),
.B(n_1834),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2463),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2390),
.B(n_1761),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2467),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2467),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2344),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2355),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2550),
.B(n_1743),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2328),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2404),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2406),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2550),
.B(n_1743),
.Y(n_2748)
);

OR2x2_ASAP7_75t_L g2749 ( 
.A(n_2424),
.B(n_1846),
.Y(n_2749)
);

CKINVDCx20_ASAP7_75t_R g2750 ( 
.A(n_2521),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2472),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2556),
.B(n_1743),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2408),
.Y(n_2753)
);

INVx4_ASAP7_75t_L g2754 ( 
.A(n_2465),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2409),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2412),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2472),
.Y(n_2757)
);

INVxp67_ASAP7_75t_L g2758 ( 
.A(n_2337),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2413),
.B(n_1761),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2427),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2328),
.Y(n_2761)
);

HB1xp67_ASAP7_75t_L g2762 ( 
.A(n_2454),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2556),
.B(n_1747),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2429),
.B(n_1782),
.Y(n_2764)
);

AND2x4_ASAP7_75t_L g2765 ( 
.A(n_2390),
.B(n_1782),
.Y(n_2765)
);

INVxp67_ASAP7_75t_L g2766 ( 
.A(n_2433),
.Y(n_2766)
);

BUFx6f_ASAP7_75t_L g2767 ( 
.A(n_2333),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2477),
.Y(n_2768)
);

BUFx6f_ASAP7_75t_L g2769 ( 
.A(n_2333),
.Y(n_2769)
);

AO22x2_ASAP7_75t_L g2770 ( 
.A1(n_2622),
.A2(n_2645),
.B1(n_2585),
.B2(n_2632),
.Y(n_2770)
);

AOI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2633),
.A2(n_1796),
.B1(n_1747),
.B2(n_1893),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2471),
.B(n_2439),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2431),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2465),
.B(n_2468),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2471),
.B(n_697),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2446),
.Y(n_2776)
);

OAI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_2648),
.A2(n_2679),
.B1(n_2492),
.B2(n_2334),
.C(n_2593),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2453),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2445),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2462),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2553),
.B(n_1747),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2439),
.B(n_697),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2364),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2633),
.A2(n_1796),
.B1(n_1893),
.B2(n_1718),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2466),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2469),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2330),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2330),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2490),
.B(n_698),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2477),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2335),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2335),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2445),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2336),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2336),
.Y(n_2795)
);

OR2x2_ASAP7_75t_L g2796 ( 
.A(n_2638),
.B(n_1796),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2586),
.B(n_1718),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2485),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2342),
.B(n_1718),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2333),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2340),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2340),
.Y(n_2802)
);

INVx1_ASAP7_75t_SL g2803 ( 
.A(n_2440),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2333),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2341),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2465),
.B(n_1756),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_SL g2807 ( 
.A1(n_2374),
.A2(n_2652),
.B1(n_2597),
.B2(n_2682),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2480),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2341),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2386),
.Y(n_2810)
);

NAND2x1p5_ASAP7_75t_L g2811 ( 
.A(n_2465),
.B(n_1722),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2465),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2440),
.B(n_698),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2468),
.B(n_1756),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2624),
.A2(n_1722),
.B1(n_1893),
.B2(n_1756),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2359),
.B(n_1722),
.Y(n_2816)
);

INVx4_ASAP7_75t_SL g2817 ( 
.A(n_2633),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2357),
.B(n_1722),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2468),
.Y(n_2819)
);

OA22x2_ASAP7_75t_L g2820 ( 
.A1(n_2677),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_2820)
);

AO22x2_ASAP7_75t_L g2821 ( 
.A1(n_2622),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2480),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2468),
.Y(n_2823)
);

BUFx2_ASAP7_75t_L g2824 ( 
.A(n_2332),
.Y(n_2824)
);

NOR2xp67_ASAP7_75t_L g2825 ( 
.A(n_2443),
.B(n_1893),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2423),
.B(n_1893),
.Y(n_2826)
);

AND2x6_ASAP7_75t_L g2827 ( 
.A(n_2628),
.B(n_78),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2347),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2347),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2633),
.A2(n_1756),
.B1(n_170),
.B2(n_171),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2482),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2378),
.Y(n_2832)
);

AND2x2_ASAP7_75t_SL g2833 ( 
.A(n_2595),
.B(n_169),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2482),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2486),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2486),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2624),
.A2(n_1756),
.B1(n_81),
.B2(n_79),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2487),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2334),
.B(n_2363),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2487),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2363),
.B(n_170),
.Y(n_2841)
);

OR2x6_ASAP7_75t_L g2842 ( 
.A(n_2425),
.B(n_171),
.Y(n_2842)
);

AND2x4_ASAP7_75t_L g2843 ( 
.A(n_2468),
.B(n_172),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2633),
.A2(n_173),
.B1(n_174),
.B2(n_172),
.Y(n_2844)
);

BUFx10_ASAP7_75t_L g2845 ( 
.A(n_2475),
.Y(n_2845)
);

NAND2x1p5_ASAP7_75t_L g2846 ( 
.A(n_2430),
.B(n_2448),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2555),
.B(n_80),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2513),
.Y(n_2848)
);

OAI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2624),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2849)
);

INVx5_ASAP7_75t_L g2850 ( 
.A(n_2396),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2513),
.Y(n_2851)
);

AOI22x1_ASAP7_75t_L g2852 ( 
.A1(n_2664),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2516),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2516),
.Y(n_2854)
);

AOI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2633),
.A2(n_175),
.B1(n_176),
.B2(n_174),
.Y(n_2855)
);

INVx5_ASAP7_75t_L g2856 ( 
.A(n_2396),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2546),
.B(n_2563),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2383),
.B(n_2444),
.Y(n_2858)
);

INVxp67_ASAP7_75t_SL g2859 ( 
.A(n_2331),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2527),
.Y(n_2860)
);

AND2x6_ASAP7_75t_L g2861 ( 
.A(n_2628),
.B(n_82),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2595),
.B(n_175),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2383),
.B(n_2444),
.Y(n_2863)
);

INVx2_ASAP7_75t_SL g2864 ( 
.A(n_2479),
.Y(n_2864)
);

OR2x6_ASAP7_75t_L g2865 ( 
.A(n_2600),
.B(n_176),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2430),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2527),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_SL g2868 ( 
.A(n_2624),
.B(n_177),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2420),
.B(n_2555),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2485),
.Y(n_2870)
);

INVx5_ASAP7_75t_L g2871 ( 
.A(n_2396),
.Y(n_2871)
);

NOR2xp33_ASAP7_75t_L g2872 ( 
.A(n_2456),
.B(n_701),
.Y(n_2872)
);

INVx2_ASAP7_75t_SL g2873 ( 
.A(n_2479),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2574),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_2378),
.Y(n_2875)
);

AND2x6_ASAP7_75t_L g2876 ( 
.A(n_2560),
.B(n_84),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2537),
.Y(n_2877)
);

BUFx6f_ASAP7_75t_L g2878 ( 
.A(n_2455),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2537),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2538),
.Y(n_2880)
);

INVx1_ASAP7_75t_SL g2881 ( 
.A(n_2609),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2456),
.B(n_702),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2548),
.B(n_84),
.Y(n_2883)
);

BUFx6f_ASAP7_75t_L g2884 ( 
.A(n_2455),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2538),
.Y(n_2885)
);

INVx1_ASAP7_75t_SL g2886 ( 
.A(n_2332),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2496),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2539),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2539),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2386),
.Y(n_2890)
);

INVx4_ASAP7_75t_L g2891 ( 
.A(n_2430),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2574),
.Y(n_2892)
);

INVxp67_ASAP7_75t_L g2893 ( 
.A(n_2620),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2478),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2571),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_L g2896 ( 
.A1(n_2596),
.A2(n_179),
.B1(n_180),
.B2(n_178),
.Y(n_2896)
);

INVx4_ASAP7_75t_L g2897 ( 
.A(n_2448),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2349),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2497),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2349),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2448),
.Y(n_2901)
);

AND2x6_ASAP7_75t_L g2902 ( 
.A(n_2560),
.B(n_85),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2358),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2358),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2450),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2548),
.B(n_85),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2595),
.B(n_178),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2360),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2360),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2420),
.B(n_678),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2372),
.Y(n_2911)
);

HB1xp67_ASAP7_75t_L g2912 ( 
.A(n_2572),
.Y(n_2912)
);

NOR2x1p5_ASAP7_75t_L g2913 ( 
.A(n_2600),
.B(n_2604),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2372),
.Y(n_2914)
);

INVxp67_ASAP7_75t_SL g2915 ( 
.A(n_2331),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2483),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2610),
.A2(n_181),
.B1(n_182),
.B2(n_179),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2600),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2456),
.B(n_679),
.Y(n_2919)
);

NAND2xp33_ASAP7_75t_L g2920 ( 
.A(n_2449),
.B(n_86),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2455),
.Y(n_2921)
);

INVx4_ASAP7_75t_L g2922 ( 
.A(n_2455),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2495),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2505),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2519),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2548),
.B(n_86),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_L g2927 ( 
.A(n_2367),
.B(n_680),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2535),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_L g2929 ( 
.A(n_2520),
.Y(n_2929)
);

INVxp67_ASAP7_75t_L g2930 ( 
.A(n_2579),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2507),
.B(n_680),
.Y(n_2931)
);

AND2x6_ASAP7_75t_L g2932 ( 
.A(n_2568),
.B(n_86),
.Y(n_2932)
);

INVx8_ASAP7_75t_L g2933 ( 
.A(n_2396),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2378),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2386),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2511),
.B(n_682),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2367),
.B(n_682),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2391),
.Y(n_2938)
);

AND2x4_ASAP7_75t_L g2939 ( 
.A(n_2415),
.B(n_2418),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_2520),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2526),
.B(n_683),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2526),
.B(n_683),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2458),
.Y(n_2943)
);

NAND3x1_ASAP7_75t_L g2944 ( 
.A(n_2562),
.B(n_87),
.C(n_88),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2415),
.B(n_181),
.Y(n_2945)
);

AO22x2_ASAP7_75t_L g2946 ( 
.A1(n_2645),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2526),
.B(n_182),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2476),
.Y(n_2948)
);

BUFx3_ASAP7_75t_L g2949 ( 
.A(n_2497),
.Y(n_2949)
);

AND2x6_ASAP7_75t_L g2950 ( 
.A(n_2568),
.B(n_2494),
.Y(n_2950)
);

INVxp67_ASAP7_75t_L g2951 ( 
.A(n_2579),
.Y(n_2951)
);

NOR2xp33_ASAP7_75t_L g2952 ( 
.A(n_2367),
.B(n_689),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2520),
.Y(n_2953)
);

AND2x4_ASAP7_75t_L g2954 ( 
.A(n_2418),
.B(n_183),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_L g2955 ( 
.A(n_2459),
.B(n_691),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2380),
.B(n_184),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2531),
.B(n_2541),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2624),
.A2(n_186),
.B1(n_187),
.B2(n_185),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2531),
.B(n_702),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2380),
.B(n_2426),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2481),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2489),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2450),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2541),
.B(n_705),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2450),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2457),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2381),
.B(n_87),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2457),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_2549),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2457),
.Y(n_2970)
);

AND2x4_ASAP7_75t_L g2971 ( 
.A(n_2559),
.B(n_185),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2493),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2520),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2436),
.B(n_186),
.Y(n_2974)
);

INVx2_ASAP7_75t_SL g2975 ( 
.A(n_2496),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2500),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2510),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2380),
.B(n_187),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2514),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_2719),
.A2(n_2611),
.B1(n_2605),
.B2(n_2634),
.Y(n_2980)
);

A2O1A1Ixp33_ASAP7_75t_L g2981 ( 
.A1(n_2727),
.A2(n_2578),
.B(n_2584),
.C(n_2524),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2916),
.B(n_2551),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2688),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2689),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2758),
.B(n_2602),
.Y(n_2985)
);

BUFx3_ASAP7_75t_L g2986 ( 
.A(n_2798),
.Y(n_2986)
);

AOI22xp33_ASAP7_75t_L g2987 ( 
.A1(n_2719),
.A2(n_2634),
.B1(n_2671),
.B2(n_2669),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2803),
.B(n_2602),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2898),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2777),
.B(n_2644),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2923),
.B(n_2558),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2924),
.B(n_2558),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2925),
.B(n_2346),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2900),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2803),
.B(n_2602),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2928),
.B(n_2674),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_SL g2997 ( 
.A(n_2869),
.B(n_2602),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2903),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2904),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2684),
.B(n_2533),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2908),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2943),
.B(n_2673),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2909),
.Y(n_3003)
);

INVx3_ASAP7_75t_L g3004 ( 
.A(n_2754),
.Y(n_3004)
);

AOI22xp5_ASAP7_75t_L g3005 ( 
.A1(n_2955),
.A2(n_2351),
.B1(n_2398),
.B2(n_2545),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2911),
.Y(n_3006)
);

BUFx3_ASAP7_75t_L g3007 ( 
.A(n_2870),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2699),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2707),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2894),
.B(n_2678),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2914),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2812),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2711),
.B(n_2533),
.Y(n_3013)
);

A2O1A1Ixp33_ASAP7_75t_SL g3014 ( 
.A1(n_2872),
.A2(n_2544),
.B(n_2613),
.C(n_2670),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2772),
.B(n_2678),
.Y(n_3015)
);

NAND3xp33_ASAP7_75t_SL g3016 ( 
.A(n_2868),
.B(n_2855),
.C(n_2597),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2746),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2857),
.B(n_2687),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2687),
.B(n_2579),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2789),
.B(n_2594),
.Y(n_3020)
);

BUFx3_ASAP7_75t_L g3021 ( 
.A(n_2899),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2766),
.B(n_2762),
.Y(n_3022)
);

INVxp67_ASAP7_75t_L g3023 ( 
.A(n_2713),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2712),
.A2(n_2659),
.B1(n_2368),
.B2(n_2634),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2747),
.Y(n_3025)
);

A2O1A1Ixp33_ASAP7_75t_L g3026 ( 
.A1(n_2712),
.A2(n_2377),
.B(n_2534),
.C(n_2400),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2869),
.B(n_2602),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2696),
.B(n_2616),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2697),
.B(n_2437),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2696),
.B(n_2637),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2717),
.B(n_2666),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2717),
.B(n_2666),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2723),
.B(n_2666),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2779),
.B(n_2621),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2722),
.Y(n_3035)
);

INVx1_ASAP7_75t_SL g3036 ( 
.A(n_2886),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2728),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2730),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2881),
.B(n_2666),
.Y(n_3039)
);

CKINVDCx5p33_ASAP7_75t_R g3040 ( 
.A(n_2714),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2793),
.B(n_2621),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2881),
.B(n_2603),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2817),
.B(n_2603),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2817),
.B(n_2787),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2839),
.B(n_2398),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2788),
.B(n_2661),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2753),
.Y(n_3047)
);

O2A1O1Ixp5_ASAP7_75t_L g3048 ( 
.A1(n_2826),
.A2(n_2534),
.B(n_2434),
.C(n_2419),
.Y(n_3048)
);

BUFx12f_ASAP7_75t_L g3049 ( 
.A(n_2832),
.Y(n_3049)
);

CKINVDCx8_ASAP7_75t_R g3050 ( 
.A(n_2824),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2685),
.Y(n_3051)
);

AOI22xp33_ASAP7_75t_L g3052 ( 
.A1(n_2868),
.A2(n_2659),
.B1(n_2680),
.B2(n_2657),
.Y(n_3052)
);

NAND2x1p5_ASAP7_75t_L g3053 ( 
.A(n_2754),
.B(n_2380),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2749),
.B(n_2680),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2920),
.A2(n_2380),
.B(n_2356),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2791),
.B(n_2661),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2845),
.B(n_2604),
.Y(n_3057)
);

INVx2_ASAP7_75t_SL g3058 ( 
.A(n_2949),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2845),
.B(n_2604),
.Y(n_3059)
);

OR2x2_ASAP7_75t_L g3060 ( 
.A(n_2796),
.B(n_2557),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2792),
.B(n_2655),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2698),
.B(n_2621),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2755),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2941),
.A2(n_2540),
.B1(n_2569),
.B2(n_2509),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2756),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2794),
.B(n_2655),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2795),
.B(n_2572),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2718),
.B(n_2339),
.Y(n_3068)
);

NAND2x1p5_ASAP7_75t_L g3069 ( 
.A(n_2774),
.B(n_2326),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2690),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2812),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2782),
.B(n_2659),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2698),
.B(n_2607),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2774),
.B(n_2886),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2702),
.B(n_2683),
.Y(n_3075)
);

INVx2_ASAP7_75t_SL g3076 ( 
.A(n_2969),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2706),
.B(n_2339),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2760),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2930),
.B(n_2657),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2951),
.B(n_2657),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2912),
.B(n_2388),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2773),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2833),
.B(n_2683),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2776),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2957),
.B(n_2799),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2827),
.A2(n_2680),
.B1(n_2657),
.B2(n_2572),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2813),
.B(n_2557),
.Y(n_3087)
);

BUFx2_ASAP7_75t_L g3088 ( 
.A(n_2893),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2703),
.B(n_2680),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2939),
.B(n_2607),
.Y(n_3090)
);

AOI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2942),
.A2(n_2460),
.B1(n_2499),
.B2(n_2447),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2974),
.B(n_2656),
.Y(n_3092)
);

OR2x6_ASAP7_75t_L g3093 ( 
.A(n_2812),
.B(n_2549),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2693),
.B(n_2635),
.Y(n_3094)
);

OAI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2830),
.A2(n_2855),
.B1(n_2842),
.B2(n_2917),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2691),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2797),
.B(n_2656),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_2827),
.A2(n_2656),
.B1(n_2528),
.B2(n_2652),
.Y(n_3098)
);

AND2x6_ASAP7_75t_SL g3099 ( 
.A(n_2865),
.B(n_2599),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2847),
.B(n_2656),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2692),
.Y(n_3101)
);

OR2x2_ASAP7_75t_L g3102 ( 
.A(n_2759),
.B(n_2460),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2847),
.B(n_2656),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2967),
.B(n_2778),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2967),
.B(n_2780),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2913),
.B(n_2447),
.Y(n_3106)
);

O2A1O1Ixp5_ASAP7_75t_L g3107 ( 
.A1(n_2816),
.A2(n_2434),
.B(n_2419),
.C(n_2400),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2785),
.Y(n_3108)
);

BUFx6f_ASAP7_75t_L g3109 ( 
.A(n_2819),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2786),
.B(n_2939),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2971),
.B(n_2576),
.Y(n_3111)
);

AND2x4_ASAP7_75t_L g3112 ( 
.A(n_2913),
.B(n_2565),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2701),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2931),
.B(n_2649),
.Y(n_3114)
);

NAND2x1p5_ASAP7_75t_L g3115 ( 
.A(n_2819),
.B(n_2326),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2742),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2971),
.B(n_2576),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2743),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2704),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2895),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2818),
.A2(n_2356),
.B(n_2522),
.Y(n_3121)
);

OR2x2_ASAP7_75t_L g3122 ( 
.A(n_2874),
.B(n_2589),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2827),
.A2(n_2861),
.B1(n_2947),
.B2(n_2907),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2950),
.B(n_2632),
.Y(n_3124)
);

NAND2x1_ASAP7_75t_L g3125 ( 
.A(n_2708),
.B(n_2326),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_2827),
.A2(n_2528),
.B1(n_2652),
.B2(n_2591),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2705),
.Y(n_3127)
);

AOI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2700),
.A2(n_2374),
.B1(n_2451),
.B2(n_2543),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2801),
.B(n_2371),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2892),
.B(n_2614),
.Y(n_3130)
);

NOR3xp33_ASAP7_75t_L g3131 ( 
.A(n_2862),
.B(n_2580),
.C(n_2573),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2802),
.B(n_2371),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2715),
.Y(n_3133)
);

OAI22xp5_ASAP7_75t_L g3134 ( 
.A1(n_2830),
.A2(n_2946),
.B1(n_2821),
.B2(n_2844),
.Y(n_3134)
);

NOR3xp33_ASAP7_75t_L g3135 ( 
.A(n_2882),
.B(n_2573),
.C(n_2564),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2805),
.B(n_2387),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2919),
.A2(n_2646),
.B1(n_2512),
.B2(n_2619),
.Y(n_3137)
);

NOR2xp33_ASAP7_75t_L g3138 ( 
.A(n_2927),
.B(n_2614),
.Y(n_3138)
);

OR2x6_ASAP7_75t_L g3139 ( 
.A(n_2819),
.B(n_2590),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_2858),
.B(n_2590),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2716),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2720),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2861),
.A2(n_2528),
.B1(n_2652),
.B2(n_2676),
.Y(n_3143)
);

AOI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2937),
.A2(n_2619),
.B1(n_2528),
.B2(n_2658),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2936),
.B(n_2663),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2809),
.B(n_2387),
.Y(n_3146)
);

NOR3xp33_ASAP7_75t_L g3147 ( 
.A(n_2952),
.B(n_2582),
.C(n_2601),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_2861),
.A2(n_2528),
.B1(n_2676),
.B2(n_2654),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2724),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2828),
.B(n_2663),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2841),
.B(n_2663),
.Y(n_3151)
);

NAND3xp33_ASAP7_75t_L g3152 ( 
.A(n_2958),
.B(n_2392),
.C(n_2665),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2775),
.B(n_2647),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2829),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2729),
.B(n_2391),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2818),
.A2(n_2356),
.B(n_2522),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2823),
.B(n_2494),
.Y(n_3157)
);

OR2x6_ASAP7_75t_L g3158 ( 
.A(n_2823),
.B(n_2651),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2731),
.B(n_2391),
.Y(n_3159)
);

AO22x1_ASAP7_75t_L g3160 ( 
.A1(n_2861),
.A2(n_2682),
.B1(n_2588),
.B2(n_2606),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2734),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2823),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2738),
.B(n_2401),
.Y(n_3163)
);

OR2x2_ASAP7_75t_L g3164 ( 
.A(n_2979),
.B(n_2588),
.Y(n_3164)
);

AOI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_2821),
.A2(n_2528),
.B1(n_2654),
.B2(n_2643),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2740),
.B(n_2401),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_2858),
.B(n_2494),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2741),
.B(n_2401),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2950),
.B(n_2494),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2807),
.B(n_2682),
.Y(n_3170)
);

AOI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_2710),
.A2(n_2525),
.B(n_2508),
.Y(n_3171)
);

INVx4_ASAP7_75t_L g3172 ( 
.A(n_2878),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2950),
.A2(n_2441),
.B1(n_2654),
.B2(n_2643),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_2863),
.B(n_2536),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2950),
.B(n_2343),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2751),
.Y(n_3176)
);

NAND2xp33_ASAP7_75t_L g3177 ( 
.A(n_2929),
.B(n_2940),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2781),
.B(n_2664),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2757),
.Y(n_3179)
);

AOI22xp33_ASAP7_75t_L g3180 ( 
.A1(n_2946),
.A2(n_2676),
.B1(n_2643),
.B2(n_2650),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2768),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2790),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2863),
.B(n_2474),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2781),
.B(n_2350),
.Y(n_3184)
);

INVxp67_ASAP7_75t_L g3185 ( 
.A(n_2864),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2808),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_2708),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2849),
.A2(n_2650),
.B1(n_2647),
.B2(n_2672),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_SL g3189 ( 
.A(n_2843),
.B(n_2515),
.Y(n_3189)
);

NAND2x1_ASAP7_75t_L g3190 ( 
.A(n_2709),
.B(n_2354),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2744),
.B(n_2647),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_2918),
.Y(n_3192)
);

OAI21xp33_ASAP7_75t_L g3193 ( 
.A1(n_2896),
.A2(n_2606),
.B(n_2592),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2822),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2843),
.B(n_2554),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2834),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2744),
.B(n_2650),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_2807),
.B(n_2592),
.Y(n_3198)
);

O2A1O1Ixp33_ASAP7_75t_L g3199 ( 
.A1(n_2837),
.A2(n_2601),
.B(n_2625),
.C(n_2675),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2831),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2748),
.B(n_2361),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2929),
.B(n_2345),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2748),
.B(n_2362),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2725),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2948),
.B(n_2641),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3017),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3025),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3047),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_3064),
.B(n_2929),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_3140),
.B(n_2940),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3063),
.Y(n_3211)
);

INVx4_ASAP7_75t_L g3212 ( 
.A(n_3040),
.Y(n_3212)
);

INVxp67_ASAP7_75t_SL g3213 ( 
.A(n_3042),
.Y(n_3213)
);

AND2x4_ASAP7_75t_L g3214 ( 
.A(n_3140),
.B(n_2940),
.Y(n_3214)
);

AOI22xp5_ASAP7_75t_L g3215 ( 
.A1(n_3138),
.A2(n_2944),
.B1(n_2842),
.B2(n_2934),
.Y(n_3215)
);

INVx2_ASAP7_75t_SL g3216 ( 
.A(n_2986),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_3049),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_3112),
.B(n_2953),
.Y(n_3218)
);

INVx2_ASAP7_75t_SL g3219 ( 
.A(n_3007),
.Y(n_3219)
);

NOR2xp33_ASAP7_75t_L g3220 ( 
.A(n_3000),
.B(n_2842),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3065),
.Y(n_3221)
);

HB1xp67_ASAP7_75t_L g3222 ( 
.A(n_3042),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2983),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3018),
.B(n_2686),
.Y(n_3224)
);

A2O1A1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_3029),
.A2(n_2825),
.B(n_2917),
.C(n_2639),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_3050),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2984),
.Y(n_3227)
);

BUFx6f_ASAP7_75t_L g3228 ( 
.A(n_3204),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3078),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3082),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3084),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3204),
.Y(n_3232)
);

AOI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2990),
.A2(n_2875),
.B1(n_2750),
.B2(n_2721),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3020),
.B(n_2910),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_3034),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3008),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_3204),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2981),
.B(n_2686),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3108),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_3041),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3028),
.B(n_2770),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3009),
.Y(n_3242)
);

BUFx2_ASAP7_75t_L g3243 ( 
.A(n_3036),
.Y(n_3243)
);

HB1xp67_ASAP7_75t_L g3244 ( 
.A(n_3039),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3030),
.B(n_2770),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_3035),
.Y(n_3246)
);

AO22x1_ASAP7_75t_L g3247 ( 
.A1(n_3057),
.A2(n_2837),
.B1(n_2902),
.B2(n_2876),
.Y(n_3247)
);

INVx3_ASAP7_75t_L g3248 ( 
.A(n_3012),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3005),
.B(n_2953),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3031),
.B(n_2405),
.Y(n_3250)
);

INVx2_ASAP7_75t_SL g3251 ( 
.A(n_3021),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_3012),
.Y(n_3252)
);

OR2x2_ASAP7_75t_SL g3253 ( 
.A(n_3016),
.B(n_2694),
.Y(n_3253)
);

AND2x4_ASAP7_75t_L g3254 ( 
.A(n_3112),
.B(n_2953),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3032),
.B(n_2405),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_3060),
.Y(n_3256)
);

INVx2_ASAP7_75t_SL g3257 ( 
.A(n_3058),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3116),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3118),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_3033),
.B(n_2975),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_3012),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3164),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2996),
.B(n_2980),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3205),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3196),
.Y(n_3265)
);

BUFx3_ASAP7_75t_L g3266 ( 
.A(n_3076),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2989),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2994),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2998),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_3093),
.B(n_2973),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3091),
.A2(n_2721),
.B1(n_2956),
.B2(n_2978),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3037),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2999),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_3088),
.Y(n_3274)
);

INVx5_ASAP7_75t_L g3275 ( 
.A(n_3071),
.Y(n_3275)
);

BUFx12f_ASAP7_75t_L g3276 ( 
.A(n_3099),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3001),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_3102),
.B(n_2883),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_L g3279 ( 
.A(n_3081),
.B(n_2873),
.Y(n_3279)
);

CKINVDCx8_ASAP7_75t_R g3280 ( 
.A(n_3093),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3003),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3006),
.Y(n_3282)
);

BUFx2_ASAP7_75t_L g3283 ( 
.A(n_3192),
.Y(n_3283)
);

BUFx6f_ASAP7_75t_L g3284 ( 
.A(n_3071),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2996),
.B(n_2405),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3095),
.A2(n_2902),
.B1(n_2932),
.B2(n_2876),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3038),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3011),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3051),
.Y(n_3289)
);

BUFx2_ASAP7_75t_L g3290 ( 
.A(n_3023),
.Y(n_3290)
);

INVx4_ASAP7_75t_L g3291 ( 
.A(n_3093),
.Y(n_3291)
);

HB1xp67_ASAP7_75t_L g3292 ( 
.A(n_3120),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3104),
.B(n_2883),
.Y(n_3293)
);

INVxp67_ASAP7_75t_L g3294 ( 
.A(n_3022),
.Y(n_3294)
);

INVx2_ASAP7_75t_SL g3295 ( 
.A(n_3139),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3154),
.Y(n_3296)
);

BUFx3_ASAP7_75t_L g3297 ( 
.A(n_3139),
.Y(n_3297)
);

INVx4_ASAP7_75t_L g3298 ( 
.A(n_3139),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3070),
.Y(n_3299)
);

INVx3_ASAP7_75t_L g3300 ( 
.A(n_3071),
.Y(n_3300)
);

BUFx2_ASAP7_75t_L g3301 ( 
.A(n_3185),
.Y(n_3301)
);

INVx3_ASAP7_75t_L g3302 ( 
.A(n_3109),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_3109),
.Y(n_3303)
);

AND2x4_ASAP7_75t_L g3304 ( 
.A(n_3106),
.B(n_2973),
.Y(n_3304)
);

INVxp67_ASAP7_75t_L g3305 ( 
.A(n_3122),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3114),
.B(n_2959),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3105),
.B(n_2926),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2982),
.B(n_2973),
.Y(n_3308)
);

BUFx8_ASAP7_75t_L g3309 ( 
.A(n_3109),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3096),
.Y(n_3310)
);

BUFx2_ASAP7_75t_L g3311 ( 
.A(n_3075),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3013),
.B(n_2887),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3191),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3002),
.B(n_2982),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_3162),
.Y(n_3315)
);

AND2x4_ASAP7_75t_L g3316 ( 
.A(n_3106),
.B(n_2732),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_2987),
.A2(n_2865),
.B1(n_2825),
.B2(n_2876),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3046),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3046),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3056),
.Y(n_3320)
);

INVx5_ASAP7_75t_L g3321 ( 
.A(n_3162),
.Y(n_3321)
);

NOR2xp33_ASAP7_75t_SL g3322 ( 
.A(n_3134),
.B(n_2856),
.Y(n_3322)
);

AOI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_3152),
.A2(n_2865),
.B1(n_2902),
.B2(n_2876),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3056),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3083),
.B(n_2964),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3061),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3061),
.Y(n_3327)
);

NOR2xp67_ASAP7_75t_L g3328 ( 
.A(n_3059),
.B(n_2961),
.Y(n_3328)
);

INVx3_ASAP7_75t_L g3329 ( 
.A(n_3162),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3072),
.B(n_2945),
.Y(n_3330)
);

A2O1A1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_3026),
.A2(n_2639),
.B(n_2488),
.C(n_2675),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_3172),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3066),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3066),
.Y(n_3334)
);

CKINVDCx20_ASAP7_75t_R g3335 ( 
.A(n_3094),
.Y(n_3335)
);

NOR2xp33_ASAP7_75t_R g3336 ( 
.A(n_3177),
.B(n_2878),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3002),
.B(n_2906),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3010),
.B(n_2906),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_3069),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3087),
.B(n_2945),
.Y(n_3340)
);

INVx1_ASAP7_75t_SL g3341 ( 
.A(n_3110),
.Y(n_3341)
);

CKINVDCx20_ASAP7_75t_R g3342 ( 
.A(n_3128),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3101),
.Y(n_3343)
);

BUFx3_ASAP7_75t_L g3344 ( 
.A(n_3130),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_3137),
.B(n_2598),
.Y(n_3345)
);

INVx5_ASAP7_75t_L g3346 ( 
.A(n_3158),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3113),
.Y(n_3347)
);

INVx2_ASAP7_75t_SL g3348 ( 
.A(n_3090),
.Y(n_3348)
);

BUFx12f_ASAP7_75t_L g3349 ( 
.A(n_3172),
.Y(n_3349)
);

HB1xp67_ASAP7_75t_L g3350 ( 
.A(n_3191),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3119),
.Y(n_3351)
);

BUFx12f_ASAP7_75t_L g3352 ( 
.A(n_3069),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_3054),
.B(n_2962),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3010),
.B(n_2926),
.Y(n_3354)
);

BUFx3_ASAP7_75t_L g3355 ( 
.A(n_3115),
.Y(n_3355)
);

HB1xp67_ASAP7_75t_L g3356 ( 
.A(n_3197),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3127),
.Y(n_3357)
);

INVxp67_ASAP7_75t_SL g3358 ( 
.A(n_3197),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3133),
.Y(n_3359)
);

INVx2_ASAP7_75t_SL g3360 ( 
.A(n_3111),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3085),
.B(n_2612),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2993),
.B(n_2612),
.Y(n_3362)
);

BUFx6f_ASAP7_75t_L g3363 ( 
.A(n_3117),
.Y(n_3363)
);

INVx3_ASAP7_75t_L g3364 ( 
.A(n_3115),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3141),
.Y(n_3365)
);

INVx2_ASAP7_75t_SL g3366 ( 
.A(n_3074),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3142),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_2993),
.B(n_2972),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3149),
.Y(n_3369)
);

INVx5_ASAP7_75t_L g3370 ( 
.A(n_3158),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3024),
.B(n_2617),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3161),
.Y(n_3372)
);

INVx2_ASAP7_75t_SL g3373 ( 
.A(n_3073),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3024),
.B(n_2617),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3176),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3147),
.B(n_3045),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_2997),
.B(n_2732),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3068),
.B(n_2976),
.Y(n_3378)
);

INVx1_ASAP7_75t_SL g3379 ( 
.A(n_3145),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_3027),
.B(n_2739),
.Y(n_3380)
);

AO21x2_ASAP7_75t_L g3381 ( 
.A1(n_3171),
.A2(n_2525),
.B(n_2508),
.Y(n_3381)
);

OR2x2_ASAP7_75t_L g3382 ( 
.A(n_3015),
.B(n_2623),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3100),
.B(n_2623),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_3089),
.B(n_2977),
.Y(n_3384)
);

BUFx2_ASAP7_75t_L g3385 ( 
.A(n_3151),
.Y(n_3385)
);

INVx2_ASAP7_75t_SL g3386 ( 
.A(n_3044),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_3097),
.B(n_2710),
.Y(n_3387)
);

INVxp67_ASAP7_75t_SL g3388 ( 
.A(n_3150),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3179),
.Y(n_3389)
);

HB1xp67_ASAP7_75t_L g3390 ( 
.A(n_3175),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3103),
.B(n_2631),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3181),
.Y(n_3392)
);

BUFx3_ASAP7_75t_L g3393 ( 
.A(n_3169),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3153),
.B(n_2954),
.Y(n_3394)
);

INVxp67_ASAP7_75t_L g3395 ( 
.A(n_2991),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3182),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3186),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3194),
.Y(n_3398)
);

OR2x6_ASAP7_75t_L g3399 ( 
.A(n_3160),
.B(n_2933),
.Y(n_3399)
);

BUFx3_ASAP7_75t_L g3400 ( 
.A(n_3169),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3134),
.A2(n_2932),
.B1(n_2902),
.B2(n_2432),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3200),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3150),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3184),
.B(n_2631),
.Y(n_3404)
);

BUFx2_ASAP7_75t_L g3405 ( 
.A(n_3124),
.Y(n_3405)
);

BUFx4f_ASAP7_75t_L g3406 ( 
.A(n_3158),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3129),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_L g3408 ( 
.A1(n_3131),
.A2(n_2932),
.B1(n_2432),
.B2(n_2577),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3077),
.B(n_2954),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2991),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_3193),
.A2(n_2852),
.B1(n_2820),
.B2(n_2932),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3184),
.B(n_2641),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_3092),
.B(n_2710),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3129),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3132),
.Y(n_3415)
);

AND2x2_ASAP7_75t_L g3416 ( 
.A(n_3325),
.B(n_3198),
.Y(n_3416)
);

BUFx6f_ASAP7_75t_L g3417 ( 
.A(n_3228),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3289),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_3225),
.A2(n_3055),
.B(n_3195),
.Y(n_3419)
);

BUFx6f_ASAP7_75t_L g3420 ( 
.A(n_3228),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_3328),
.B(n_3314),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_3331),
.A2(n_2501),
.B(n_3121),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3314),
.B(n_3014),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3206),
.Y(n_3424)
);

INVx4_ASAP7_75t_L g3425 ( 
.A(n_3275),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3256),
.B(n_3052),
.Y(n_3426)
);

OAI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3376),
.A2(n_3135),
.B(n_3107),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_3279),
.B(n_3170),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_3406),
.A2(n_2501),
.B(n_3156),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3406),
.A2(n_3189),
.B(n_2428),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3256),
.B(n_3019),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_3376),
.B(n_3144),
.Y(n_3432)
);

NOR2xp33_ASAP7_75t_L g3433 ( 
.A(n_3344),
.B(n_3062),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3363),
.B(n_3123),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3330),
.B(n_3143),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3341),
.B(n_2992),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3341),
.B(n_2992),
.Y(n_3437)
);

BUFx6f_ASAP7_75t_L g3438 ( 
.A(n_3228),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_3393),
.B(n_2985),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3294),
.B(n_3079),
.Y(n_3440)
);

AO32x1_ASAP7_75t_L g3441 ( 
.A1(n_3318),
.A2(n_3324),
.A3(n_3326),
.B1(n_3320),
.B2(n_3319),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3299),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3207),
.Y(n_3443)
);

O2A1O1Ixp5_ASAP7_75t_L g3444 ( 
.A1(n_3249),
.A2(n_3048),
.B(n_3183),
.C(n_2428),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3294),
.B(n_3080),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3208),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3211),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3220),
.B(n_3043),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3274),
.B(n_3043),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3337),
.A2(n_2856),
.B(n_2850),
.Y(n_3450)
);

O2A1O1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_3345),
.A2(n_3199),
.B(n_2988),
.C(n_2995),
.Y(n_3451)
);

OAI22x1_ASAP7_75t_L g3452 ( 
.A1(n_3215),
.A2(n_3323),
.B1(n_3317),
.B2(n_3378),
.Y(n_3452)
);

AOI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_3337),
.A2(n_2856),
.B(n_2850),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3342),
.A2(n_3098),
.B1(n_3086),
.B2(n_3126),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3353),
.B(n_3180),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_SL g3456 ( 
.A(n_3363),
.B(n_3263),
.Y(n_3456)
);

O2A1O1Ixp33_ASAP7_75t_L g3457 ( 
.A1(n_3209),
.A2(n_3360),
.B(n_3263),
.C(n_3361),
.Y(n_3457)
);

OR2x2_ASAP7_75t_SL g3458 ( 
.A(n_3363),
.B(n_2642),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3293),
.A2(n_2871),
.B(n_2850),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3293),
.A2(n_2871),
.B(n_2435),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3307),
.A2(n_2871),
.B(n_2435),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3307),
.A2(n_2353),
.B(n_2327),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_3232),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3399),
.A2(n_2353),
.B(n_2327),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3286),
.A2(n_3165),
.B1(n_3188),
.B2(n_3148),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3244),
.B(n_2642),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3399),
.A2(n_2933),
.B(n_2815),
.Y(n_3467)
);

CKINVDCx5p33_ASAP7_75t_R g3468 ( 
.A(n_3226),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_SL g3469 ( 
.A1(n_3312),
.A2(n_3260),
.B(n_3411),
.C(n_3339),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3361),
.A2(n_3174),
.B(n_3167),
.C(n_3044),
.Y(n_3470)
);

AOI22xp5_ASAP7_75t_L g3471 ( 
.A1(n_3271),
.A2(n_3173),
.B1(n_2432),
.B2(n_3067),
.Y(n_3471)
);

BUFx3_ASAP7_75t_L g3472 ( 
.A(n_3266),
.Y(n_3472)
);

NAND3xp33_ASAP7_75t_L g3473 ( 
.A(n_3411),
.B(n_2577),
.C(n_2506),
.Y(n_3473)
);

AOI21x1_ASAP7_75t_L g3474 ( 
.A1(n_3247),
.A2(n_3178),
.B(n_3175),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_L g3475 ( 
.A1(n_3387),
.A2(n_3178),
.B(n_2411),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_3373),
.B(n_3067),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_3399),
.A2(n_2933),
.B(n_2815),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3244),
.B(n_3132),
.Y(n_3478)
);

OAI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3233),
.A2(n_2660),
.B1(n_2567),
.B2(n_2629),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3395),
.B(n_3136),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3338),
.A2(n_2960),
.B(n_2566),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3306),
.B(n_2577),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3234),
.B(n_2577),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3395),
.B(n_3136),
.Y(n_3484)
);

O2A1O1Ixp33_ASAP7_75t_L g3485 ( 
.A1(n_3413),
.A2(n_2630),
.B(n_3157),
.C(n_2667),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3310),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3343),
.Y(n_3487)
);

O2A1O1Ixp33_ASAP7_75t_SL g3488 ( 
.A1(n_3308),
.A2(n_2630),
.B(n_3125),
.C(n_3190),
.Y(n_3488)
);

NAND2x1p5_ASAP7_75t_L g3489 ( 
.A(n_3275),
.B(n_2709),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3407),
.B(n_3146),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3414),
.B(n_3146),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3338),
.A2(n_2566),
.B(n_2552),
.Y(n_3492)
);

INVx4_ASAP7_75t_L g3493 ( 
.A(n_3275),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3415),
.B(n_3201),
.Y(n_3494)
);

AOI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3322),
.A2(n_2561),
.B1(n_2765),
.B2(n_2739),
.Y(n_3495)
);

OAI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3368),
.A2(n_2608),
.B(n_2461),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3322),
.A2(n_2570),
.B1(n_2764),
.B2(n_2587),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3354),
.A2(n_2552),
.B(n_2461),
.Y(n_3498)
);

OAI22xp5_ASAP7_75t_L g3499 ( 
.A1(n_3401),
.A2(n_2615),
.B1(n_2771),
.B2(n_3201),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3366),
.B(n_3004),
.Y(n_3500)
);

AOI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3409),
.A2(n_2636),
.B1(n_2369),
.B2(n_2379),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_3348),
.A2(n_2441),
.B(n_2636),
.C(n_2529),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3354),
.A2(n_2366),
.B(n_2345),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3221),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_3410),
.B(n_3004),
.Y(n_3505)
);

OAI22x1_ASAP7_75t_L g3506 ( 
.A1(n_3305),
.A2(n_3202),
.B1(n_2771),
.B2(n_3187),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3311),
.B(n_3203),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3276),
.A2(n_2581),
.B1(n_2583),
.B2(n_2438),
.Y(n_3508)
);

INVxp67_ASAP7_75t_L g3509 ( 
.A(n_3243),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_3238),
.A2(n_2438),
.B1(n_2530),
.B2(n_2523),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_3358),
.A2(n_2366),
.B(n_2345),
.Y(n_3511)
);

OAI22xp5_ASAP7_75t_L g3512 ( 
.A1(n_3280),
.A2(n_3203),
.B1(n_2784),
.B2(n_2922),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_L g3513 ( 
.A(n_3235),
.B(n_2878),
.Y(n_3513)
);

BUFx12f_ASAP7_75t_L g3514 ( 
.A(n_3217),
.Y(n_3514)
);

O2A1O1Ixp33_ASAP7_75t_L g3515 ( 
.A1(n_3305),
.A2(n_3384),
.B(n_3362),
.C(n_3383),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3229),
.Y(n_3516)
);

INVx4_ASAP7_75t_L g3517 ( 
.A(n_3275),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3240),
.B(n_2884),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3358),
.A2(n_2376),
.B(n_2366),
.Y(n_3519)
);

OR2x6_ASAP7_75t_L g3520 ( 
.A(n_3238),
.B(n_3053),
.Y(n_3520)
);

NAND3xp33_ASAP7_75t_L g3521 ( 
.A(n_3408),
.B(n_2532),
.C(n_2470),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3213),
.B(n_3155),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3385),
.B(n_2905),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3230),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3213),
.B(n_3155),
.Y(n_3525)
);

NAND2x1p5_ASAP7_75t_L g3526 ( 
.A(n_3321),
.B(n_2783),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3278),
.B(n_2884),
.Y(n_3527)
);

NOR3xp33_ASAP7_75t_L g3528 ( 
.A(n_3291),
.B(n_2922),
.C(n_2736),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3365),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3369),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3388),
.A2(n_2376),
.B(n_2575),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3388),
.A2(n_2376),
.B(n_3053),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3335),
.A2(n_2765),
.B1(n_2449),
.B2(n_2396),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3223),
.Y(n_3534)
);

CKINVDCx5p33_ASAP7_75t_R g3535 ( 
.A(n_3212),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3379),
.B(n_3159),
.Y(n_3536)
);

AOI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3340),
.A2(n_2365),
.B1(n_2397),
.B2(n_2382),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3231),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_3297),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_L g3540 ( 
.A(n_3212),
.B(n_2884),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3301),
.B(n_2921),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3379),
.B(n_3159),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3346),
.B(n_2921),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3290),
.B(n_2921),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3346),
.A2(n_2859),
.B(n_2726),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3253),
.A2(n_2668),
.B1(n_3166),
.B2(n_3163),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3346),
.A2(n_2915),
.B(n_3163),
.Y(n_3547)
);

O2A1O1Ixp5_ASAP7_75t_L g3548 ( 
.A1(n_3285),
.A2(n_2653),
.B(n_3168),
.C(n_3166),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_3400),
.B(n_3187),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3264),
.B(n_3168),
.Y(n_3550)
);

A2O1A1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_3371),
.A2(n_2640),
.B(n_2662),
.C(n_2783),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3346),
.A2(n_2348),
.B(n_2354),
.Y(n_3552)
);

BUFx2_ASAP7_75t_L g3553 ( 
.A(n_3283),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3222),
.B(n_2835),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3222),
.B(n_2838),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3370),
.A2(n_2354),
.B(n_2421),
.Y(n_3556)
);

AOI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3285),
.A2(n_2626),
.B(n_2752),
.Y(n_3557)
);

OAI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3371),
.A2(n_2811),
.B1(n_2846),
.B2(n_2866),
.Y(n_3558)
);

O2A1O1Ixp33_ASAP7_75t_L g3559 ( 
.A1(n_3362),
.A2(n_2752),
.B(n_2763),
.C(n_2733),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3370),
.A2(n_3381),
.B(n_3224),
.Y(n_3560)
);

HB1xp67_ASAP7_75t_L g3561 ( 
.A(n_3292),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3262),
.B(n_2840),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3390),
.B(n_2851),
.Y(n_3563)
);

BUFx6f_ASAP7_75t_L g3564 ( 
.A(n_3232),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3239),
.Y(n_3565)
);

O2A1O1Ixp33_ASAP7_75t_L g3566 ( 
.A1(n_3383),
.A2(n_2763),
.B(n_2733),
.C(n_2853),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3258),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3259),
.Y(n_3568)
);

BUFx6f_ASAP7_75t_L g3569 ( 
.A(n_3232),
.Y(n_3569)
);

BUFx12f_ASAP7_75t_L g3570 ( 
.A(n_3349),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_SL g3571 ( 
.A1(n_3295),
.A2(n_3298),
.B1(n_3291),
.B2(n_3219),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_3216),
.B(n_2836),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3390),
.B(n_2854),
.Y(n_3573)
);

BUFx3_ASAP7_75t_L g3574 ( 
.A(n_3251),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3327),
.B(n_2877),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3333),
.B(n_2879),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_3270),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3265),
.Y(n_3578)
);

INVx2_ASAP7_75t_SL g3579 ( 
.A(n_3257),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3334),
.B(n_3391),
.Y(n_3580)
);

O2A1O1Ixp33_ASAP7_75t_L g3581 ( 
.A1(n_3391),
.A2(n_2880),
.B(n_2888),
.C(n_2885),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3316),
.B(n_2848),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3394),
.B(n_2860),
.Y(n_3583)
);

OAI22xp5_ASAP7_75t_SL g3584 ( 
.A1(n_3298),
.A2(n_2891),
.B1(n_2897),
.B2(n_2866),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_3370),
.B(n_2810),
.Y(n_3585)
);

BUFx6f_ASAP7_75t_L g3586 ( 
.A(n_3237),
.Y(n_3586)
);

OR2x6_ASAP7_75t_L g3587 ( 
.A(n_3224),
.B(n_2891),
.Y(n_3587)
);

NAND2xp33_ASAP7_75t_L g3588 ( 
.A(n_3336),
.B(n_2449),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3405),
.B(n_2867),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3313),
.B(n_2889),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3370),
.A2(n_2422),
.B(n_2421),
.Y(n_3591)
);

HB1xp67_ASAP7_75t_L g3592 ( 
.A(n_3292),
.Y(n_3592)
);

NAND2x1p5_ASAP7_75t_L g3593 ( 
.A(n_3321),
.B(n_2897),
.Y(n_3593)
);

AOI22xp33_ASAP7_75t_L g3594 ( 
.A1(n_3377),
.A2(n_2438),
.B1(n_2449),
.B2(n_2695),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3316),
.B(n_2810),
.Y(n_3595)
);

AOI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3377),
.A2(n_2449),
.B1(n_2438),
.B2(n_2695),
.Y(n_3596)
);

AO21x1_ASAP7_75t_L g3597 ( 
.A1(n_3374),
.A2(n_2503),
.B(n_2484),
.Y(n_3597)
);

AND2x4_ASAP7_75t_L g3598 ( 
.A(n_3304),
.B(n_2725),
.Y(n_3598)
);

INVx3_ASAP7_75t_L g3599 ( 
.A(n_3270),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3313),
.B(n_2963),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3267),
.Y(n_3601)
);

AND2x4_ASAP7_75t_SL g3602 ( 
.A(n_3210),
.B(n_2806),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3304),
.B(n_2965),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3350),
.B(n_3356),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3210),
.B(n_2890),
.Y(n_3605)
);

AOI33xp33_ASAP7_75t_L g3606 ( 
.A1(n_3268),
.A2(n_112),
.A3(n_96),
.B1(n_121),
.B2(n_104),
.B3(n_88),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3214),
.B(n_2890),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3350),
.B(n_2966),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_3214),
.B(n_2935),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3381),
.A2(n_2422),
.B(n_2421),
.Y(n_3610)
);

AO21x1_ASAP7_75t_L g3611 ( 
.A1(n_3374),
.A2(n_3245),
.B(n_3241),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3241),
.A2(n_2422),
.B(n_2411),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3245),
.A2(n_2411),
.B(n_2402),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3218),
.A2(n_2901),
.B1(n_2725),
.B2(n_2745),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3356),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3227),
.Y(n_3616)
);

HB1xp67_ASAP7_75t_L g3617 ( 
.A(n_3382),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_L g3618 ( 
.A(n_3386),
.B(n_2935),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3403),
.B(n_2968),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3404),
.B(n_2970),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3404),
.B(n_2938),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3218),
.B(n_3254),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3269),
.Y(n_3623)
);

INVx3_ASAP7_75t_L g3624 ( 
.A(n_3252),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3412),
.B(n_2938),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3419),
.A2(n_3255),
.B(n_3250),
.Y(n_3626)
);

OAI21x1_ASAP7_75t_L g3627 ( 
.A1(n_3422),
.A2(n_3255),
.B(n_3250),
.Y(n_3627)
);

AOI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_3588),
.A2(n_3412),
.B(n_3339),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3617),
.B(n_3273),
.Y(n_3629)
);

OAI21x1_ASAP7_75t_L g3630 ( 
.A1(n_3429),
.A2(n_2414),
.B(n_2402),
.Y(n_3630)
);

INVxp67_ASAP7_75t_SL g3631 ( 
.A(n_3561),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3610),
.A2(n_2414),
.B(n_2402),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3427),
.A2(n_3380),
.B(n_3351),
.Y(n_3633)
);

OAI21x1_ASAP7_75t_L g3634 ( 
.A1(n_3460),
.A2(n_2414),
.B(n_3277),
.Y(n_3634)
);

AO31x2_ASAP7_75t_L g3635 ( 
.A1(n_3597),
.A2(n_3282),
.A3(n_3288),
.B(n_3281),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3423),
.B(n_3296),
.Y(n_3636)
);

AO21x2_ASAP7_75t_L g3637 ( 
.A1(n_3461),
.A2(n_3357),
.B(n_3347),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3428),
.B(n_3254),
.Y(n_3638)
);

OAI21x1_ASAP7_75t_L g3639 ( 
.A1(n_3531),
.A2(n_3367),
.B(n_3359),
.Y(n_3639)
);

OAI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3471),
.A2(n_3380),
.B1(n_3355),
.B2(n_3332),
.Y(n_3640)
);

OAI22xp5_ASAP7_75t_L g3641 ( 
.A1(n_3508),
.A2(n_3352),
.B1(n_3364),
.B2(n_3372),
.Y(n_3641)
);

OAI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3455),
.A2(n_3364),
.B1(n_3321),
.B2(n_3389),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3467),
.A2(n_3397),
.B(n_3392),
.Y(n_3643)
);

OAI21x1_ASAP7_75t_L g3644 ( 
.A1(n_3477),
.A2(n_3402),
.B(n_3242),
.Y(n_3644)
);

INVx2_ASAP7_75t_SL g3645 ( 
.A(n_3472),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3424),
.Y(n_3646)
);

AOI21xp5_ASAP7_75t_SL g3647 ( 
.A1(n_3502),
.A2(n_2814),
.B(n_2806),
.Y(n_3647)
);

NAND2x1p5_ASAP7_75t_L g3648 ( 
.A(n_3425),
.B(n_3321),
.Y(n_3648)
);

AO22x2_ASAP7_75t_L g3649 ( 
.A1(n_3560),
.A2(n_3236),
.B1(n_3272),
.B2(n_3246),
.Y(n_3649)
);

OA21x2_ASAP7_75t_L g3650 ( 
.A1(n_3548),
.A2(n_3375),
.B(n_3287),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_3457),
.B(n_3396),
.Y(n_3651)
);

OAI21x1_ASAP7_75t_L g3652 ( 
.A1(n_3557),
.A2(n_3398),
.B(n_2502),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3612),
.A2(n_2473),
.B(n_2491),
.Y(n_3653)
);

O2A1O1Ixp5_ASAP7_75t_SL g3654 ( 
.A1(n_3456),
.A2(n_3300),
.B(n_3302),
.C(n_3248),
.Y(n_3654)
);

BUFx6f_ASAP7_75t_L g3655 ( 
.A(n_3417),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_SL g3656 ( 
.A(n_3432),
.B(n_3252),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3478),
.B(n_3248),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3552),
.A2(n_2518),
.B(n_2901),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3507),
.B(n_3300),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3443),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3448),
.B(n_3302),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3431),
.B(n_3440),
.Y(n_3662)
);

AND2x4_ASAP7_75t_L g3663 ( 
.A(n_3592),
.B(n_3303),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3445),
.B(n_3303),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_L g3665 ( 
.A1(n_3613),
.A2(n_2498),
.B(n_2491),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3436),
.B(n_3315),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3492),
.A2(n_2814),
.B(n_2503),
.Y(n_3667)
);

AOI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3506),
.A2(n_2438),
.B(n_3309),
.Y(n_3668)
);

AOI211x1_ASAP7_75t_L g3669 ( 
.A1(n_3611),
.A2(n_203),
.B(n_212),
.C(n_195),
.Y(n_3669)
);

BUFx6f_ASAP7_75t_L g3670 ( 
.A(n_3417),
.Y(n_3670)
);

OAI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3430),
.A2(n_2438),
.B(n_2449),
.Y(n_3671)
);

NAND2x1p5_ASAP7_75t_L g3672 ( 
.A(n_3425),
.B(n_3315),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3417),
.Y(n_3673)
);

OAI21x1_ASAP7_75t_L g3674 ( 
.A1(n_3532),
.A2(n_2498),
.B(n_2491),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3437),
.B(n_3329),
.Y(n_3675)
);

AOI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3474),
.A2(n_3309),
.B(n_2695),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3446),
.Y(n_3677)
);

INVx3_ASAP7_75t_L g3678 ( 
.A(n_3439),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3580),
.B(n_3329),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_3439),
.Y(n_3680)
);

OAI21x1_ASAP7_75t_L g3681 ( 
.A1(n_3475),
.A2(n_2517),
.B(n_2498),
.Y(n_3681)
);

CKINVDCx6p67_ASAP7_75t_R g3682 ( 
.A(n_3514),
.Y(n_3682)
);

NOR2xp67_ASAP7_75t_SL g3683 ( 
.A(n_3570),
.B(n_3252),
.Y(n_3683)
);

OAI21x1_ASAP7_75t_L g3684 ( 
.A1(n_3511),
.A2(n_2517),
.B(n_2695),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3421),
.B(n_3261),
.Y(n_3685)
);

NOR2xp67_ASAP7_75t_L g3686 ( 
.A(n_3447),
.B(n_3261),
.Y(n_3686)
);

O2A1O1Ixp5_ASAP7_75t_L g3687 ( 
.A1(n_3444),
.A2(n_2503),
.B(n_2484),
.C(n_2517),
.Y(n_3687)
);

OR2x6_ASAP7_75t_L g3688 ( 
.A(n_3571),
.B(n_3261),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3604),
.B(n_3284),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_SL g3690 ( 
.A1(n_3451),
.A2(n_2484),
.B(n_89),
.Y(n_3690)
);

OAI21x1_ASAP7_75t_SL g3691 ( 
.A1(n_3515),
.A2(n_89),
.B(n_90),
.Y(n_3691)
);

AOI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3434),
.A2(n_2737),
.B(n_3284),
.Y(n_3692)
);

OAI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3469),
.A2(n_2737),
.B(n_3284),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3416),
.B(n_3237),
.Y(n_3694)
);

AOI21xp5_ASAP7_75t_L g3695 ( 
.A1(n_3481),
.A2(n_2745),
.B(n_2735),
.Y(n_3695)
);

OA22x2_ASAP7_75t_L g3696 ( 
.A1(n_3452),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3480),
.B(n_3237),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3546),
.A2(n_2737),
.B(n_90),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3483),
.B(n_188),
.Y(n_3699)
);

OAI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3519),
.A2(n_2737),
.B(n_2735),
.Y(n_3700)
);

AOI221xp5_ASAP7_75t_L g3701 ( 
.A1(n_3479),
.A2(n_93),
.B1(n_95),
.B2(n_92),
.C(n_94),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3464),
.A2(n_2745),
.B(n_2735),
.Y(n_3702)
);

INVx1_ASAP7_75t_SL g3703 ( 
.A(n_3553),
.Y(n_3703)
);

NAND2x1p5_ASAP7_75t_L g3704 ( 
.A(n_3493),
.B(n_2761),
.Y(n_3704)
);

INVxp67_ASAP7_75t_L g3705 ( 
.A(n_3579),
.Y(n_3705)
);

AOI21xp33_ASAP7_75t_L g3706 ( 
.A1(n_3470),
.A2(n_2767),
.B(n_2761),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3473),
.A2(n_91),
.B(n_92),
.Y(n_3707)
);

CKINVDCx20_ASAP7_75t_R g3708 ( 
.A(n_3468),
.Y(n_3708)
);

AO21x2_ASAP7_75t_L g3709 ( 
.A1(n_3496),
.A2(n_2767),
.B(n_2761),
.Y(n_3709)
);

INVxp67_ASAP7_75t_SL g3710 ( 
.A(n_3615),
.Y(n_3710)
);

AOI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3543),
.A2(n_2769),
.B(n_2767),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3484),
.B(n_188),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3536),
.B(n_189),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3591),
.A2(n_2800),
.B(n_2769),
.Y(n_3714)
);

INVx4_ASAP7_75t_L g3715 ( 
.A(n_3493),
.Y(n_3715)
);

A2O1A1Ixp33_ASAP7_75t_L g3716 ( 
.A1(n_3606),
.A2(n_2804),
.B(n_2800),
.C(n_2769),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3450),
.A2(n_2804),
.B(n_2800),
.Y(n_3717)
);

BUFx2_ASAP7_75t_L g3718 ( 
.A(n_3458),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3495),
.A2(n_2804),
.B1(n_94),
.B2(n_91),
.Y(n_3719)
);

INVx4_ASAP7_75t_L g3720 ( 
.A(n_3517),
.Y(n_3720)
);

OAI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3485),
.A2(n_93),
.B(n_95),
.Y(n_3721)
);

AO21x2_ASAP7_75t_L g3722 ( 
.A1(n_3498),
.A2(n_93),
.B(n_95),
.Y(n_3722)
);

OAI21x1_ASAP7_75t_SL g3723 ( 
.A1(n_3581),
.A2(n_96),
.B(n_97),
.Y(n_3723)
);

OAI21x1_ASAP7_75t_L g3724 ( 
.A1(n_3453),
.A2(n_96),
.B(n_97),
.Y(n_3724)
);

OR2x2_ASAP7_75t_L g3725 ( 
.A(n_3504),
.B(n_190),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3542),
.B(n_192),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3482),
.B(n_192),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3494),
.B(n_193),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3503),
.A2(n_3566),
.B(n_3556),
.Y(n_3729)
);

INVx3_ASAP7_75t_L g3730 ( 
.A(n_3577),
.Y(n_3730)
);

OAI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3459),
.A2(n_97),
.B(n_98),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3426),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3732)
);

INVx3_ASAP7_75t_L g3733 ( 
.A(n_3577),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3547),
.A2(n_98),
.B(n_99),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3516),
.Y(n_3735)
);

OAI21x1_ASAP7_75t_SL g3736 ( 
.A1(n_3462),
.A2(n_99),
.B(n_101),
.Y(n_3736)
);

OAI22x1_ASAP7_75t_L g3737 ( 
.A1(n_3524),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3490),
.B(n_3491),
.Y(n_3738)
);

OAI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3433),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3739)
);

OAI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3512),
.A2(n_103),
.B(n_105),
.Y(n_3740)
);

INVx5_ASAP7_75t_L g3741 ( 
.A(n_3517),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3522),
.B(n_194),
.Y(n_3742)
);

INVx2_ASAP7_75t_SL g3743 ( 
.A(n_3574),
.Y(n_3743)
);

OR2x6_ASAP7_75t_L g3744 ( 
.A(n_3587),
.B(n_194),
.Y(n_3744)
);

NAND2x1_ASAP7_75t_L g3745 ( 
.A(n_3587),
.B(n_196),
.Y(n_3745)
);

INVx1_ASAP7_75t_SL g3746 ( 
.A(n_3527),
.Y(n_3746)
);

OAI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3501),
.A2(n_105),
.B(n_106),
.Y(n_3747)
);

CKINVDCx20_ASAP7_75t_R g3748 ( 
.A(n_3535),
.Y(n_3748)
);

NOR2xp33_ASAP7_75t_L g3749 ( 
.A(n_3449),
.B(n_197),
.Y(n_3749)
);

OAI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3501),
.A2(n_3521),
.B(n_3551),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3538),
.Y(n_3751)
);

OAI21x1_ASAP7_75t_L g3752 ( 
.A1(n_3559),
.A2(n_105),
.B(n_106),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3565),
.B(n_106),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_SL g3754 ( 
.A1(n_3466),
.A2(n_107),
.B(n_108),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3525),
.B(n_197),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3545),
.A2(n_107),
.B(n_108),
.Y(n_3756)
);

BUFx6f_ASAP7_75t_L g3757 ( 
.A(n_3420),
.Y(n_3757)
);

OAI21x1_ASAP7_75t_L g3758 ( 
.A1(n_3558),
.A2(n_107),
.B(n_108),
.Y(n_3758)
);

AO31x2_ASAP7_75t_L g3759 ( 
.A1(n_3499),
.A2(n_111),
.A3(n_109),
.B(n_110),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3509),
.B(n_198),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3567),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3568),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3621),
.A2(n_109),
.B(n_110),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3563),
.A2(n_109),
.B(n_111),
.Y(n_3764)
);

AO31x2_ASAP7_75t_L g3765 ( 
.A1(n_3578),
.A2(n_113),
.A3(n_111),
.B(n_112),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3465),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3585),
.A2(n_113),
.B(n_114),
.Y(n_3767)
);

BUFx6f_ASAP7_75t_L g3768 ( 
.A(n_3420),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3573),
.A2(n_116),
.B(n_117),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3550),
.B(n_198),
.Y(n_3770)
);

NOR2xp67_ASAP7_75t_L g3771 ( 
.A(n_3601),
.B(n_199),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3623),
.Y(n_3772)
);

OAI21x1_ASAP7_75t_L g3773 ( 
.A1(n_3625),
.A2(n_3620),
.B(n_3576),
.Y(n_3773)
);

A2O1A1Ixp33_ASAP7_75t_L g3774 ( 
.A1(n_3454),
.A2(n_201),
.B(n_202),
.C(n_200),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3505),
.A2(n_116),
.B(n_117),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3575),
.A2(n_117),
.B(n_118),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3441),
.Y(n_3777)
);

OA21x2_ASAP7_75t_L g3778 ( 
.A1(n_3510),
.A2(n_118),
.B(n_119),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3418),
.B(n_3442),
.Y(n_3779)
);

INVxp67_ASAP7_75t_L g3780 ( 
.A(n_3541),
.Y(n_3780)
);

OAI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_3476),
.A2(n_119),
.B(n_120),
.Y(n_3781)
);

BUFx3_ASAP7_75t_L g3782 ( 
.A(n_3539),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3486),
.B(n_203),
.Y(n_3783)
);

OAI21x1_ASAP7_75t_L g3784 ( 
.A1(n_3596),
.A2(n_120),
.B(n_121),
.Y(n_3784)
);

OAI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3497),
.A2(n_122),
.B(n_123),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3441),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3590),
.A2(n_122),
.B(n_123),
.Y(n_3787)
);

A2O1A1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3533),
.A2(n_206),
.B(n_207),
.C(n_205),
.Y(n_3788)
);

CKINVDCx20_ASAP7_75t_R g3789 ( 
.A(n_3622),
.Y(n_3789)
);

OAI21x1_ASAP7_75t_L g3790 ( 
.A1(n_3600),
.A2(n_122),
.B(n_124),
.Y(n_3790)
);

OAI21x1_ASAP7_75t_L g3791 ( 
.A1(n_3608),
.A2(n_124),
.B(n_126),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3537),
.A2(n_3500),
.B(n_3528),
.Y(n_3792)
);

BUFx3_ASAP7_75t_L g3793 ( 
.A(n_3420),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3487),
.B(n_207),
.Y(n_3794)
);

NAND3xp33_ASAP7_75t_L g3795 ( 
.A(n_3537),
.B(n_124),
.C(n_126),
.Y(n_3795)
);

BUFx4f_ASAP7_75t_L g3796 ( 
.A(n_3438),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3441),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3438),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3619),
.A2(n_126),
.B(n_127),
.Y(n_3799)
);

AO21x1_ASAP7_75t_L g3800 ( 
.A1(n_3618),
.A2(n_127),
.B(n_128),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3549),
.B(n_208),
.Y(n_3801)
);

O2A1O1Ixp5_ASAP7_75t_SL g3802 ( 
.A1(n_3599),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_3802)
);

AOI211x1_ASAP7_75t_L g3803 ( 
.A1(n_3583),
.A2(n_209),
.B(n_210),
.C(n_208),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3554),
.A2(n_128),
.B(n_129),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3488),
.A2(n_129),
.B(n_130),
.Y(n_3805)
);

OAI21x1_ASAP7_75t_SL g3806 ( 
.A1(n_3555),
.A2(n_130),
.B(n_131),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3594),
.A2(n_130),
.B(n_131),
.Y(n_3807)
);

INVx3_ASAP7_75t_L g3808 ( 
.A(n_3599),
.Y(n_3808)
);

AOI21xp5_ASAP7_75t_L g3809 ( 
.A1(n_3614),
.A2(n_131),
.B(n_132),
.Y(n_3809)
);

AO31x2_ASAP7_75t_L g3810 ( 
.A1(n_3529),
.A2(n_132),
.A3(n_211),
.B(n_210),
.Y(n_3810)
);

NAND2x1_ASAP7_75t_L g3811 ( 
.A(n_3587),
.B(n_211),
.Y(n_3811)
);

BUFx2_ASAP7_75t_L g3812 ( 
.A(n_3624),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3530),
.A2(n_132),
.B(n_212),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_3544),
.B(n_213),
.Y(n_3814)
);

OAI21x1_ASAP7_75t_L g3815 ( 
.A1(n_3534),
.A2(n_213),
.B(n_214),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3584),
.A2(n_215),
.B(n_216),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3589),
.B(n_216),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3616),
.B(n_217),
.Y(n_3818)
);

BUFx2_ASAP7_75t_L g3819 ( 
.A(n_3624),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3562),
.A2(n_217),
.B(n_218),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3523),
.B(n_219),
.Y(n_3821)
);

CKINVDCx20_ASAP7_75t_R g3822 ( 
.A(n_3540),
.Y(n_3822)
);

CKINVDCx5p33_ASAP7_75t_R g3823 ( 
.A(n_3438),
.Y(n_3823)
);

OR2x6_ASAP7_75t_L g3824 ( 
.A(n_3520),
.B(n_220),
.Y(n_3824)
);

OAI21x1_ASAP7_75t_L g3825 ( 
.A1(n_3489),
.A2(n_220),
.B(n_221),
.Y(n_3825)
);

AO32x2_ASAP7_75t_L g3826 ( 
.A1(n_3520),
.A2(n_224),
.A3(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_3826)
);

INVx4_ASAP7_75t_L g3827 ( 
.A(n_3463),
.Y(n_3827)
);

AO31x2_ASAP7_75t_L g3828 ( 
.A1(n_3595),
.A2(n_225),
.A3(n_222),
.B(n_224),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3435),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3520),
.Y(n_3830)
);

A2O1A1Ixp33_ASAP7_75t_L g3831 ( 
.A1(n_3582),
.A2(n_232),
.B(n_229),
.C(n_231),
.Y(n_3831)
);

OAI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3526),
.A2(n_233),
.B(n_235),
.Y(n_3832)
);

OAI21x1_ASAP7_75t_L g3833 ( 
.A1(n_3593),
.A2(n_233),
.B(n_236),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3513),
.A2(n_236),
.B(n_237),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3518),
.A2(n_237),
.B(n_238),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3572),
.B(n_238),
.Y(n_3836)
);

AOI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3602),
.A2(n_240),
.B(n_242),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3603),
.B(n_242),
.Y(n_3838)
);

INVx4_ASAP7_75t_L g3839 ( 
.A(n_3463),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3605),
.A2(n_243),
.B(n_244),
.Y(n_3840)
);

OAI21x1_ASAP7_75t_L g3841 ( 
.A1(n_3607),
.A2(n_243),
.B(n_244),
.Y(n_3841)
);

OA21x2_ASAP7_75t_L g3842 ( 
.A1(n_3609),
.A2(n_245),
.B(n_246),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3463),
.B(n_245),
.Y(n_3843)
);

OAI21x1_ASAP7_75t_L g3844 ( 
.A1(n_3564),
.A2(n_247),
.B(n_249),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3564),
.Y(n_3845)
);

OAI21x1_ASAP7_75t_L g3846 ( 
.A1(n_3564),
.A2(n_3586),
.B(n_3569),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3569),
.B(n_708),
.Y(n_3847)
);

AOI21x1_ASAP7_75t_L g3848 ( 
.A1(n_3598),
.A2(n_250),
.B(n_251),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3598),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3849)
);

BUFx2_ASAP7_75t_L g3850 ( 
.A(n_3569),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3586),
.A2(n_253),
.B(n_254),
.Y(n_3851)
);

INVx3_ASAP7_75t_L g3852 ( 
.A(n_3586),
.Y(n_3852)
);

OAI21x1_ASAP7_75t_L g3853 ( 
.A1(n_3729),
.A2(n_253),
.B(n_255),
.Y(n_3853)
);

NAND3xp33_ASAP7_75t_L g3854 ( 
.A(n_3701),
.B(n_255),
.C(n_256),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3646),
.Y(n_3855)
);

OAI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3774),
.A2(n_257),
.B(n_258),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3636),
.B(n_257),
.Y(n_3857)
);

BUFx2_ASAP7_75t_L g3858 ( 
.A(n_3678),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3647),
.A2(n_258),
.B(n_259),
.Y(n_3859)
);

NOR2x1_ASAP7_75t_L g3860 ( 
.A(n_3662),
.B(n_3782),
.Y(n_3860)
);

INVx3_ASAP7_75t_SL g3861 ( 
.A(n_3748),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3707),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_3862)
);

NAND2x1p5_ASAP7_75t_L g3863 ( 
.A(n_3741),
.B(n_260),
.Y(n_3863)
);

OAI22xp5_ASAP7_75t_L g3864 ( 
.A1(n_3766),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_3864)
);

OAI21x1_ASAP7_75t_L g3865 ( 
.A1(n_3652),
.A2(n_262),
.B(n_263),
.Y(n_3865)
);

AND2x4_ASAP7_75t_L g3866 ( 
.A(n_3830),
.B(n_264),
.Y(n_3866)
);

O2A1O1Ixp33_ASAP7_75t_L g3867 ( 
.A1(n_3831),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3750),
.A2(n_265),
.B(n_267),
.Y(n_3868)
);

A2O1A1Ixp33_ASAP7_75t_L g3869 ( 
.A1(n_3721),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_3869)
);

OAI21x1_ASAP7_75t_L g3870 ( 
.A1(n_3653),
.A2(n_268),
.B(n_269),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3698),
.A2(n_270),
.B(n_271),
.Y(n_3871)
);

NOR2xp33_ASAP7_75t_L g3872 ( 
.A(n_3822),
.B(n_3780),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3631),
.B(n_271),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3660),
.Y(n_3874)
);

OR2x2_ASAP7_75t_L g3875 ( 
.A(n_3710),
.B(n_272),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3667),
.A2(n_272),
.B(n_273),
.Y(n_3876)
);

INVx3_ASAP7_75t_L g3877 ( 
.A(n_3655),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3795),
.A2(n_273),
.B(n_274),
.Y(n_3878)
);

OAI21xp33_ASAP7_75t_L g3879 ( 
.A1(n_3766),
.A2(n_274),
.B(n_275),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_L g3880 ( 
.A(n_3789),
.B(n_275),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3629),
.B(n_276),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3795),
.A2(n_276),
.B(n_277),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3772),
.Y(n_3883)
);

A2O1A1Ixp33_ASAP7_75t_L g3884 ( 
.A1(n_3740),
.A2(n_280),
.B(n_277),
.C(n_279),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3805),
.A2(n_3671),
.B(n_3687),
.Y(n_3885)
);

CKINVDCx5p33_ASAP7_75t_R g3886 ( 
.A(n_3708),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3677),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3677),
.Y(n_3888)
);

CKINVDCx11_ASAP7_75t_R g3889 ( 
.A(n_3682),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3738),
.B(n_281),
.Y(n_3890)
);

OAI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3756),
.A2(n_281),
.B(n_282),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3659),
.B(n_3657),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3689),
.B(n_283),
.Y(n_3893)
);

NOR4xp25_ASAP7_75t_L g3894 ( 
.A(n_3747),
.B(n_286),
.C(n_284),
.D(n_285),
.Y(n_3894)
);

OAI21x1_ASAP7_75t_L g3895 ( 
.A1(n_3668),
.A2(n_287),
.B(n_288),
.Y(n_3895)
);

OAI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3676),
.A2(n_287),
.B(n_288),
.Y(n_3896)
);

OAI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3851),
.A2(n_289),
.B(n_291),
.Y(n_3897)
);

INVxp67_ASAP7_75t_L g3898 ( 
.A(n_3661),
.Y(n_3898)
);

O2A1O1Ixp33_ASAP7_75t_SL g3899 ( 
.A1(n_3788),
.A2(n_293),
.B(n_289),
.C(n_292),
.Y(n_3899)
);

OAI22x1_ASAP7_75t_L g3900 ( 
.A1(n_3718),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3696),
.A2(n_299),
.B1(n_294),
.B2(n_297),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3703),
.B(n_299),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3830),
.B(n_301),
.Y(n_3903)
);

OAI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3834),
.A2(n_301),
.B(n_302),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_3655),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3658),
.A2(n_302),
.B(n_303),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3651),
.A2(n_303),
.B(n_304),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_3663),
.Y(n_3908)
);

OAI22xp5_ASAP7_75t_L g3909 ( 
.A1(n_3829),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3909)
);

O2A1O1Ixp5_ASAP7_75t_L g3910 ( 
.A1(n_3800),
.A2(n_3732),
.B(n_3811),
.C(n_3745),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3773),
.B(n_305),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3785),
.A2(n_306),
.B(n_307),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3633),
.B(n_307),
.Y(n_3913)
);

AO31x2_ASAP7_75t_L g3914 ( 
.A1(n_3777),
.A2(n_310),
.A3(n_308),
.B(n_309),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3694),
.B(n_308),
.Y(n_3915)
);

AO31x2_ASAP7_75t_L g3916 ( 
.A1(n_3777),
.A2(n_311),
.A3(n_309),
.B(n_310),
.Y(n_3916)
);

OAI21x1_ASAP7_75t_L g3917 ( 
.A1(n_3634),
.A2(n_311),
.B(n_312),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3735),
.Y(n_3918)
);

BUFx3_ASAP7_75t_L g3919 ( 
.A(n_3645),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3666),
.B(n_312),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3675),
.B(n_313),
.Y(n_3921)
);

O2A1O1Ixp5_ASAP7_75t_L g3922 ( 
.A1(n_3781),
.A2(n_317),
.B(n_314),
.C(n_315),
.Y(n_3922)
);

OAI21x1_ASAP7_75t_L g3923 ( 
.A1(n_3681),
.A2(n_3684),
.B(n_3632),
.Y(n_3923)
);

BUFx8_ASAP7_75t_L g3924 ( 
.A(n_3847),
.Y(n_3924)
);

OAI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3829),
.A2(n_317),
.B1(n_314),
.B2(n_315),
.Y(n_3925)
);

OAI21x1_ASAP7_75t_L g3926 ( 
.A1(n_3630),
.A2(n_319),
.B(n_320),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3679),
.B(n_3697),
.Y(n_3927)
);

OR2x2_ASAP7_75t_L g3928 ( 
.A(n_3735),
.B(n_319),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3751),
.B(n_320),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3664),
.B(n_321),
.Y(n_3930)
);

OAI21x1_ASAP7_75t_L g3931 ( 
.A1(n_3702),
.A2(n_321),
.B(n_322),
.Y(n_3931)
);

INVx5_ASAP7_75t_L g3932 ( 
.A(n_3824),
.Y(n_3932)
);

BUFx3_ASAP7_75t_L g3933 ( 
.A(n_3743),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3751),
.Y(n_3934)
);

OAI21x1_ASAP7_75t_L g3935 ( 
.A1(n_3665),
.A2(n_322),
.B(n_323),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3761),
.B(n_324),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3749),
.B(n_324),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3761),
.Y(n_3938)
);

A2O1A1Ixp33_ASAP7_75t_L g3939 ( 
.A1(n_3816),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_3939)
);

OAI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3849),
.A2(n_329),
.B1(n_325),
.B2(n_328),
.Y(n_3940)
);

AO21x1_ASAP7_75t_L g3941 ( 
.A1(n_3656),
.A2(n_3685),
.B(n_3753),
.Y(n_3941)
);

OAI21x1_ASAP7_75t_L g3942 ( 
.A1(n_3700),
.A2(n_330),
.B(n_331),
.Y(n_3942)
);

OAI21x1_ASAP7_75t_L g3943 ( 
.A1(n_3654),
.A2(n_330),
.B(n_332),
.Y(n_3943)
);

AO31x2_ASAP7_75t_L g3944 ( 
.A1(n_3786),
.A2(n_335),
.A3(n_332),
.B(n_334),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3678),
.B(n_334),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3762),
.B(n_336),
.Y(n_3946)
);

OAI22x1_ASAP7_75t_L g3947 ( 
.A1(n_3849),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.Y(n_3947)
);

O2A1O1Ixp33_ASAP7_75t_L g3948 ( 
.A1(n_3691),
.A2(n_341),
.B(n_337),
.C(n_340),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3628),
.A2(n_341),
.B(n_342),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3762),
.Y(n_3950)
);

A2O1A1Ixp33_ASAP7_75t_L g3951 ( 
.A1(n_3809),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_3951)
);

A2O1A1Ixp33_ASAP7_75t_L g3952 ( 
.A1(n_3775),
.A2(n_3835),
.B(n_3767),
.C(n_3792),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3649),
.Y(n_3953)
);

OAI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_3744),
.A2(n_346),
.B1(n_343),
.B2(n_344),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3663),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3637),
.A2(n_3649),
.B(n_3695),
.Y(n_3956)
);

OAI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3734),
.A2(n_346),
.B(n_347),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3680),
.B(n_347),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3680),
.B(n_348),
.Y(n_3959)
);

OAI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3744),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3779),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3812),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3746),
.B(n_350),
.Y(n_3963)
);

AO31x2_ASAP7_75t_L g3964 ( 
.A1(n_3786),
.A2(n_354),
.A3(n_352),
.B(n_353),
.Y(n_3964)
);

A2O1A1Ixp33_ASAP7_75t_L g3965 ( 
.A1(n_3837),
.A2(n_3752),
.B(n_3784),
.C(n_3758),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_L g3966 ( 
.A(n_3638),
.B(n_352),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3635),
.Y(n_3967)
);

CKINVDCx20_ASAP7_75t_R g3968 ( 
.A(n_3823),
.Y(n_3968)
);

AOI22xp5_ASAP7_75t_L g3969 ( 
.A1(n_3640),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3635),
.Y(n_3970)
);

CKINVDCx20_ASAP7_75t_R g3971 ( 
.A(n_3793),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3746),
.B(n_3626),
.Y(n_3972)
);

NOR2xp67_ASAP7_75t_SL g3973 ( 
.A(n_3741),
.B(n_356),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3730),
.B(n_356),
.Y(n_3974)
);

AO31x2_ASAP7_75t_L g3975 ( 
.A1(n_3797),
.A2(n_359),
.A3(n_357),
.B(n_358),
.Y(n_3975)
);

AOI221x1_ASAP7_75t_L g3976 ( 
.A1(n_3737),
.A2(n_361),
.B1(n_357),
.B2(n_359),
.C(n_362),
.Y(n_3976)
);

OR2x2_ASAP7_75t_L g3977 ( 
.A(n_3627),
.B(n_363),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3819),
.Y(n_3978)
);

AOI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3637),
.A2(n_363),
.B(n_366),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3635),
.Y(n_3980)
);

AO31x2_ASAP7_75t_L g3981 ( 
.A1(n_3797),
.A2(n_368),
.A3(n_366),
.B(n_367),
.Y(n_3981)
);

O2A1O1Ixp33_ASAP7_75t_SL g3982 ( 
.A1(n_3801),
.A2(n_370),
.B(n_367),
.C(n_369),
.Y(n_3982)
);

OAI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3639),
.A2(n_369),
.B(n_370),
.Y(n_3983)
);

AOI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3717),
.A2(n_371),
.B(n_372),
.Y(n_3984)
);

A2O1A1Ixp33_ASAP7_75t_L g3985 ( 
.A1(n_3719),
.A2(n_374),
.B(n_371),
.C(n_372),
.Y(n_3985)
);

A2O1A1Ixp33_ASAP7_75t_L g3986 ( 
.A1(n_3771),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3730),
.B(n_3733),
.Y(n_3987)
);

NAND2x1_ASAP7_75t_L g3988 ( 
.A(n_3715),
.B(n_376),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3821),
.B(n_377),
.Y(n_3989)
);

AOI221x1_ASAP7_75t_L g3990 ( 
.A1(n_3806),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.C(n_381),
.Y(n_3990)
);

AO31x2_ASAP7_75t_L g3991 ( 
.A1(n_3642),
.A2(n_381),
.A3(n_379),
.B(n_380),
.Y(n_3991)
);

AOI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3722),
.A2(n_382),
.B(n_383),
.Y(n_3992)
);

CKINVDCx5p33_ASAP7_75t_R g3993 ( 
.A(n_3850),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3722),
.A2(n_382),
.B(n_384),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3733),
.B(n_384),
.Y(n_3995)
);

INVx4_ASAP7_75t_L g3996 ( 
.A(n_3688),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3845),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3693),
.A2(n_385),
.B(n_386),
.Y(n_3998)
);

A2O1A1Ixp33_ASAP7_75t_L g3999 ( 
.A1(n_3771),
.A2(n_3716),
.B(n_3814),
.C(n_3739),
.Y(n_3999)
);

AO31x2_ASAP7_75t_L g4000 ( 
.A1(n_3641),
.A2(n_388),
.A3(n_385),
.B(n_386),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_L g4001 ( 
.A(n_3705),
.B(n_388),
.Y(n_4001)
);

AOI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3824),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_4002)
);

BUFx6f_ASAP7_75t_L g4003 ( 
.A(n_3655),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3845),
.Y(n_4004)
);

OAI21x1_ASAP7_75t_L g4005 ( 
.A1(n_3674),
.A2(n_389),
.B(n_392),
.Y(n_4005)
);

OAI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3803),
.A2(n_396),
.B1(n_392),
.B2(n_394),
.Y(n_4006)
);

OAI21x1_ASAP7_75t_L g4007 ( 
.A1(n_3643),
.A2(n_394),
.B(n_396),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3650),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3650),
.Y(n_4009)
);

OA21x2_ASAP7_75t_L g4010 ( 
.A1(n_3731),
.A2(n_397),
.B(n_398),
.Y(n_4010)
);

OAI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3802),
.A2(n_398),
.B(n_399),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3706),
.A2(n_3778),
.B(n_3709),
.Y(n_4012)
);

OAI21x1_ASAP7_75t_L g4013 ( 
.A1(n_3692),
.A2(n_399),
.B(n_400),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3778),
.A2(n_401),
.B(n_402),
.Y(n_4014)
);

AO22x1_ASAP7_75t_L g4015 ( 
.A1(n_3753),
.A2(n_3741),
.B1(n_3712),
.B2(n_3726),
.Y(n_4015)
);

A2O1A1Ixp33_ASAP7_75t_L g4016 ( 
.A1(n_3820),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_4016)
);

INVxp67_ASAP7_75t_L g4017 ( 
.A(n_3760),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3690),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_4018)
);

BUFx6f_ASAP7_75t_L g4019 ( 
.A(n_3670),
.Y(n_4019)
);

AO31x2_ASAP7_75t_L g4020 ( 
.A1(n_3715),
.A2(n_406),
.A3(n_404),
.B(n_405),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3810),
.Y(n_4021)
);

BUFx6f_ASAP7_75t_L g4022 ( 
.A(n_3670),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3709),
.A2(n_406),
.B(n_407),
.Y(n_4023)
);

INVx5_ASAP7_75t_L g4024 ( 
.A(n_3688),
.Y(n_4024)
);

BUFx3_ASAP7_75t_L g4025 ( 
.A(n_3670),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3711),
.A2(n_407),
.B(n_408),
.Y(n_4026)
);

AOI31xp67_ASAP7_75t_L g4027 ( 
.A1(n_3742),
.A2(n_411),
.A3(n_408),
.B(n_409),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3644),
.A2(n_409),
.B(n_411),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_SL g4029 ( 
.A(n_3755),
.B(n_412),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3810),
.Y(n_4030)
);

OAI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3803),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_4031)
);

O2A1O1Ixp33_ASAP7_75t_SL g4032 ( 
.A1(n_3836),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_4032)
);

AND2x2_ASAP7_75t_SL g4033 ( 
.A(n_3842),
.B(n_417),
.Y(n_4033)
);

INVx3_ASAP7_75t_L g4034 ( 
.A(n_3997),
.Y(n_4034)
);

OAI21x1_ASAP7_75t_L g4035 ( 
.A1(n_3956),
.A2(n_3870),
.B(n_4012),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_4004),
.Y(n_4036)
);

OAI21x1_ASAP7_75t_L g4037 ( 
.A1(n_3865),
.A2(n_3724),
.B(n_3736),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3860),
.B(n_3686),
.Y(n_4038)
);

OAI21x1_ASAP7_75t_L g4039 ( 
.A1(n_4008),
.A2(n_3763),
.B(n_3787),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3961),
.B(n_3764),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3887),
.Y(n_4041)
);

INVx2_ASAP7_75t_SL g4042 ( 
.A(n_3919),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3918),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_SL g4044 ( 
.A1(n_3941),
.A2(n_3754),
.B(n_3848),
.Y(n_4044)
);

OAI21x1_ASAP7_75t_L g4045 ( 
.A1(n_4009),
.A2(n_3791),
.B(n_3790),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3885),
.A2(n_3804),
.B(n_3799),
.Y(n_4046)
);

OAI21x1_ASAP7_75t_L g4047 ( 
.A1(n_3967),
.A2(n_3776),
.B(n_3815),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3950),
.Y(n_4048)
);

INVx3_ASAP7_75t_L g4049 ( 
.A(n_3955),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3888),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3934),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3953),
.B(n_3764),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3938),
.Y(n_4053)
);

BUFx3_ASAP7_75t_L g4054 ( 
.A(n_3968),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3970),
.A2(n_3813),
.B(n_3714),
.Y(n_4055)
);

OAI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3980),
.A2(n_3853),
.B(n_3923),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3868),
.A2(n_3844),
.B(n_3841),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_L g4058 ( 
.A1(n_3879),
.A2(n_3723),
.B1(n_3769),
.B2(n_3842),
.Y(n_4058)
);

OAI21x1_ASAP7_75t_L g4059 ( 
.A1(n_4021),
.A2(n_3840),
.B(n_3648),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_4033),
.B(n_4024),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3855),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3874),
.Y(n_4062)
);

BUFx12f_ASAP7_75t_L g4063 ( 
.A(n_3889),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3908),
.B(n_3808),
.Y(n_4064)
);

AOI222xp33_ASAP7_75t_L g4065 ( 
.A1(n_3856),
.A2(n_3854),
.B1(n_3891),
.B2(n_3904),
.C1(n_3864),
.C2(n_3909),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3962),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3978),
.Y(n_4067)
);

OAI21x1_ASAP7_75t_SL g4068 ( 
.A1(n_3996),
.A2(n_3713),
.B(n_3770),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3925),
.A2(n_3940),
.B1(n_3871),
.B2(n_4006),
.Y(n_4069)
);

OAI21x1_ASAP7_75t_L g4070 ( 
.A1(n_4030),
.A2(n_3833),
.B(n_3832),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_SL g4071 ( 
.A1(n_3932),
.A2(n_3769),
.B1(n_3826),
.B2(n_3725),
.Y(n_4071)
);

OAI21x1_ASAP7_75t_L g4072 ( 
.A1(n_3979),
.A2(n_3825),
.B(n_3808),
.Y(n_4072)
);

OA21x2_ASAP7_75t_L g4073 ( 
.A1(n_3972),
.A2(n_3686),
.B(n_3846),
.Y(n_4073)
);

OR2x6_ASAP7_75t_L g4074 ( 
.A(n_3996),
.B(n_3720),
.Y(n_4074)
);

OAI21x1_ASAP7_75t_L g4075 ( 
.A1(n_4007),
.A2(n_3672),
.B(n_3704),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3883),
.Y(n_4076)
);

INVx4_ASAP7_75t_L g4077 ( 
.A(n_3932),
.Y(n_4077)
);

AO21x1_ASAP7_75t_L g4078 ( 
.A1(n_4031),
.A2(n_3826),
.B(n_3817),
.Y(n_4078)
);

BUFx2_ASAP7_75t_L g4079 ( 
.A(n_3858),
.Y(n_4079)
);

OAI21x1_ASAP7_75t_L g4080 ( 
.A1(n_3917),
.A2(n_3807),
.B(n_3794),
.Y(n_4080)
);

AOI22x1_ASAP7_75t_L g4081 ( 
.A1(n_3859),
.A2(n_3947),
.B1(n_3900),
.B2(n_3998),
.Y(n_4081)
);

OAI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3926),
.A2(n_3818),
.B(n_3783),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3927),
.Y(n_4083)
);

OR2x2_ASAP7_75t_L g4084 ( 
.A(n_3892),
.B(n_3699),
.Y(n_4084)
);

AO21x2_ASAP7_75t_L g4085 ( 
.A1(n_3992),
.A2(n_3728),
.B(n_3843),
.Y(n_4085)
);

INVxp67_ASAP7_75t_SL g4086 ( 
.A(n_3911),
.Y(n_4086)
);

AND2x4_ASAP7_75t_L g4087 ( 
.A(n_3987),
.B(n_3852),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_4025),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3993),
.B(n_3727),
.Y(n_4089)
);

OA21x2_ASAP7_75t_L g4090 ( 
.A1(n_3994),
.A2(n_3838),
.B(n_3826),
.Y(n_4090)
);

OAI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_3952),
.A2(n_3683),
.B(n_3796),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3914),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3977),
.Y(n_4093)
);

OAI21x1_ASAP7_75t_L g4094 ( 
.A1(n_3983),
.A2(n_3852),
.B(n_3810),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4017),
.B(n_3759),
.Y(n_4095)
);

OAI21x1_ASAP7_75t_L g4096 ( 
.A1(n_3935),
.A2(n_3765),
.B(n_3759),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_3898),
.B(n_4015),
.Y(n_4097)
);

OAI21x1_ASAP7_75t_L g4098 ( 
.A1(n_4005),
.A2(n_3765),
.B(n_3759),
.Y(n_4098)
);

OR2x6_ASAP7_75t_L g4099 ( 
.A(n_4014),
.B(n_3720),
.Y(n_4099)
);

INVxp67_ASAP7_75t_L g4100 ( 
.A(n_3963),
.Y(n_4100)
);

OAI21x1_ASAP7_75t_L g4101 ( 
.A1(n_4028),
.A2(n_3765),
.B(n_3828),
.Y(n_4101)
);

INVxp67_ASAP7_75t_L g4102 ( 
.A(n_3857),
.Y(n_4102)
);

AO21x2_ASAP7_75t_L g4103 ( 
.A1(n_4023),
.A2(n_3669),
.B(n_3828),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3933),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3877),
.Y(n_4105)
);

CKINVDCx20_ASAP7_75t_R g4106 ( 
.A(n_3861),
.Y(n_4106)
);

OAI21x1_ASAP7_75t_L g4107 ( 
.A1(n_3895),
.A2(n_3828),
.B(n_3669),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3931),
.A2(n_3839),
.B(n_3827),
.Y(n_4108)
);

AO31x2_ASAP7_75t_L g4109 ( 
.A1(n_3976),
.A2(n_3827),
.A3(n_3839),
.B(n_3796),
.Y(n_4109)
);

OR2x2_ASAP7_75t_L g4110 ( 
.A(n_3873),
.B(n_3673),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3914),
.Y(n_4111)
);

AOI22xp33_ASAP7_75t_L g4112 ( 
.A1(n_3912),
.A2(n_3757),
.B1(n_3768),
.B2(n_3673),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_3867),
.A2(n_3798),
.B(n_3757),
.C(n_3768),
.Y(n_4113)
);

OAI21xp33_ASAP7_75t_SL g4114 ( 
.A1(n_3894),
.A2(n_3757),
.B(n_3673),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3914),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3905),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3916),
.B(n_3944),
.Y(n_4117)
);

INVx1_ASAP7_75t_SL g4118 ( 
.A(n_3875),
.Y(n_4118)
);

HB1xp67_ASAP7_75t_L g4119 ( 
.A(n_3916),
.Y(n_4119)
);

BUFx3_ASAP7_75t_L g4120 ( 
.A(n_3971),
.Y(n_4120)
);

A2O1A1Ixp33_ASAP7_75t_L g4121 ( 
.A1(n_3878),
.A2(n_3798),
.B(n_3768),
.C(n_419),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3916),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3937),
.A2(n_3798),
.B1(n_419),
.B2(n_417),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3913),
.A2(n_418),
.B(n_420),
.Y(n_4124)
);

AO31x2_ASAP7_75t_L g4125 ( 
.A1(n_3990),
.A2(n_421),
.A3(n_418),
.B(n_420),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3944),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3942),
.A2(n_421),
.B(n_422),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3944),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_L g4129 ( 
.A1(n_3882),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4129)
);

NAND2x1p5_ASAP7_75t_L g4130 ( 
.A(n_4024),
.B(n_423),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_3896),
.A2(n_426),
.B(n_427),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3964),
.Y(n_4132)
);

CKINVDCx6p67_ASAP7_75t_R g4133 ( 
.A(n_3932),
.Y(n_4133)
);

AO31x2_ASAP7_75t_L g4134 ( 
.A1(n_3965),
.A2(n_428),
.A3(n_426),
.B(n_427),
.Y(n_4134)
);

NAND2x1p5_ASAP7_75t_L g4135 ( 
.A(n_4024),
.B(n_428),
.Y(n_4135)
);

AOI21x1_ASAP7_75t_L g4136 ( 
.A1(n_3929),
.A2(n_429),
.B(n_430),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3905),
.Y(n_4137)
);

OAI22xp33_ASAP7_75t_L g4138 ( 
.A1(n_3969),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_4138)
);

OAI21x1_ASAP7_75t_L g4139 ( 
.A1(n_3943),
.A2(n_432),
.B(n_433),
.Y(n_4139)
);

NAND2x1p5_ASAP7_75t_L g4140 ( 
.A(n_3973),
.B(n_433),
.Y(n_4140)
);

NAND2x1p5_ASAP7_75t_L g4141 ( 
.A(n_4010),
.B(n_3945),
.Y(n_4141)
);

OAI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_4002),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3964),
.B(n_3975),
.Y(n_4143)
);

OAI21x1_ASAP7_75t_L g4144 ( 
.A1(n_4026),
.A2(n_434),
.B(n_435),
.Y(n_4144)
);

OAI21x1_ASAP7_75t_L g4145 ( 
.A1(n_3876),
.A2(n_436),
.B(n_437),
.Y(n_4145)
);

CKINVDCx20_ASAP7_75t_R g4146 ( 
.A(n_3886),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3964),
.Y(n_4147)
);

BUFx2_ASAP7_75t_L g4148 ( 
.A(n_3905),
.Y(n_4148)
);

OAI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_3869),
.A2(n_3862),
.B1(n_3901),
.B2(n_3884),
.Y(n_4149)
);

OAI21x1_ASAP7_75t_L g4150 ( 
.A1(n_4013),
.A2(n_437),
.B(n_438),
.Y(n_4150)
);

AND2x4_ASAP7_75t_L g4151 ( 
.A(n_3945),
.B(n_439),
.Y(n_4151)
);

O2A1O1Ixp33_ASAP7_75t_L g4152 ( 
.A1(n_3939),
.A2(n_442),
.B(n_440),
.C(n_441),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3975),
.Y(n_4153)
);

OAI21x1_ASAP7_75t_L g4154 ( 
.A1(n_3949),
.A2(n_441),
.B(n_442),
.Y(n_4154)
);

AOI22xp33_ASAP7_75t_L g4155 ( 
.A1(n_3897),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_4155)
);

BUFx3_ASAP7_75t_L g4156 ( 
.A(n_3924),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4003),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4003),
.Y(n_4158)
);

OR2x6_ASAP7_75t_L g4159 ( 
.A(n_3863),
.B(n_445),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3975),
.B(n_446),
.Y(n_4160)
);

OAI21x1_ASAP7_75t_L g4161 ( 
.A1(n_3936),
.A2(n_446),
.B(n_447),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3981),
.B(n_447),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3954),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3981),
.B(n_448),
.Y(n_4164)
);

AND2x4_ASAP7_75t_L g4165 ( 
.A(n_3974),
.B(n_449),
.Y(n_4165)
);

HB1xp67_ASAP7_75t_L g4166 ( 
.A(n_3981),
.Y(n_4166)
);

BUFx2_ASAP7_75t_L g4167 ( 
.A(n_4003),
.Y(n_4167)
);

AOI21x1_ASAP7_75t_L g4168 ( 
.A1(n_3946),
.A2(n_450),
.B(n_451),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_3872),
.B(n_451),
.Y(n_4169)
);

OR2x6_ASAP7_75t_SL g4170 ( 
.A(n_3903),
.B(n_452),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3928),
.Y(n_4171)
);

O2A1O1Ixp33_ASAP7_75t_L g4172 ( 
.A1(n_3951),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_4172)
);

OAI21x1_ASAP7_75t_L g4173 ( 
.A1(n_3984),
.A2(n_453),
.B(n_454),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4020),
.Y(n_4174)
);

OAI21x1_ASAP7_75t_L g4175 ( 
.A1(n_3906),
.A2(n_455),
.B(n_456),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4020),
.Y(n_4176)
);

OAI21x1_ASAP7_75t_L g4177 ( 
.A1(n_3957),
.A2(n_458),
.B(n_459),
.Y(n_4177)
);

NAND2x1p5_ASAP7_75t_L g4178 ( 
.A(n_4010),
.B(n_458),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_3924),
.Y(n_4179)
);

OAI21x1_ASAP7_75t_L g4180 ( 
.A1(n_3910),
.A2(n_459),
.B(n_460),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4019),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3915),
.B(n_460),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_4019),
.Y(n_4183)
);

AOI21x1_ASAP7_75t_L g4184 ( 
.A1(n_4029),
.A2(n_461),
.B(n_462),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4041),
.Y(n_4185)
);

AO31x2_ASAP7_75t_L g4186 ( 
.A1(n_4117),
.A2(n_4143),
.A3(n_4078),
.B(n_4111),
.Y(n_4186)
);

OR2x6_ASAP7_75t_L g4187 ( 
.A(n_4077),
.B(n_3988),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4043),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4073),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4048),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_4141),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4086),
.B(n_4083),
.Y(n_4192)
);

BUFx4f_ASAP7_75t_L g4193 ( 
.A(n_4063),
.Y(n_4193)
);

OA21x2_ASAP7_75t_L g4194 ( 
.A1(n_4035),
.A2(n_3881),
.B(n_3920),
.Y(n_4194)
);

OAI21x1_ASAP7_75t_SL g4195 ( 
.A1(n_4077),
.A2(n_3921),
.B(n_3893),
.Y(n_4195)
);

OAI21x1_ASAP7_75t_L g4196 ( 
.A1(n_4056),
.A2(n_3907),
.B(n_3958),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_4152),
.A2(n_3899),
.B(n_4016),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4119),
.Y(n_4198)
);

CKINVDCx20_ASAP7_75t_R g4199 ( 
.A(n_4146),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4086),
.B(n_3930),
.Y(n_4200)
);

OA21x2_ASAP7_75t_L g4201 ( 
.A1(n_4117),
.A2(n_3890),
.B(n_4011),
.Y(n_4201)
);

OAI21x1_ASAP7_75t_L g4202 ( 
.A1(n_4039),
.A2(n_3959),
.B(n_3995),
.Y(n_4202)
);

AND2x4_ASAP7_75t_L g4203 ( 
.A(n_4074),
.B(n_3866),
.Y(n_4203)
);

OAI21x1_ASAP7_75t_L g4204 ( 
.A1(n_4045),
.A2(n_3989),
.B(n_3922),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4119),
.Y(n_4205)
);

AO31x2_ASAP7_75t_L g4206 ( 
.A1(n_4143),
.A2(n_3986),
.A3(n_3999),
.B(n_3960),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4073),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4093),
.B(n_4100),
.Y(n_4208)
);

OA21x2_ASAP7_75t_L g4209 ( 
.A1(n_4092),
.A2(n_4001),
.B(n_3902),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4100),
.B(n_3991),
.Y(n_4210)
);

OR2x2_ASAP7_75t_L g4211 ( 
.A(n_4052),
.B(n_3991),
.Y(n_4211)
);

BUFx3_ASAP7_75t_L g4212 ( 
.A(n_4106),
.Y(n_4212)
);

OAI21x1_ASAP7_75t_L g4213 ( 
.A1(n_4094),
.A2(n_3948),
.B(n_4018),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_4152),
.A2(n_4032),
.B(n_3982),
.Y(n_4214)
);

OAI21x1_ASAP7_75t_L g4215 ( 
.A1(n_4101),
.A2(n_3966),
.B(n_3880),
.Y(n_4215)
);

AO31x2_ASAP7_75t_L g4216 ( 
.A1(n_4115),
.A2(n_3985),
.A3(n_4027),
.B(n_4000),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_4172),
.A2(n_4113),
.B(n_4060),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_4172),
.A2(n_3974),
.B(n_3866),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4141),
.Y(n_4219)
);

AOI21x1_ASAP7_75t_L g4220 ( 
.A1(n_4060),
.A2(n_4020),
.B(n_4000),
.Y(n_4220)
);

BUFx3_ASAP7_75t_L g4221 ( 
.A(n_4106),
.Y(n_4221)
);

OAI21x1_ASAP7_75t_L g4222 ( 
.A1(n_4055),
.A2(n_3991),
.B(n_4000),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4166),
.Y(n_4223)
);

NAND2x1p5_ASAP7_75t_L g4224 ( 
.A(n_4079),
.B(n_4019),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4102),
.B(n_4022),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4166),
.Y(n_4226)
);

AO31x2_ASAP7_75t_L g4227 ( 
.A1(n_4122),
.A2(n_4022),
.A3(n_465),
.B(n_463),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_4113),
.A2(n_4022),
.B(n_463),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4102),
.B(n_4146),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4050),
.Y(n_4230)
);

AO21x2_ASAP7_75t_L g4231 ( 
.A1(n_4160),
.A2(n_464),
.B(n_465),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4133),
.Y(n_4232)
);

OA21x2_ASAP7_75t_L g4233 ( 
.A1(n_4126),
.A2(n_464),
.B(n_466),
.Y(n_4233)
);

NAND2x1p5_ASAP7_75t_L g4234 ( 
.A(n_4042),
.B(n_466),
.Y(n_4234)
);

AOI21xp5_ASAP7_75t_L g4235 ( 
.A1(n_4149),
.A2(n_467),
.B(n_468),
.Y(n_4235)
);

HB1xp67_ASAP7_75t_L g4236 ( 
.A(n_4052),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4087),
.B(n_467),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4149),
.A2(n_708),
.B(n_468),
.Y(n_4238)
);

OAI21x1_ASAP7_75t_L g4239 ( 
.A1(n_4096),
.A2(n_4098),
.B(n_4047),
.Y(n_4239)
);

INVxp67_ASAP7_75t_L g4240 ( 
.A(n_4170),
.Y(n_4240)
);

AO21x1_ASAP7_75t_L g4241 ( 
.A1(n_4160),
.A2(n_469),
.B(n_471),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4051),
.Y(n_4242)
);

AO31x2_ASAP7_75t_L g4243 ( 
.A1(n_4128),
.A2(n_474),
.A3(n_472),
.B(n_473),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_4040),
.Y(n_4244)
);

CKINVDCx20_ASAP7_75t_R g4245 ( 
.A(n_4054),
.Y(n_4245)
);

AO31x2_ASAP7_75t_L g4246 ( 
.A1(n_4132),
.A2(n_477),
.A3(n_474),
.B(n_475),
.Y(n_4246)
);

BUFx3_ASAP7_75t_L g4247 ( 
.A(n_4120),
.Y(n_4247)
);

INVx4_ASAP7_75t_SL g4248 ( 
.A(n_4156),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_4095),
.B(n_478),
.Y(n_4249)
);

AO31x2_ASAP7_75t_L g4250 ( 
.A1(n_4147),
.A2(n_480),
.A3(n_478),
.B(n_479),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4034),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_4034),
.Y(n_4252)
);

BUFx2_ASAP7_75t_L g4253 ( 
.A(n_4038),
.Y(n_4253)
);

HB1xp67_ASAP7_75t_L g4254 ( 
.A(n_4040),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4053),
.Y(n_4255)
);

CKINVDCx14_ASAP7_75t_R g4256 ( 
.A(n_4179),
.Y(n_4256)
);

OR2x6_ASAP7_75t_L g4257 ( 
.A(n_4074),
.B(n_480),
.Y(n_4257)
);

OAI21x1_ASAP7_75t_L g4258 ( 
.A1(n_4059),
.A2(n_483),
.B(n_484),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4153),
.Y(n_4259)
);

AO222x2_ASAP7_75t_L g4260 ( 
.A1(n_4169),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.C1(n_486),
.C2(n_487),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4179),
.B(n_485),
.Y(n_4261)
);

AO21x2_ASAP7_75t_L g4262 ( 
.A1(n_4162),
.A2(n_4164),
.B(n_4095),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4118),
.B(n_486),
.Y(n_4263)
);

OR2x2_ASAP7_75t_L g4264 ( 
.A(n_4097),
.B(n_489),
.Y(n_4264)
);

BUFx3_ASAP7_75t_L g4265 ( 
.A(n_4104),
.Y(n_4265)
);

BUFx2_ASAP7_75t_L g4266 ( 
.A(n_4038),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4118),
.B(n_4171),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4061),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4062),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4036),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4162),
.Y(n_4271)
);

HB1xp67_ASAP7_75t_L g4272 ( 
.A(n_4174),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4049),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4090),
.B(n_490),
.Y(n_4274)
);

INVxp33_ASAP7_75t_L g4275 ( 
.A(n_4089),
.Y(n_4275)
);

BUFx6f_ASAP7_75t_L g4276 ( 
.A(n_4130),
.Y(n_4276)
);

AOI22xp33_ASAP7_75t_L g4277 ( 
.A1(n_4065),
.A2(n_4081),
.B1(n_4069),
.B2(n_4155),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4090),
.B(n_490),
.Y(n_4278)
);

OAI21x1_ASAP7_75t_L g4279 ( 
.A1(n_4070),
.A2(n_491),
.B(n_492),
.Y(n_4279)
);

AND2x4_ASAP7_75t_L g4280 ( 
.A(n_4074),
.B(n_491),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4084),
.B(n_492),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_4065),
.A2(n_493),
.B(n_494),
.Y(n_4282)
);

AOI21x1_ASAP7_75t_L g4283 ( 
.A1(n_4164),
.A2(n_493),
.B(n_494),
.Y(n_4283)
);

OA21x2_ASAP7_75t_L g4284 ( 
.A1(n_4176),
.A2(n_496),
.B(n_497),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4049),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4085),
.B(n_496),
.Y(n_4286)
);

OAI21x1_ASAP7_75t_L g4287 ( 
.A1(n_4046),
.A2(n_497),
.B(n_498),
.Y(n_4287)
);

OA21x2_ASAP7_75t_L g4288 ( 
.A1(n_4108),
.A2(n_498),
.B(n_499),
.Y(n_4288)
);

AND2x4_ASAP7_75t_L g4289 ( 
.A(n_4087),
.B(n_499),
.Y(n_4289)
);

OAI21x1_ASAP7_75t_L g4290 ( 
.A1(n_4072),
.A2(n_500),
.B(n_501),
.Y(n_4290)
);

OA21x2_ASAP7_75t_L g4291 ( 
.A1(n_4044),
.A2(n_500),
.B(n_501),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4076),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4064),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4148),
.Y(n_4294)
);

NAND3xp33_ASAP7_75t_L g4295 ( 
.A(n_4071),
.B(n_502),
.C(n_503),
.Y(n_4295)
);

NOR2xp33_ASAP7_75t_R g4296 ( 
.A(n_4184),
.B(n_502),
.Y(n_4296)
);

NAND2x1p5_ASAP7_75t_L g4297 ( 
.A(n_4167),
.B(n_503),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4178),
.Y(n_4298)
);

INVx1_ASAP7_75t_SL g4299 ( 
.A(n_4110),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4116),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4178),
.Y(n_4301)
);

OAI21x1_ASAP7_75t_L g4302 ( 
.A1(n_4082),
.A2(n_504),
.B(n_505),
.Y(n_4302)
);

AO31x2_ASAP7_75t_L g4303 ( 
.A1(n_4137),
.A2(n_504),
.A3(n_507),
.B(n_508),
.Y(n_4303)
);

HB1xp67_ASAP7_75t_L g4304 ( 
.A(n_4066),
.Y(n_4304)
);

CKINVDCx5p33_ASAP7_75t_R g4305 ( 
.A(n_4157),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4067),
.Y(n_4306)
);

NOR2x1_ASAP7_75t_R g4307 ( 
.A(n_4151),
.B(n_507),
.Y(n_4307)
);

AOI21x1_ASAP7_75t_L g4308 ( 
.A1(n_4068),
.A2(n_508),
.B(n_509),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4134),
.Y(n_4309)
);

AOI211xp5_ASAP7_75t_L g4310 ( 
.A1(n_4142),
.A2(n_509),
.B(n_510),
.C(n_511),
.Y(n_4310)
);

OAI21x1_ASAP7_75t_L g4311 ( 
.A1(n_4107),
.A2(n_510),
.B(n_512),
.Y(n_4311)
);

OAI21x1_ASAP7_75t_L g4312 ( 
.A1(n_4080),
.A2(n_512),
.B(n_513),
.Y(n_4312)
);

BUFx2_ASAP7_75t_L g4313 ( 
.A(n_4099),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4158),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4134),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_4105),
.B(n_694),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4134),
.Y(n_4317)
);

OAI21x1_ASAP7_75t_L g4318 ( 
.A1(n_4075),
.A2(n_514),
.B(n_515),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4181),
.Y(n_4319)
);

AND2x4_ASAP7_75t_L g4320 ( 
.A(n_4183),
.B(n_514),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_4091),
.A2(n_516),
.B(n_517),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4088),
.Y(n_4322)
);

OAI21x1_ASAP7_75t_L g4323 ( 
.A1(n_4057),
.A2(n_517),
.B(n_518),
.Y(n_4323)
);

BUFx3_ASAP7_75t_L g4324 ( 
.A(n_4165),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_4091),
.A2(n_518),
.B(n_519),
.Y(n_4325)
);

HB1xp67_ASAP7_75t_L g4326 ( 
.A(n_4085),
.Y(n_4326)
);

OA21x2_ASAP7_75t_L g4327 ( 
.A1(n_4057),
.A2(n_519),
.B(n_520),
.Y(n_4327)
);

AO31x2_ASAP7_75t_L g4328 ( 
.A1(n_4121),
.A2(n_521),
.A3(n_522),
.B(n_523),
.Y(n_4328)
);

INVx1_ASAP7_75t_SL g4329 ( 
.A(n_4182),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4071),
.B(n_521),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_4232),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4185),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4185),
.Y(n_4333)
);

AOI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4277),
.A2(n_4155),
.B1(n_4103),
.B2(n_4138),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_L g4335 ( 
.A1(n_4295),
.A2(n_4103),
.B1(n_4138),
.B2(n_4142),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4294),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_SL g4337 ( 
.A1(n_4217),
.A2(n_4135),
.B1(n_4130),
.B2(n_4140),
.Y(n_4337)
);

OAI22xp5_ASAP7_75t_L g4338 ( 
.A1(n_4240),
.A2(n_4058),
.B1(n_4121),
.B2(n_4123),
.Y(n_4338)
);

BUFx12f_ASAP7_75t_L g4339 ( 
.A(n_4234),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_4193),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4188),
.Y(n_4341)
);

NAND3xp33_ASAP7_75t_L g4342 ( 
.A(n_4282),
.B(n_4129),
.C(n_4124),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4188),
.Y(n_4343)
);

OAI22xp33_ASAP7_75t_L g4344 ( 
.A1(n_4330),
.A2(n_4099),
.B1(n_4159),
.B2(n_4135),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4197),
.A2(n_4058),
.B1(n_4112),
.B2(n_4129),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4190),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4276),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4203),
.B(n_4099),
.Y(n_4348)
);

OAI22xp5_ASAP7_75t_L g4349 ( 
.A1(n_4310),
.A2(n_4274),
.B1(n_4278),
.B2(n_4321),
.Y(n_4349)
);

INVx2_ASAP7_75t_SL g4350 ( 
.A(n_4193),
.Y(n_4350)
);

OAI21xp5_ASAP7_75t_SL g4351 ( 
.A1(n_4325),
.A2(n_4123),
.B(n_4124),
.Y(n_4351)
);

HB1xp67_ASAP7_75t_L g4352 ( 
.A(n_4288),
.Y(n_4352)
);

AOI22xp5_ASAP7_75t_L g4353 ( 
.A1(n_4241),
.A2(n_4114),
.B1(n_4112),
.B2(n_4163),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4286),
.A2(n_4163),
.B1(n_4140),
.B2(n_4159),
.Y(n_4354)
);

OAI22xp33_ASAP7_75t_L g4355 ( 
.A1(n_4276),
.A2(n_4159),
.B1(n_4168),
.B2(n_4136),
.Y(n_4355)
);

AOI22xp33_ASAP7_75t_L g4356 ( 
.A1(n_4201),
.A2(n_4238),
.B1(n_4235),
.B2(n_4327),
.Y(n_4356)
);

AOI22xp33_ASAP7_75t_L g4357 ( 
.A1(n_4201),
.A2(n_4177),
.B1(n_4154),
.B2(n_4175),
.Y(n_4357)
);

BUFx3_ASAP7_75t_L g4358 ( 
.A(n_4212),
.Y(n_4358)
);

BUFx12f_ASAP7_75t_L g4359 ( 
.A(n_4257),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4276),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4190),
.Y(n_4361)
);

AOI211xp5_ASAP7_75t_L g4362 ( 
.A1(n_4260),
.A2(n_4180),
.B(n_4173),
.C(n_4145),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4259),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4259),
.Y(n_4364)
);

AOI22xp33_ASAP7_75t_SL g4365 ( 
.A1(n_4327),
.A2(n_4151),
.B1(n_4161),
.B2(n_4165),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_4291),
.A2(n_4037),
.B1(n_4139),
.B2(n_4127),
.Y(n_4366)
);

AOI22xp33_ASAP7_75t_SL g4367 ( 
.A1(n_4215),
.A2(n_4131),
.B1(n_4144),
.B2(n_4150),
.Y(n_4367)
);

AOI22xp33_ASAP7_75t_SL g4368 ( 
.A1(n_4296),
.A2(n_4213),
.B1(n_4291),
.B2(n_4209),
.Y(n_4368)
);

AOI21xp33_ASAP7_75t_L g4369 ( 
.A1(n_4194),
.A2(n_4109),
.B(n_4125),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4198),
.Y(n_4370)
);

INVx3_ASAP7_75t_L g4371 ( 
.A(n_4232),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_L g4372 ( 
.A1(n_4262),
.A2(n_4125),
.B1(n_4109),
.B2(n_525),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4262),
.A2(n_4125),
.B1(n_4109),
.B2(n_526),
.Y(n_4373)
);

OAI22xp33_ASAP7_75t_L g4374 ( 
.A1(n_4257),
.A2(n_523),
.B1(n_524),
.B2(n_526),
.Y(n_4374)
);

BUFx12f_ASAP7_75t_L g4375 ( 
.A(n_4264),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_4313),
.A2(n_524),
.B1(n_527),
.B2(n_528),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_SL g4377 ( 
.A1(n_4209),
.A2(n_690),
.B1(n_530),
.B2(n_531),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4300),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4271),
.A2(n_529),
.B1(n_531),
.B2(n_532),
.Y(n_4379)
);

AOI22xp33_ASAP7_75t_SL g4380 ( 
.A1(n_4200),
.A2(n_529),
.B1(n_532),
.B2(n_533),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4198),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_SL g4382 ( 
.A1(n_4231),
.A2(n_687),
.B1(n_535),
.B2(n_536),
.Y(n_4382)
);

AOI22xp33_ASAP7_75t_L g4383 ( 
.A1(n_4271),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4205),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4205),
.Y(n_4385)
);

OAI21xp33_ASAP7_75t_L g4386 ( 
.A1(n_4214),
.A2(n_4210),
.B(n_4220),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4194),
.A2(n_537),
.B1(n_538),
.B2(n_540),
.Y(n_4387)
);

BUFx6f_ASAP7_75t_L g4388 ( 
.A(n_4280),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_SL g4389 ( 
.A1(n_4231),
.A2(n_685),
.B1(n_538),
.B2(n_540),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4298),
.B(n_537),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4203),
.B(n_541),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4298),
.B(n_4301),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_L g4393 ( 
.A1(n_4299),
.A2(n_541),
.B1(n_542),
.B2(n_543),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4223),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4314),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_4319),
.Y(n_4396)
);

BUFx6f_ASAP7_75t_L g4397 ( 
.A(n_4280),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_SL g4398 ( 
.A(n_4192),
.B(n_4229),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4293),
.B(n_543),
.Y(n_4399)
);

OAI21xp5_ASAP7_75t_SL g4400 ( 
.A1(n_4228),
.A2(n_544),
.B(n_545),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4223),
.Y(n_4401)
);

INVx3_ASAP7_75t_L g4402 ( 
.A(n_4224),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4301),
.B(n_544),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_4195),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_4404)
);

INVx4_ASAP7_75t_L g4405 ( 
.A(n_4248),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4208),
.B(n_546),
.Y(n_4406)
);

INVx8_ASAP7_75t_L g4407 ( 
.A(n_4320),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4226),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4218),
.A2(n_547),
.B1(n_548),
.B2(n_549),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4226),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4275),
.A2(n_4315),
.B1(n_4317),
.B2(n_4309),
.Y(n_4411)
);

INVx2_ASAP7_75t_SL g4412 ( 
.A(n_4248),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4268),
.Y(n_4413)
);

CKINVDCx5p33_ASAP7_75t_R g4414 ( 
.A(n_4199),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4309),
.A2(n_549),
.B1(n_550),
.B2(n_551),
.Y(n_4415)
);

OAI21xp5_ASAP7_75t_SL g4416 ( 
.A1(n_4261),
.A2(n_550),
.B(n_551),
.Y(n_4416)
);

OAI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4233),
.A2(n_552),
.B1(n_553),
.B2(n_554),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4273),
.Y(n_4418)
);

OAI22xp5_ASAP7_75t_L g4419 ( 
.A1(n_4249),
.A2(n_552),
.B1(n_554),
.B2(n_555),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4253),
.B(n_555),
.Y(n_4420)
);

AOI22xp5_ASAP7_75t_L g4421 ( 
.A1(n_4187),
.A2(n_556),
.B1(n_557),
.B2(n_558),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4315),
.A2(n_556),
.B1(n_558),
.B2(n_559),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4285),
.Y(n_4423)
);

AOI22xp33_ASAP7_75t_SL g4424 ( 
.A1(n_4288),
.A2(n_681),
.B1(n_560),
.B2(n_561),
.Y(n_4424)
);

OAI22xp5_ASAP7_75t_L g4425 ( 
.A1(n_4187),
.A2(n_559),
.B1(n_561),
.B2(n_562),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4317),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_L g4427 ( 
.A1(n_4204),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4268),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4269),
.Y(n_4429)
);

AOI22xp33_ASAP7_75t_L g4430 ( 
.A1(n_4266),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_4430)
);

AOI211xp5_ASAP7_75t_SL g4431 ( 
.A1(n_4326),
.A2(n_566),
.B(n_567),
.C(n_568),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_L g4432 ( 
.A1(n_4233),
.A2(n_569),
.B1(n_571),
.B2(n_572),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4269),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_4221),
.B(n_569),
.Y(n_4434)
);

OAI21xp5_ASAP7_75t_SL g4435 ( 
.A1(n_4256),
.A2(n_571),
.B(n_572),
.Y(n_4435)
);

AOI22xp33_ASAP7_75t_L g4436 ( 
.A1(n_4196),
.A2(n_573),
.B1(n_574),
.B2(n_576),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4202),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_SL g4438 ( 
.A1(n_4323),
.A2(n_573),
.B1(n_574),
.B2(n_576),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4230),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4230),
.Y(n_4440)
);

AOI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_4324),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4251),
.Y(n_4442)
);

HB1xp67_ASAP7_75t_L g4443 ( 
.A(n_4186),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4252),
.Y(n_4444)
);

AOI22xp33_ASAP7_75t_L g4445 ( 
.A1(n_4329),
.A2(n_577),
.B1(n_580),
.B2(n_581),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4322),
.B(n_4191),
.Y(n_4446)
);

OAI21xp5_ASAP7_75t_SL g4447 ( 
.A1(n_4297),
.A2(n_4308),
.B(n_4283),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_4284),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_4448)
);

AOI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4284),
.A2(n_583),
.B1(n_584),
.B2(n_585),
.Y(n_4449)
);

INVx4_ASAP7_75t_L g4450 ( 
.A(n_4320),
.Y(n_4450)
);

HB1xp67_ASAP7_75t_L g4451 ( 
.A(n_4186),
.Y(n_4451)
);

INVx4_ASAP7_75t_L g4452 ( 
.A(n_4289),
.Y(n_4452)
);

OAI22xp33_ASAP7_75t_L g4453 ( 
.A1(n_4211),
.A2(n_584),
.B1(n_586),
.B2(n_587),
.Y(n_4453)
);

AOI22xp33_ASAP7_75t_SL g4454 ( 
.A1(n_4219),
.A2(n_586),
.B1(n_587),
.B2(n_588),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4242),
.Y(n_4455)
);

INVx3_ASAP7_75t_L g4456 ( 
.A(n_4289),
.Y(n_4456)
);

OAI21xp33_ASAP7_75t_L g4457 ( 
.A1(n_4267),
.A2(n_588),
.B(n_589),
.Y(n_4457)
);

OAI22xp5_ASAP7_75t_L g4458 ( 
.A1(n_4225),
.A2(n_589),
.B1(n_590),
.B2(n_591),
.Y(n_4458)
);

OAI22xp5_ASAP7_75t_L g4459 ( 
.A1(n_4305),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_4459)
);

AOI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4265),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4242),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4255),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_4281),
.B(n_597),
.Y(n_4463)
);

OAI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4263),
.A2(n_4316),
.B1(n_4247),
.B2(n_4189),
.Y(n_4464)
);

OAI21xp33_ASAP7_75t_L g4465 ( 
.A1(n_4222),
.A2(n_597),
.B(n_598),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_L g4466 ( 
.A1(n_4312),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.Y(n_4466)
);

OAI22xp5_ASAP7_75t_L g4467 ( 
.A1(n_4245),
.A2(n_599),
.B1(n_600),
.B2(n_601),
.Y(n_4467)
);

AOI22xp33_ASAP7_75t_L g4468 ( 
.A1(n_4237),
.A2(n_602),
.B1(n_603),
.B2(n_604),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4186),
.B(n_602),
.Y(n_4469)
);

OAI22xp5_ASAP7_75t_L g4470 ( 
.A1(n_4236),
.A2(n_604),
.B1(n_605),
.B2(n_606),
.Y(n_4470)
);

INVx4_ASAP7_75t_L g4471 ( 
.A(n_4307),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4388),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4331),
.B(n_4244),
.Y(n_4473)
);

AND2x2_ASAP7_75t_L g4474 ( 
.A(n_4331),
.B(n_4304),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4332),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4371),
.B(n_4254),
.Y(n_4476)
);

INVx3_ASAP7_75t_L g4477 ( 
.A(n_4405),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_4371),
.B(n_4255),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4333),
.Y(n_4479)
);

BUFx2_ASAP7_75t_SL g4480 ( 
.A(n_4405),
.Y(n_4480)
);

OR2x2_ASAP7_75t_L g4481 ( 
.A(n_4336),
.B(n_4216),
.Y(n_4481)
);

INVx2_ASAP7_75t_SL g4482 ( 
.A(n_4412),
.Y(n_4482)
);

HB1xp67_ASAP7_75t_L g4483 ( 
.A(n_4443),
.Y(n_4483)
);

HB1xp67_ASAP7_75t_L g4484 ( 
.A(n_4451),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4388),
.Y(n_4485)
);

INVx3_ASAP7_75t_L g4486 ( 
.A(n_4388),
.Y(n_4486)
);

OR2x2_ASAP7_75t_L g4487 ( 
.A(n_4378),
.B(n_4216),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4397),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4341),
.Y(n_4489)
);

BUFx3_ASAP7_75t_L g4490 ( 
.A(n_4340),
.Y(n_4490)
);

NAND3x1_ASAP7_75t_L g4491 ( 
.A(n_4469),
.B(n_4243),
.C(n_4246),
.Y(n_4491)
);

HB1xp67_ASAP7_75t_L g4492 ( 
.A(n_4352),
.Y(n_4492)
);

HB1xp67_ASAP7_75t_L g4493 ( 
.A(n_4343),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4397),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4397),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4365),
.B(n_4206),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_4349),
.B(n_4206),
.Y(n_4497)
);

INVxp67_ASAP7_75t_L g4498 ( 
.A(n_4456),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4346),
.Y(n_4499)
);

AND2x2_ASAP7_75t_L g4500 ( 
.A(n_4348),
.B(n_4306),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4361),
.Y(n_4501)
);

AO21x2_ASAP7_75t_L g4502 ( 
.A1(n_4386),
.A2(n_4207),
.B(n_4239),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4456),
.B(n_4306),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4413),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_4471),
.B(n_4292),
.Y(n_4505)
);

AOI21x1_ASAP7_75t_L g4506 ( 
.A1(n_4420),
.A2(n_4272),
.B(n_4258),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4428),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_4450),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4429),
.Y(n_4509)
);

HB1xp67_ASAP7_75t_L g4510 ( 
.A(n_4363),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4452),
.B(n_4270),
.Y(n_4511)
);

OAI21x1_ASAP7_75t_L g4512 ( 
.A1(n_4411),
.A2(n_4437),
.B(n_4402),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4450),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4433),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4452),
.B(n_4292),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4439),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_4364),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4347),
.B(n_4206),
.Y(n_4518)
);

BUFx2_ASAP7_75t_L g4519 ( 
.A(n_4359),
.Y(n_4519)
);

OAI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4335),
.A2(n_4216),
.B1(n_4328),
.B2(n_4243),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4355),
.B(n_4447),
.Y(n_4521)
);

AO21x1_ASAP7_75t_SL g4522 ( 
.A1(n_4353),
.A2(n_4328),
.B(n_4227),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4360),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4395),
.Y(n_4524)
);

OA21x2_ASAP7_75t_L g4525 ( 
.A1(n_4369),
.A2(n_4356),
.B(n_4447),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4440),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4338),
.B(n_4328),
.Y(n_4527)
);

OAI21xp5_ASAP7_75t_L g4528 ( 
.A1(n_4368),
.A2(n_4290),
.B(n_4311),
.Y(n_4528)
);

INVx2_ASAP7_75t_SL g4529 ( 
.A(n_4407),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4446),
.B(n_4227),
.Y(n_4530)
);

INVxp67_ASAP7_75t_L g4531 ( 
.A(n_4398),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4402),
.B(n_4227),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4396),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4455),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4461),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4462),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_4418),
.Y(n_4537)
);

AO21x2_ASAP7_75t_L g4538 ( 
.A1(n_4417),
.A2(n_4432),
.B(n_4453),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4423),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_4442),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4444),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4370),
.Y(n_4542)
);

INVx2_ASAP7_75t_SL g4543 ( 
.A(n_4407),
.Y(n_4543)
);

INVxp67_ASAP7_75t_L g4544 ( 
.A(n_4338),
.Y(n_4544)
);

INVx4_ASAP7_75t_L g4545 ( 
.A(n_4340),
.Y(n_4545)
);

AOI22xp33_ASAP7_75t_L g4546 ( 
.A1(n_4342),
.A2(n_4302),
.B1(n_4287),
.B2(n_4279),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4381),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4384),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4345),
.B(n_4318),
.Y(n_4549)
);

AOI221xp5_ASAP7_75t_L g4550 ( 
.A1(n_4334),
.A2(n_4342),
.B1(n_4351),
.B2(n_4362),
.C(n_4409),
.Y(n_4550)
);

BUFx3_ASAP7_75t_L g4551 ( 
.A(n_4340),
.Y(n_4551)
);

AND2x4_ASAP7_75t_L g4552 ( 
.A(n_4385),
.B(n_4243),
.Y(n_4552)
);

OR2x6_ASAP7_75t_L g4553 ( 
.A(n_4435),
.B(n_4246),
.Y(n_4553)
);

OR2x6_ASAP7_75t_L g4554 ( 
.A(n_4435),
.B(n_4409),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4394),
.Y(n_4555)
);

INVx3_ASAP7_75t_L g4556 ( 
.A(n_4375),
.Y(n_4556)
);

OAI221xp5_ASAP7_75t_L g4557 ( 
.A1(n_4351),
.A2(n_4250),
.B1(n_4246),
.B2(n_4303),
.C(n_608),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4401),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_4354),
.A2(n_4250),
.B1(n_4303),
.B2(n_607),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4408),
.B(n_4250),
.Y(n_4560)
);

OAI21x1_ASAP7_75t_L g4561 ( 
.A1(n_4392),
.A2(n_4303),
.B(n_606),
.Y(n_4561)
);

OAI21x1_ASAP7_75t_L g4562 ( 
.A1(n_4410),
.A2(n_4366),
.B(n_4357),
.Y(n_4562)
);

INVx3_ASAP7_75t_L g4563 ( 
.A(n_4407),
.Y(n_4563)
);

BUFx2_ASAP7_75t_L g4564 ( 
.A(n_4339),
.Y(n_4564)
);

BUFx6f_ASAP7_75t_L g4565 ( 
.A(n_4350),
.Y(n_4565)
);

AO21x2_ASAP7_75t_L g4566 ( 
.A1(n_4417),
.A2(n_605),
.B(n_608),
.Y(n_4566)
);

INVx3_ASAP7_75t_L g4567 ( 
.A(n_4471),
.Y(n_4567)
);

BUFx5_ASAP7_75t_L g4568 ( 
.A(n_4391),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_4358),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4337),
.B(n_609),
.Y(n_4570)
);

BUFx3_ASAP7_75t_L g4571 ( 
.A(n_4414),
.Y(n_4571)
);

BUFx6f_ASAP7_75t_L g4572 ( 
.A(n_4399),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4367),
.B(n_610),
.Y(n_4573)
);

AND2x4_ASAP7_75t_L g4574 ( 
.A(n_4372),
.B(n_610),
.Y(n_4574)
);

INVx3_ASAP7_75t_L g4575 ( 
.A(n_4390),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4432),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4464),
.B(n_611),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4403),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4377),
.B(n_611),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_4406),
.B(n_612),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4463),
.Y(n_4581)
);

INVx2_ASAP7_75t_SL g4582 ( 
.A(n_4434),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4436),
.B(n_612),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4373),
.B(n_613),
.Y(n_4584)
);

AO21x2_ASAP7_75t_L g4585 ( 
.A1(n_4344),
.A2(n_614),
.B(n_615),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4427),
.B(n_615),
.Y(n_4586)
);

AO21x1_ASAP7_75t_SL g4587 ( 
.A1(n_4421),
.A2(n_616),
.B(n_617),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4362),
.B(n_616),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4425),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4465),
.Y(n_4590)
);

AOI21xp5_ASAP7_75t_SL g4591 ( 
.A1(n_4467),
.A2(n_619),
.B(n_620),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4470),
.Y(n_4592)
);

INVx3_ASAP7_75t_L g4593 ( 
.A(n_4431),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4404),
.B(n_619),
.Y(n_4594)
);

HB1xp67_ASAP7_75t_L g4595 ( 
.A(n_4431),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4458),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4387),
.B(n_620),
.Y(n_4597)
);

INVx2_ASAP7_75t_SL g4598 ( 
.A(n_4459),
.Y(n_4598)
);

INVxp67_ASAP7_75t_SL g4599 ( 
.A(n_4416),
.Y(n_4599)
);

OR2x6_ASAP7_75t_L g4600 ( 
.A(n_4416),
.B(n_621),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4424),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4419),
.Y(n_4602)
);

BUFx2_ASAP7_75t_L g4603 ( 
.A(n_4374),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4448),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4486),
.Y(n_4605)
);

INVx2_ASAP7_75t_SL g4606 ( 
.A(n_4477),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4492),
.Y(n_4607)
);

OAI21x1_ASAP7_75t_L g4608 ( 
.A1(n_4512),
.A2(n_4562),
.B(n_4506),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4595),
.B(n_4400),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4492),
.Y(n_4610)
);

BUFx6f_ASAP7_75t_L g4611 ( 
.A(n_4490),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4482),
.B(n_4454),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4482),
.B(n_4382),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4493),
.Y(n_4614)
);

BUFx3_ASAP7_75t_L g4615 ( 
.A(n_4571),
.Y(n_4615)
);

BUFx2_ASAP7_75t_L g4616 ( 
.A(n_4593),
.Y(n_4616)
);

AOI221xp5_ASAP7_75t_L g4617 ( 
.A1(n_4550),
.A2(n_4400),
.B1(n_4457),
.B2(n_4389),
.C(n_4380),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4486),
.B(n_4563),
.Y(n_4618)
);

OR2x2_ASAP7_75t_L g4619 ( 
.A(n_4576),
.B(n_4449),
.Y(n_4619)
);

BUFx6f_ASAP7_75t_L g4620 ( 
.A(n_4490),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4486),
.B(n_4438),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_4567),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4567),
.Y(n_4623)
);

OR2x2_ASAP7_75t_L g4624 ( 
.A(n_4524),
.B(n_4393),
.Y(n_4624)
);

BUFx12f_ASAP7_75t_L g4625 ( 
.A(n_4545),
.Y(n_4625)
);

BUFx3_ASAP7_75t_L g4626 ( 
.A(n_4571),
.Y(n_4626)
);

INVxp67_ASAP7_75t_L g4627 ( 
.A(n_4595),
.Y(n_4627)
);

INVx2_ASAP7_75t_SL g4628 ( 
.A(n_4477),
.Y(n_4628)
);

NOR2xp33_ASAP7_75t_L g4629 ( 
.A(n_4545),
.B(n_4445),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_4572),
.Y(n_4630)
);

AND2x4_ASAP7_75t_L g4631 ( 
.A(n_4477),
.B(n_4430),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4567),
.Y(n_4632)
);

AND2x4_ASAP7_75t_L g4633 ( 
.A(n_4472),
.B(n_4376),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4493),
.Y(n_4634)
);

AND2x2_ASAP7_75t_L g4635 ( 
.A(n_4563),
.B(n_4466),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4563),
.B(n_4468),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4593),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4472),
.B(n_4415),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4593),
.B(n_4441),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4510),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4485),
.B(n_4488),
.Y(n_4641)
);

INVxp67_ASAP7_75t_L g4642 ( 
.A(n_4480),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4485),
.B(n_4488),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4551),
.Y(n_4644)
);

BUFx6f_ASAP7_75t_L g4645 ( 
.A(n_4551),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4510),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_SL g4647 ( 
.A(n_4572),
.B(n_4460),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4572),
.Y(n_4648)
);

OA21x2_ASAP7_75t_L g4649 ( 
.A1(n_4562),
.A2(n_4426),
.B(n_4422),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4572),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4483),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4565),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4483),
.Y(n_4653)
);

AND2x4_ASAP7_75t_L g4654 ( 
.A(n_4494),
.B(n_4379),
.Y(n_4654)
);

BUFx2_ASAP7_75t_L g4655 ( 
.A(n_4553),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4484),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4524),
.B(n_4533),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4494),
.B(n_4495),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4495),
.B(n_4383),
.Y(n_4659)
);

NAND3xp33_ASAP7_75t_L g4660 ( 
.A(n_4497),
.B(n_622),
.C(n_623),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4565),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4529),
.B(n_622),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4565),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4565),
.Y(n_4664)
);

OAI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4554),
.A2(n_4553),
.B1(n_4599),
.B2(n_4559),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4484),
.Y(n_4666)
);

HB1xp67_ASAP7_75t_L g4667 ( 
.A(n_4498),
.Y(n_4667)
);

BUFx3_ASAP7_75t_L g4668 ( 
.A(n_4519),
.Y(n_4668)
);

NOR2x1_ASAP7_75t_L g4669 ( 
.A(n_4585),
.B(n_624),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4517),
.Y(n_4670)
);

CKINVDCx5p33_ASAP7_75t_R g4671 ( 
.A(n_4556),
.Y(n_4671)
);

INVx3_ASAP7_75t_L g4672 ( 
.A(n_4545),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4517),
.Y(n_4673)
);

HB1xp67_ASAP7_75t_L g4674 ( 
.A(n_4552),
.Y(n_4674)
);

BUFx6f_ASAP7_75t_L g4675 ( 
.A(n_4588),
.Y(n_4675)
);

INVx2_ASAP7_75t_L g4676 ( 
.A(n_4569),
.Y(n_4676)
);

HB1xp67_ASAP7_75t_L g4677 ( 
.A(n_4552),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4529),
.B(n_624),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4535),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4543),
.B(n_4508),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4543),
.B(n_625),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4535),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4508),
.B(n_625),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4475),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4552),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4569),
.Y(n_4686)
);

CKINVDCx11_ASAP7_75t_R g4687 ( 
.A(n_4564),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4513),
.B(n_626),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4568),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4479),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4513),
.B(n_626),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4568),
.Y(n_4692)
);

OA21x2_ASAP7_75t_L g4693 ( 
.A1(n_4521),
.A2(n_627),
.B(n_628),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4474),
.B(n_629),
.Y(n_4694)
);

INVx2_ASAP7_75t_L g4695 ( 
.A(n_4568),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4489),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4568),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4499),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4501),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4533),
.B(n_630),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4530),
.B(n_631),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4568),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4538),
.B(n_631),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4530),
.B(n_632),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4511),
.B(n_632),
.Y(n_4705)
);

HB1xp67_ASAP7_75t_L g4706 ( 
.A(n_4560),
.Y(n_4706)
);

INVx2_ASAP7_75t_R g4707 ( 
.A(n_4573),
.Y(n_4707)
);

INVx2_ASAP7_75t_SL g4708 ( 
.A(n_4611),
.Y(n_4708)
);

BUFx6f_ASAP7_75t_L g4709 ( 
.A(n_4625),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4668),
.B(n_4556),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4703),
.Y(n_4711)
);

INVx4_ASAP7_75t_L g4712 ( 
.A(n_4671),
.Y(n_4712)
);

HB1xp67_ASAP7_75t_L g4713 ( 
.A(n_4616),
.Y(n_4713)
);

NAND2x1_ASAP7_75t_L g4714 ( 
.A(n_4703),
.B(n_4553),
.Y(n_4714)
);

INVx4_ASAP7_75t_L g4715 ( 
.A(n_4671),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4616),
.Y(n_4716)
);

AND2x4_ASAP7_75t_L g4717 ( 
.A(n_4606),
.B(n_4556),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4627),
.B(n_4538),
.Y(n_4718)
);

INVx3_ASAP7_75t_L g4719 ( 
.A(n_4625),
.Y(n_4719)
);

INVxp67_ASAP7_75t_SL g4720 ( 
.A(n_4669),
.Y(n_4720)
);

BUFx2_ASAP7_75t_L g4721 ( 
.A(n_4655),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4634),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4611),
.Y(n_4723)
);

INVx3_ASAP7_75t_L g4724 ( 
.A(n_4611),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4634),
.Y(n_4725)
);

INVx4_ASAP7_75t_L g4726 ( 
.A(n_4611),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4611),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4668),
.B(n_4515),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4640),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4640),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4637),
.B(n_4531),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4637),
.B(n_4532),
.Y(n_4732)
);

OR2x2_ASAP7_75t_L g4733 ( 
.A(n_4609),
.B(n_4525),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4612),
.B(n_4532),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4620),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4707),
.B(n_4525),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4620),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4674),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4707),
.B(n_4525),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4646),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4646),
.Y(n_4741)
);

BUFx2_ASAP7_75t_L g4742 ( 
.A(n_4655),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4620),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4651),
.Y(n_4744)
);

HB1xp67_ASAP7_75t_L g4745 ( 
.A(n_4677),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4651),
.Y(n_4746)
);

OR2x2_ASAP7_75t_L g4747 ( 
.A(n_4619),
.B(n_4607),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4653),
.Y(n_4748)
);

BUFx6f_ASAP7_75t_L g4749 ( 
.A(n_4687),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4620),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4620),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4653),
.Y(n_4752)
);

BUFx2_ASAP7_75t_L g4753 ( 
.A(n_4672),
.Y(n_4753)
);

AND2x4_ASAP7_75t_L g4754 ( 
.A(n_4606),
.B(n_4560),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4644),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4644),
.Y(n_4756)
);

INVx3_ASAP7_75t_L g4757 ( 
.A(n_4644),
.Y(n_4757)
);

BUFx2_ASAP7_75t_L g4758 ( 
.A(n_4672),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4612),
.B(n_4603),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4644),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4613),
.B(n_4598),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4613),
.B(n_4500),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4656),
.Y(n_4763)
);

BUFx2_ASAP7_75t_L g4764 ( 
.A(n_4672),
.Y(n_4764)
);

OR2x2_ASAP7_75t_L g4765 ( 
.A(n_4619),
.B(n_4544),
.Y(n_4765)
);

AOI22xp33_ASAP7_75t_L g4766 ( 
.A1(n_4665),
.A2(n_4649),
.B1(n_4675),
.B2(n_4554),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4656),
.Y(n_4767)
);

INVxp67_ASAP7_75t_R g4768 ( 
.A(n_4701),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4644),
.Y(n_4769)
);

INVx1_ASAP7_75t_SL g4770 ( 
.A(n_4736),
.Y(n_4770)
);

NAND3xp33_ASAP7_75t_L g4771 ( 
.A(n_4766),
.B(n_4675),
.C(n_4617),
.Y(n_4771)
);

NOR2x1_ASAP7_75t_L g4772 ( 
.A(n_4736),
.B(n_4615),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4749),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4713),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4716),
.Y(n_4775)
);

INVxp67_ASAP7_75t_L g4776 ( 
.A(n_4749),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4749),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_4749),
.Y(n_4778)
);

HB1xp67_ASAP7_75t_L g4779 ( 
.A(n_4753),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4749),
.Y(n_4780)
);

INVxp67_ASAP7_75t_L g4781 ( 
.A(n_4720),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4716),
.Y(n_4782)
);

OAI21xp5_ASAP7_75t_SL g4783 ( 
.A1(n_4718),
.A2(n_4639),
.B(n_4527),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_SL g4784 ( 
.A(n_4710),
.B(n_4645),
.Y(n_4784)
);

AND2x4_ASAP7_75t_L g4785 ( 
.A(n_4708),
.B(n_4615),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4761),
.B(n_4676),
.Y(n_4786)
);

OR2x2_ASAP7_75t_L g4787 ( 
.A(n_4759),
.B(n_4676),
.Y(n_4787)
);

AND2x4_ASAP7_75t_L g4788 ( 
.A(n_4708),
.B(n_4626),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4738),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4745),
.Y(n_4790)
);

OR2x2_ASAP7_75t_L g4791 ( 
.A(n_4747),
.B(n_4765),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4753),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4711),
.B(n_4701),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4747),
.B(n_4686),
.Y(n_4794)
);

AOI22xp33_ASAP7_75t_L g4795 ( 
.A1(n_4710),
.A2(n_4675),
.B1(n_4649),
.B2(n_4554),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4711),
.B(n_4704),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4758),
.Y(n_4797)
);

INVx2_ASAP7_75t_SL g4798 ( 
.A(n_4717),
.Y(n_4798)
);

OR2x2_ASAP7_75t_L g4799 ( 
.A(n_4765),
.B(n_4686),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4768),
.B(n_4626),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4758),
.Y(n_4801)
);

OR2x2_ASAP7_75t_L g4802 ( 
.A(n_4718),
.B(n_4667),
.Y(n_4802)
);

AND2x2_ASAP7_75t_L g4803 ( 
.A(n_4768),
.B(n_4642),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4721),
.B(n_4704),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4721),
.B(n_4675),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4742),
.B(n_4675),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4742),
.B(n_4693),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4764),
.Y(n_4808)
);

AND2x2_ASAP7_75t_L g4809 ( 
.A(n_4762),
.B(n_4621),
.Y(n_4809)
);

INVx2_ASAP7_75t_SL g4810 ( 
.A(n_4717),
.Y(n_4810)
);

NOR2x1_ASAP7_75t_SL g4811 ( 
.A(n_4739),
.B(n_4585),
.Y(n_4811)
);

NOR2xp33_ASAP7_75t_R g4812 ( 
.A(n_4719),
.B(n_4645),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4764),
.Y(n_4813)
);

BUFx2_ASAP7_75t_L g4814 ( 
.A(n_4717),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4733),
.B(n_4693),
.Y(n_4815)
);

BUFx3_ASAP7_75t_L g4816 ( 
.A(n_4717),
.Y(n_4816)
);

AND2x4_ASAP7_75t_SL g4817 ( 
.A(n_4712),
.B(n_4645),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4762),
.B(n_4621),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4744),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4733),
.B(n_4693),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4734),
.B(n_4630),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4734),
.B(n_4693),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4726),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4739),
.B(n_4610),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_SL g4825 ( 
.A(n_4770),
.B(n_4712),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4779),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4814),
.Y(n_4827)
);

OR2x2_ASAP7_75t_L g4828 ( 
.A(n_4770),
.B(n_4714),
.Y(n_4828)
);

NOR2xp33_ASAP7_75t_L g4829 ( 
.A(n_4776),
.B(n_4712),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4809),
.B(n_4728),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4792),
.Y(n_4831)
);

INVx3_ASAP7_75t_L g4832 ( 
.A(n_4816),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4797),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4798),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4818),
.B(n_4728),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4801),
.Y(n_4836)
);

INVx2_ASAP7_75t_L g4837 ( 
.A(n_4810),
.Y(n_4837)
);

NOR2xp33_ASAP7_75t_L g4838 ( 
.A(n_4773),
.B(n_4715),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4813),
.Y(n_4839)
);

BUFx2_ASAP7_75t_L g4840 ( 
.A(n_4772),
.Y(n_4840)
);

HB1xp67_ASAP7_75t_L g4841 ( 
.A(n_4785),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4777),
.B(n_4618),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4808),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4778),
.B(n_4731),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4780),
.B(n_4618),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4794),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4800),
.B(n_4652),
.Y(n_4847)
);

OR2x2_ASAP7_75t_L g4848 ( 
.A(n_4791),
.B(n_4714),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4805),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4803),
.B(n_4652),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4785),
.B(n_4788),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4805),
.Y(n_4852)
);

BUFx2_ASAP7_75t_L g4853 ( 
.A(n_4812),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4788),
.B(n_4661),
.Y(n_4854)
);

AOI22xp5_ASAP7_75t_L g4855 ( 
.A1(n_4771),
.A2(n_4649),
.B1(n_4496),
.B2(n_4520),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4817),
.B(n_4661),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4806),
.Y(n_4857)
);

AND2x2_ASAP7_75t_SL g4858 ( 
.A(n_4795),
.B(n_4715),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4774),
.B(n_4731),
.Y(n_4859)
);

NAND4xp25_ASAP7_75t_L g4860 ( 
.A(n_4821),
.B(n_4715),
.C(n_4719),
.D(n_4629),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4789),
.B(n_4663),
.Y(n_4861)
);

HB1xp67_ASAP7_75t_L g4862 ( 
.A(n_4806),
.Y(n_4862)
);

AND2x4_ASAP7_75t_L g4863 ( 
.A(n_4823),
.B(n_4726),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4799),
.Y(n_4864)
);

AND2x2_ASAP7_75t_L g4865 ( 
.A(n_4790),
.B(n_4663),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4781),
.A2(n_4649),
.B1(n_4608),
.B2(n_4600),
.Y(n_4866)
);

BUFx2_ASAP7_75t_SL g4867 ( 
.A(n_4784),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4841),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4828),
.Y(n_4869)
);

HB1xp67_ASAP7_75t_L g4870 ( 
.A(n_4840),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4828),
.Y(n_4871)
);

OR2x2_ASAP7_75t_L g4872 ( 
.A(n_4844),
.B(n_4804),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4834),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4834),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4837),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4830),
.B(n_4715),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4837),
.Y(n_4877)
);

AND2x4_ASAP7_75t_L g4878 ( 
.A(n_4832),
.B(n_4726),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4830),
.B(n_4680),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4840),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4855),
.B(n_4783),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4827),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4862),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4850),
.B(n_4680),
.Y(n_4884)
);

AOI21xp33_ASAP7_75t_L g4885 ( 
.A1(n_4825),
.A2(n_4820),
.B(n_4815),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4848),
.Y(n_4886)
);

NOR2xp33_ASAP7_75t_L g4887 ( 
.A(n_4860),
.B(n_4709),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4861),
.B(n_4783),
.Y(n_4888)
);

AND2x4_ASAP7_75t_SL g4889 ( 
.A(n_4856),
.B(n_4709),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4850),
.B(n_4719),
.Y(n_4890)
);

OR2x6_ASAP7_75t_L g4891 ( 
.A(n_4825),
.B(n_4709),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4848),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4861),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_SL g4894 ( 
.A(n_4853),
.B(n_4645),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_SL g4895 ( 
.A(n_4853),
.B(n_4645),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4865),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4847),
.B(n_4636),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4870),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4870),
.B(n_4842),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4897),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4879),
.B(n_4847),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4886),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4892),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4884),
.B(n_4842),
.Y(n_4904)
);

OR2x2_ASAP7_75t_L g4905 ( 
.A(n_4868),
.B(n_4804),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4890),
.B(n_4854),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4878),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4893),
.B(n_4854),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4896),
.B(n_4845),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4869),
.B(n_4845),
.Y(n_4910)
);

OR2x2_ASAP7_75t_L g4911 ( 
.A(n_4888),
.B(n_4793),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4871),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4876),
.B(n_4856),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4873),
.Y(n_4914)
);

INVx1_ASAP7_75t_SL g4915 ( 
.A(n_4889),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4874),
.Y(n_4916)
);

OR2x2_ASAP7_75t_L g4917 ( 
.A(n_4888),
.B(n_4793),
.Y(n_4917)
);

OR2x2_ASAP7_75t_L g4918 ( 
.A(n_4872),
.B(n_4796),
.Y(n_4918)
);

INVx2_ASAP7_75t_SL g4919 ( 
.A(n_4878),
.Y(n_4919)
);

AND2x2_ASAP7_75t_L g4920 ( 
.A(n_4887),
.B(n_4858),
.Y(n_4920)
);

AND2x2_ASAP7_75t_L g4921 ( 
.A(n_4901),
.B(n_4858),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4899),
.A2(n_4881),
.B(n_4885),
.Y(n_4922)
);

NAND2x1p5_ASAP7_75t_L g4923 ( 
.A(n_4915),
.B(n_4709),
.Y(n_4923)
);

INVxp67_ASAP7_75t_L g4924 ( 
.A(n_4899),
.Y(n_4924)
);

OR2x2_ASAP7_75t_L g4925 ( 
.A(n_4906),
.B(n_4835),
.Y(n_4925)
);

NOR2x1_ASAP7_75t_R g4926 ( 
.A(n_4919),
.B(n_4709),
.Y(n_4926)
);

INVxp67_ASAP7_75t_L g4927 ( 
.A(n_4913),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4904),
.B(n_4832),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4908),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4915),
.B(n_4832),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4910),
.Y(n_4931)
);

INVx2_ASAP7_75t_SL g4932 ( 
.A(n_4907),
.Y(n_4932)
);

OR2x2_ASAP7_75t_L g4933 ( 
.A(n_4910),
.B(n_4796),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4898),
.Y(n_4934)
);

OR2x2_ASAP7_75t_L g4935 ( 
.A(n_4909),
.B(n_4859),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4900),
.B(n_4723),
.Y(n_4936)
);

INVxp67_ASAP7_75t_L g4937 ( 
.A(n_4909),
.Y(n_4937)
);

OAI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4920),
.A2(n_4881),
.B(n_4866),
.Y(n_4938)
);

NOR2xp33_ASAP7_75t_SL g4939 ( 
.A(n_4926),
.B(n_4928),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4930),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4923),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4927),
.A2(n_4851),
.B1(n_4787),
.B2(n_4664),
.Y(n_4942)
);

INVx1_ASAP7_75t_SL g4943 ( 
.A(n_4921),
.Y(n_4943)
);

OR2x2_ASAP7_75t_L g4944 ( 
.A(n_4932),
.B(n_4867),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4934),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4936),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4938),
.B(n_4867),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4934),
.Y(n_4948)
);

OAI22xp33_ASAP7_75t_L g4949 ( 
.A1(n_4922),
.A2(n_4820),
.B1(n_4815),
.B2(n_4807),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4924),
.B(n_4865),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4937),
.B(n_4826),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4944),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4947),
.B(n_4829),
.Y(n_4953)
);

AOI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4943),
.A2(n_4838),
.B1(n_4664),
.B2(n_4628),
.Y(n_4954)
);

OAI21xp33_ASAP7_75t_SL g4955 ( 
.A1(n_4950),
.A2(n_4608),
.B(n_4807),
.Y(n_4955)
);

HB1xp67_ASAP7_75t_L g4956 ( 
.A(n_4941),
.Y(n_4956)
);

OAI22xp5_ASAP7_75t_L g4957 ( 
.A1(n_4943),
.A2(n_4650),
.B1(n_4648),
.B2(n_4786),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4942),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4940),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4951),
.Y(n_4960)
);

AOI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_4953),
.A2(n_4939),
.B1(n_4843),
.B2(n_4882),
.Y(n_4961)
);

OAI221xp5_ASAP7_75t_L g4962 ( 
.A1(n_4954),
.A2(n_4939),
.B1(n_4885),
.B2(n_4891),
.C(n_4824),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4957),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4956),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4958),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4952),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4959),
.B(n_4863),
.Y(n_4967)
);

AOI211xp5_ASAP7_75t_L g4968 ( 
.A1(n_4955),
.A2(n_4949),
.B(n_4895),
.C(n_4894),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4960),
.Y(n_4969)
);

AOI221xp5_ASAP7_75t_L g4970 ( 
.A1(n_4957),
.A2(n_4880),
.B1(n_4824),
.B2(n_4877),
.C(n_4875),
.Y(n_4970)
);

OAI21xp33_ASAP7_75t_L g4971 ( 
.A1(n_4953),
.A2(n_4925),
.B(n_4822),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4954),
.Y(n_4972)
);

OR2x2_ASAP7_75t_L g4973 ( 
.A(n_4957),
.B(n_4802),
.Y(n_4973)
);

AOI221x1_ASAP7_75t_L g4974 ( 
.A1(n_4958),
.A2(n_4912),
.B1(n_4914),
.B2(n_4916),
.C(n_4931),
.Y(n_4974)
);

NOR2xp33_ASAP7_75t_L g4975 ( 
.A(n_4962),
.B(n_4849),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4973),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4964),
.B(n_4864),
.Y(n_4977)
);

AOI33xp33_ASAP7_75t_L g4978 ( 
.A1(n_4972),
.A2(n_4836),
.A3(n_4839),
.B1(n_4833),
.B2(n_4831),
.B3(n_4883),
.Y(n_4978)
);

A2O1A1Ixp33_ASAP7_75t_L g4979 ( 
.A1(n_4971),
.A2(n_4724),
.B(n_4757),
.C(n_4727),
.Y(n_4979)
);

O2A1O1Ixp33_ASAP7_75t_SL g4980 ( 
.A1(n_4968),
.A2(n_4905),
.B(n_4917),
.C(n_4911),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4967),
.Y(n_4981)
);

AOI22xp5_ASAP7_75t_L g4982 ( 
.A1(n_4961),
.A2(n_4891),
.B1(n_4857),
.B2(n_4852),
.Y(n_4982)
);

OR2x2_ASAP7_75t_L g4983 ( 
.A(n_4963),
.B(n_4891),
.Y(n_4983)
);

AOI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4966),
.A2(n_4918),
.B(n_4933),
.Y(n_4984)
);

AOI21xp5_ASAP7_75t_L g4985 ( 
.A1(n_4970),
.A2(n_4935),
.B(n_4945),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4965),
.B(n_4863),
.Y(n_4986)
);

OAI22xp33_ASAP7_75t_L g4987 ( 
.A1(n_4974),
.A2(n_4757),
.B1(n_4724),
.B2(n_4622),
.Y(n_4987)
);

AOI222xp33_ASAP7_75t_L g4988 ( 
.A1(n_4969),
.A2(n_4811),
.B1(n_4775),
.B2(n_4782),
.C1(n_4846),
.C2(n_4902),
.Y(n_4988)
);

INVx1_ASAP7_75t_SL g4989 ( 
.A(n_4973),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4964),
.B(n_4863),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4973),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4973),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4973),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4968),
.B(n_4903),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4973),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_4973),
.Y(n_4996)
);

OAI221xp5_ASAP7_75t_L g4997 ( 
.A1(n_4982),
.A2(n_4757),
.B1(n_4724),
.B2(n_4743),
.C(n_4723),
.Y(n_4997)
);

NOR3xp33_ASAP7_75t_L g4998 ( 
.A(n_4976),
.B(n_4929),
.C(n_4946),
.Y(n_4998)
);

OAI22xp5_ASAP7_75t_L g4999 ( 
.A1(n_4982),
.A2(n_4650),
.B1(n_4648),
.B2(n_4727),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4990),
.Y(n_5000)
);

OAI222xp33_ASAP7_75t_L g5001 ( 
.A1(n_4989),
.A2(n_4735),
.B1(n_4743),
.B2(n_4750),
.C1(n_4769),
.C2(n_4751),
.Y(n_5001)
);

NOR2xp33_ASAP7_75t_L g5002 ( 
.A(n_4986),
.B(n_4948),
.Y(n_5002)
);

AOI21xp33_ASAP7_75t_L g5003 ( 
.A1(n_4988),
.A2(n_4737),
.B(n_4735),
.Y(n_5003)
);

AOI22xp5_ASAP7_75t_L g5004 ( 
.A1(n_4992),
.A2(n_4760),
.B1(n_4750),
.B2(n_4769),
.Y(n_5004)
);

OAI221xp5_ASAP7_75t_L g5005 ( 
.A1(n_4979),
.A2(n_4755),
.B1(n_4751),
.B2(n_4737),
.C(n_4756),
.Y(n_5005)
);

OAI221xp5_ASAP7_75t_L g5006 ( 
.A1(n_4994),
.A2(n_4756),
.B1(n_4755),
.B2(n_4760),
.C(n_4763),
.Y(n_5006)
);

OAI21xp5_ASAP7_75t_SL g5007 ( 
.A1(n_4993),
.A2(n_4819),
.B(n_4746),
.Y(n_5007)
);

AOI211x1_ASAP7_75t_L g5008 ( 
.A1(n_4987),
.A2(n_4746),
.B(n_4767),
.C(n_4763),
.Y(n_5008)
);

AOI321xp33_ASAP7_75t_L g5009 ( 
.A1(n_4975),
.A2(n_4744),
.A3(n_4767),
.B1(n_4748),
.B2(n_4752),
.C(n_4722),
.Y(n_5009)
);

AOI221xp5_ASAP7_75t_L g5010 ( 
.A1(n_4980),
.A2(n_4748),
.B1(n_4752),
.B2(n_4722),
.C(n_4729),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4978),
.B(n_4977),
.Y(n_5011)
);

A2O1A1Ixp33_ASAP7_75t_L g5012 ( 
.A1(n_4984),
.A2(n_4730),
.B(n_4741),
.C(n_4740),
.Y(n_5012)
);

OAI21xp33_ASAP7_75t_L g5013 ( 
.A1(n_4995),
.A2(n_4822),
.B(n_4729),
.Y(n_5013)
);

CKINVDCx5p33_ASAP7_75t_R g5014 ( 
.A(n_4991),
.Y(n_5014)
);

AOI222xp33_ASAP7_75t_L g5015 ( 
.A1(n_4996),
.A2(n_4725),
.B1(n_4741),
.B2(n_4740),
.C1(n_4730),
.C2(n_4666),
.Y(n_5015)
);

OAI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4985),
.A2(n_4725),
.B(n_4623),
.Y(n_5016)
);

AOI211xp5_ASAP7_75t_L g5017 ( 
.A1(n_4983),
.A2(n_4622),
.B(n_4623),
.C(n_4632),
.Y(n_5017)
);

OR2x2_ASAP7_75t_L g5018 ( 
.A(n_4981),
.B(n_4632),
.Y(n_5018)
);

OAI22xp5_ASAP7_75t_L g5019 ( 
.A1(n_4982),
.A2(n_4628),
.B1(n_4605),
.B2(n_4614),
.Y(n_5019)
);

AOI21xp33_ASAP7_75t_SL g5020 ( 
.A1(n_4987),
.A2(n_4700),
.B(n_4577),
.Y(n_5020)
);

INVxp67_ASAP7_75t_L g5021 ( 
.A(n_4990),
.Y(n_5021)
);

AOI22xp33_ASAP7_75t_L g5022 ( 
.A1(n_4991),
.A2(n_4732),
.B1(n_4754),
.B2(n_4605),
.Y(n_5022)
);

A2O1A1Ixp33_ASAP7_75t_L g5023 ( 
.A1(n_5013),
.A2(n_4754),
.B(n_4732),
.C(n_4688),
.Y(n_5023)
);

OAI211xp5_ASAP7_75t_L g5024 ( 
.A1(n_5003),
.A2(n_4685),
.B(n_4706),
.C(n_4689),
.Y(n_5024)
);

AO21x1_ASAP7_75t_L g5025 ( 
.A1(n_5002),
.A2(n_4754),
.B(n_4692),
.Y(n_5025)
);

AOI211xp5_ASAP7_75t_L g5026 ( 
.A1(n_5001),
.A2(n_4754),
.B(n_4683),
.C(n_4688),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_5004),
.B(n_5022),
.Y(n_5027)
);

AOI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_5014),
.A2(n_4643),
.B1(n_4641),
.B2(n_4658),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_5000),
.B(n_4641),
.Y(n_5029)
);

AOI21x1_ASAP7_75t_L g5030 ( 
.A1(n_5011),
.A2(n_5018),
.B(n_4999),
.Y(n_5030)
);

NAND3xp33_ASAP7_75t_L g5031 ( 
.A(n_4998),
.B(n_4700),
.C(n_4691),
.Y(n_5031)
);

NOR3xp33_ASAP7_75t_SL g5032 ( 
.A(n_5006),
.B(n_4660),
.C(n_4647),
.Y(n_5032)
);

AOI21xp5_ASAP7_75t_L g5033 ( 
.A1(n_5012),
.A2(n_4691),
.B(n_4683),
.Y(n_5033)
);

OAI21xp33_ASAP7_75t_L g5034 ( 
.A1(n_5021),
.A2(n_4658),
.B(n_4643),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_5020),
.B(n_4631),
.Y(n_5035)
);

NOR3xp33_ASAP7_75t_L g5036 ( 
.A(n_5007),
.B(n_4581),
.C(n_4662),
.Y(n_5036)
);

NOR2xp33_ASAP7_75t_SL g5037 ( 
.A(n_4997),
.B(n_4662),
.Y(n_5037)
);

NOR5xp2_ASAP7_75t_L g5038 ( 
.A(n_5005),
.B(n_4679),
.C(n_4673),
.D(n_4682),
.E(n_4696),
.Y(n_5038)
);

OAI32xp33_ASAP7_75t_L g5039 ( 
.A1(n_5019),
.A2(n_4697),
.A3(n_4702),
.B1(n_4689),
.B2(n_4695),
.Y(n_5039)
);

NOR2xp33_ASAP7_75t_SL g5040 ( 
.A(n_5016),
.B(n_4678),
.Y(n_5040)
);

O2A1O1Ixp33_ASAP7_75t_L g5041 ( 
.A1(n_5010),
.A2(n_4692),
.B(n_4702),
.C(n_4697),
.Y(n_5041)
);

O2A1O1Ixp5_ASAP7_75t_L g5042 ( 
.A1(n_5008),
.A2(n_4695),
.B(n_4682),
.C(n_4673),
.Y(n_5042)
);

OAI221xp5_ASAP7_75t_L g5043 ( 
.A1(n_5009),
.A2(n_4696),
.B1(n_4690),
.B2(n_4698),
.C(n_4684),
.Y(n_5043)
);

AOI221xp5_ASAP7_75t_L g5044 ( 
.A1(n_5017),
.A2(n_4678),
.B1(n_4681),
.B2(n_4690),
.C(n_4679),
.Y(n_5044)
);

AOI22xp33_ASAP7_75t_SL g5045 ( 
.A1(n_5015),
.A2(n_4681),
.B1(n_4631),
.B2(n_4573),
.Y(n_5045)
);

OAI21xp33_ASAP7_75t_L g5046 ( 
.A1(n_5022),
.A2(n_4631),
.B(n_4505),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_5028),
.Y(n_5047)
);

AOI221xp5_ASAP7_75t_SL g5048 ( 
.A1(n_5034),
.A2(n_4670),
.B1(n_4699),
.B2(n_4657),
.C(n_4694),
.Y(n_5048)
);

AOI222xp33_ASAP7_75t_L g5049 ( 
.A1(n_5046),
.A2(n_4570),
.B1(n_4601),
.B2(n_4584),
.C1(n_4604),
.C2(n_4694),
.Y(n_5049)
);

AOI211x1_ASAP7_75t_SL g5050 ( 
.A1(n_5035),
.A2(n_4602),
.B(n_4596),
.C(n_4523),
.Y(n_5050)
);

NAND3xp33_ASAP7_75t_SL g5051 ( 
.A(n_5027),
.B(n_4657),
.C(n_4570),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_SL g5052 ( 
.A(n_5026),
.B(n_4705),
.Y(n_5052)
);

AOI211x1_ASAP7_75t_SL g5053 ( 
.A1(n_5023),
.A2(n_4602),
.B(n_4596),
.C(n_4523),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_5045),
.B(n_4705),
.Y(n_5054)
);

NAND3xp33_ASAP7_75t_SL g5055 ( 
.A(n_5029),
.B(n_4624),
.C(n_4505),
.Y(n_5055)
);

OAI21xp5_ASAP7_75t_L g5056 ( 
.A1(n_5031),
.A2(n_4512),
.B(n_4636),
.Y(n_5056)
);

AOI222xp33_ASAP7_75t_L g5057 ( 
.A1(n_5044),
.A2(n_4633),
.B1(n_4635),
.B2(n_4654),
.C1(n_4580),
.C2(n_4659),
.Y(n_5057)
);

OAI21xp33_ASAP7_75t_L g5058 ( 
.A1(n_5032),
.A2(n_4635),
.B(n_4659),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_5033),
.B(n_5040),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_SL g5060 ( 
.A(n_5037),
.B(n_5025),
.Y(n_5060)
);

NOR2x1_ASAP7_75t_L g5061 ( 
.A(n_5024),
.B(n_4624),
.Y(n_5061)
);

NOR2xp33_ASAP7_75t_L g5062 ( 
.A(n_5030),
.B(n_4633),
.Y(n_5062)
);

O2A1O1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_5042),
.A2(n_4600),
.B(n_4598),
.C(n_4582),
.Y(n_5063)
);

AND2x2_ASAP7_75t_L g5064 ( 
.A(n_5057),
.B(n_5036),
.Y(n_5064)
);

NOR4xp25_ASAP7_75t_SL g5065 ( 
.A(n_5060),
.B(n_5043),
.C(n_5038),
.D(n_5041),
.Y(n_5065)
);

NAND3xp33_ASAP7_75t_L g5066 ( 
.A(n_5062),
.B(n_5039),
.C(n_4633),
.Y(n_5066)
);

AOI211xp5_ASAP7_75t_L g5067 ( 
.A1(n_5058),
.A2(n_5047),
.B(n_5051),
.C(n_5059),
.Y(n_5067)
);

NOR4xp25_ASAP7_75t_L g5068 ( 
.A(n_5052),
.B(n_4549),
.C(n_4491),
.D(n_4589),
.Y(n_5068)
);

NOR4xp25_ASAP7_75t_L g5069 ( 
.A(n_5063),
.B(n_4491),
.C(n_4589),
.D(n_4592),
.Y(n_5069)
);

BUFx2_ASAP7_75t_L g5070 ( 
.A(n_5061),
.Y(n_5070)
);

NAND3xp33_ASAP7_75t_L g5071 ( 
.A(n_5054),
.B(n_4654),
.C(n_4638),
.Y(n_5071)
);

AOI211xp5_ASAP7_75t_L g5072 ( 
.A1(n_5055),
.A2(n_4591),
.B(n_4654),
.C(n_4638),
.Y(n_5072)
);

NAND4xp25_ASAP7_75t_L g5073 ( 
.A(n_5050),
.B(n_4591),
.C(n_4638),
.D(n_4559),
.Y(n_5073)
);

O2A1O1Ixp33_ASAP7_75t_L g5074 ( 
.A1(n_5056),
.A2(n_5049),
.B(n_5053),
.C(n_5048),
.Y(n_5074)
);

AOI21xp5_ASAP7_75t_L g5075 ( 
.A1(n_5060),
.A2(n_4578),
.B(n_4575),
.Y(n_5075)
);

NOR2x1_ASAP7_75t_L g5076 ( 
.A(n_5062),
.B(n_4600),
.Y(n_5076)
);

NOR3xp33_ASAP7_75t_SL g5077 ( 
.A(n_5060),
.B(n_4557),
.C(n_4528),
.Y(n_5077)
);

AND2x2_ASAP7_75t_SL g5078 ( 
.A(n_5062),
.B(n_4574),
.Y(n_5078)
);

NAND3xp33_ASAP7_75t_L g5079 ( 
.A(n_5067),
.B(n_4592),
.C(n_4590),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_5078),
.B(n_4575),
.Y(n_5080)
);

NOR3xp33_ASAP7_75t_L g5081 ( 
.A(n_5070),
.B(n_4575),
.C(n_4582),
.Y(n_5081)
);

NOR3xp33_ASAP7_75t_SL g5082 ( 
.A(n_5066),
.B(n_633),
.C(n_634),
.Y(n_5082)
);

NOR2xp33_ASAP7_75t_L g5083 ( 
.A(n_5071),
.B(n_4568),
.Y(n_5083)
);

AOI221xp5_ASAP7_75t_SL g5084 ( 
.A1(n_5075),
.A2(n_4518),
.B1(n_4542),
.B2(n_4547),
.C(n_4548),
.Y(n_5084)
);

NOR4xp25_ASAP7_75t_L g5085 ( 
.A(n_5074),
.B(n_4555),
.C(n_4558),
.D(n_4514),
.Y(n_5085)
);

NOR2x1_ASAP7_75t_L g5086 ( 
.A(n_5076),
.B(n_4502),
.Y(n_5086)
);

HB1xp67_ASAP7_75t_L g5087 ( 
.A(n_5064),
.Y(n_5087)
);

AOI21xp33_ASAP7_75t_SL g5088 ( 
.A1(n_5069),
.A2(n_636),
.B(n_637),
.Y(n_5088)
);

NOR4xp25_ASAP7_75t_L g5089 ( 
.A(n_5065),
.B(n_4526),
.C(n_4509),
.D(n_4534),
.Y(n_5089)
);

NAND4xp25_ASAP7_75t_L g5090 ( 
.A(n_5073),
.B(n_4546),
.C(n_4574),
.D(n_4579),
.Y(n_5090)
);

AOI221xp5_ASAP7_75t_L g5091 ( 
.A1(n_5068),
.A2(n_5077),
.B1(n_5072),
.B2(n_4507),
.C(n_4504),
.Y(n_5091)
);

NOR2xp33_ASAP7_75t_SL g5092 ( 
.A(n_5070),
.B(n_4473),
.Y(n_5092)
);

AND4x2_ASAP7_75t_L g5093 ( 
.A(n_5076),
.B(n_4522),
.C(n_4502),
.D(n_4487),
.Y(n_5093)
);

OAI211xp5_ASAP7_75t_SL g5094 ( 
.A1(n_5067),
.A2(n_4546),
.B(n_4481),
.C(n_4516),
.Y(n_5094)
);

NOR2x1_ASAP7_75t_L g5095 ( 
.A(n_5070),
.B(n_4566),
.Y(n_5095)
);

AOI221xp5_ASAP7_75t_L g5096 ( 
.A1(n_5069),
.A2(n_4536),
.B1(n_4574),
.B2(n_4560),
.C(n_4539),
.Y(n_5096)
);

INVx2_ASAP7_75t_SL g5097 ( 
.A(n_5080),
.Y(n_5097)
);

HB1xp67_ASAP7_75t_L g5098 ( 
.A(n_5083),
.Y(n_5098)
);

OR2x2_ASAP7_75t_L g5099 ( 
.A(n_5090),
.B(n_4537),
.Y(n_5099)
);

AOI22xp5_ASAP7_75t_L g5100 ( 
.A1(n_5092),
.A2(n_5081),
.B1(n_5079),
.B2(n_5087),
.Y(n_5100)
);

NOR2x1_ASAP7_75t_L g5101 ( 
.A(n_5094),
.B(n_4566),
.Y(n_5101)
);

AOI22xp33_ASAP7_75t_L g5102 ( 
.A1(n_5096),
.A2(n_4541),
.B1(n_4537),
.B2(n_4539),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5082),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5088),
.Y(n_5104)
);

AOI22xp33_ASAP7_75t_L g5105 ( 
.A1(n_5086),
.A2(n_4540),
.B1(n_4541),
.B2(n_4579),
.Y(n_5105)
);

OR2x2_ASAP7_75t_L g5106 ( 
.A(n_5089),
.B(n_4540),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5091),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5085),
.Y(n_5108)
);

OAI211xp5_ASAP7_75t_SL g5109 ( 
.A1(n_5084),
.A2(n_636),
.B(n_637),
.C(n_638),
.Y(n_5109)
);

AOI22xp5_ASAP7_75t_L g5110 ( 
.A1(n_5095),
.A2(n_4473),
.B1(n_4476),
.B2(n_4503),
.Y(n_5110)
);

AND2x4_ASAP7_75t_L g5111 ( 
.A(n_5093),
.B(n_4476),
.Y(n_5111)
);

AND3x4_ASAP7_75t_L g5112 ( 
.A(n_5082),
.B(n_4597),
.C(n_4587),
.Y(n_5112)
);

NOR2x1_ASAP7_75t_L g5113 ( 
.A(n_5080),
.B(n_638),
.Y(n_5113)
);

INVxp67_ASAP7_75t_SL g5114 ( 
.A(n_5113),
.Y(n_5114)
);

NOR3xp33_ASAP7_75t_SL g5115 ( 
.A(n_5104),
.B(n_639),
.C(n_640),
.Y(n_5115)
);

NAND4xp25_ASAP7_75t_L g5116 ( 
.A(n_5100),
.B(n_4594),
.C(n_4586),
.D(n_4583),
.Y(n_5116)
);

NAND3xp33_ASAP7_75t_L g5117 ( 
.A(n_5107),
.B(n_5098),
.C(n_5108),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5111),
.B(n_4478),
.Y(n_5118)
);

NOR3xp33_ASAP7_75t_L g5119 ( 
.A(n_5097),
.B(n_4561),
.C(n_4597),
.Y(n_5119)
);

OR2x6_ASAP7_75t_L g5120 ( 
.A(n_5103),
.B(n_4561),
.Y(n_5120)
);

AOI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_5109),
.A2(n_4597),
.B1(n_641),
.B2(n_642),
.C(n_643),
.Y(n_5121)
);

NOR2x1_ASAP7_75t_L g5122 ( 
.A(n_5106),
.B(n_639),
.Y(n_5122)
);

HB1xp67_ASAP7_75t_L g5123 ( 
.A(n_5099),
.Y(n_5123)
);

NOR3xp33_ASAP7_75t_L g5124 ( 
.A(n_5101),
.B(n_642),
.C(n_643),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_5118),
.B(n_5105),
.Y(n_5125)
);

AND2x2_ASAP7_75t_SL g5126 ( 
.A(n_5124),
.B(n_5102),
.Y(n_5126)
);

OAI221xp5_ASAP7_75t_SL g5127 ( 
.A1(n_5121),
.A2(n_5110),
.B1(n_5112),
.B2(n_646),
.C(n_648),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_5115),
.B(n_644),
.Y(n_5128)
);

NOR3xp33_ASAP7_75t_L g5129 ( 
.A(n_5117),
.B(n_5114),
.C(n_5123),
.Y(n_5129)
);

NAND3xp33_ASAP7_75t_SL g5130 ( 
.A(n_5122),
.B(n_644),
.C(n_645),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_5128),
.B(n_5116),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5130),
.B(n_5127),
.Y(n_5132)
);

HB1xp67_ASAP7_75t_L g5133 ( 
.A(n_5125),
.Y(n_5133)
);

OAI22xp5_ASAP7_75t_L g5134 ( 
.A1(n_5133),
.A2(n_5126),
.B1(n_5129),
.B2(n_5120),
.Y(n_5134)
);

AOI22xp5_ASAP7_75t_L g5135 ( 
.A1(n_5131),
.A2(n_5119),
.B1(n_5120),
.B2(n_649),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_5135),
.Y(n_5136)
);

AO221x1_ASAP7_75t_L g5137 ( 
.A1(n_5136),
.A2(n_5134),
.B1(n_5132),
.B2(n_649),
.C(n_650),
.Y(n_5137)
);

OA21x2_ASAP7_75t_L g5138 ( 
.A1(n_5137),
.A2(n_645),
.B(n_648),
.Y(n_5138)
);

AOI22xp33_ASAP7_75t_R g5139 ( 
.A1(n_5138),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.Y(n_5139)
);

NAND3xp33_ASAP7_75t_L g5140 ( 
.A(n_5139),
.B(n_652),
.C(n_654),
.Y(n_5140)
);

OAI22xp5_ASAP7_75t_SL g5141 ( 
.A1(n_5140),
.A2(n_654),
.B1(n_655),
.B2(n_656),
.Y(n_5141)
);

AOI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_5141),
.A2(n_655),
.B(n_656),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5142),
.Y(n_5143)
);

AOI22xp33_ASAP7_75t_L g5144 ( 
.A1(n_5143),
.A2(n_657),
.B1(n_658),
.B2(n_659),
.Y(n_5144)
);

INVx1_ASAP7_75t_SL g5145 ( 
.A(n_5144),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5144),
.Y(n_5146)
);

AOI21xp5_ASAP7_75t_L g5147 ( 
.A1(n_5145),
.A2(n_660),
.B(n_661),
.Y(n_5147)
);

OR2x6_ASAP7_75t_L g5148 ( 
.A(n_5146),
.B(n_660),
.Y(n_5148)
);

OAI221xp5_ASAP7_75t_R g5149 ( 
.A1(n_5147),
.A2(n_661),
.B1(n_662),
.B2(n_663),
.C(n_664),
.Y(n_5149)
);

AOI221xp5_ASAP7_75t_L g5150 ( 
.A1(n_5148),
.A2(n_662),
.B1(n_664),
.B2(n_666),
.C(n_667),
.Y(n_5150)
);

AOI22xp33_ASAP7_75t_L g5151 ( 
.A1(n_5149),
.A2(n_5150),
.B1(n_667),
.B2(n_668),
.Y(n_5151)
);

AOI211xp5_ASAP7_75t_L g5152 ( 
.A1(n_5151),
.A2(n_666),
.B(n_668),
.C(n_669),
.Y(n_5152)
);


endmodule