module real_jpeg_10986_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_1),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_56),
.B1(n_58),
.B2(n_69),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_16),
.B(n_56),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_42),
.B1(n_56),
.B2(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_12),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_56),
.B1(n_58),
.B2(n_74),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_74),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_13),
.A2(n_68),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_78),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_78),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_68),
.B1(n_73),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_56),
.B1(n_58),
.B2(n_95),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_95),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_95),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_16),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_16),
.A2(n_68),
.B1(n_73),
.B2(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_76),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_16),
.A2(n_40),
.B(n_44),
.C(n_176),
.D(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_16),
.B(n_40),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_63),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_16),
.A2(n_26),
.B(n_191),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_16),
.A2(n_58),
.B(n_59),
.C(n_126),
.D(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_16),
.B(n_58),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_103),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_79),
.B2(n_80),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_38),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_35),
.B(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_26),
.A2(n_33),
.B1(n_35),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_26),
.A2(n_35),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_26),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_32),
.B1(n_120),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_27),
.A2(n_32),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_27),
.B(n_192),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_28),
.B(n_45),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_28),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_29),
.A2(n_47),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_32),
.B(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_35),
.A2(n_197),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_35),
.B(n_116),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_35),
.A2(n_205),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_43),
.B1(n_51),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_40),
.B(n_60),
.Y(n_227)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_41),
.A2(n_62),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_43),
.A2(n_51),
.B1(n_188),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_43),
.A2(n_219),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_44),
.B(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_51),
.A2(n_91),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_51),
.B(n_142),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_51),
.A2(n_140),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_51),
.B(n_116),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_72),
.B(n_75),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_69),
.B(n_116),
.C(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_94),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_96),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_123),
.B1(n_124),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_99),
.A2(n_100),
.B(n_148),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_107),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_106),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_108),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_121),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_110),
.B1(n_121),
.B2(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_118),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_168),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_152),
.B(n_167),
.Y(n_131)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_149),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_146),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_153),
.B(n_155),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_156),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_158),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_162),
.A2(n_163),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_164),
.B(n_165),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_251),
.C(n_252),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_245),
.B(n_250),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_232),
.B(n_244),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_213),
.B(n_231),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_193),
.B(n_212),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_174),
.B(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_178),
.B1(n_179),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_201),
.B(n_211),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_199),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_210),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_224),
.B2(n_230),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_223),
.C(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_234),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_240),
.C(n_242),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_239),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);


endmodule