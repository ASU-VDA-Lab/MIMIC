module fake_jpeg_27104_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_57),
.Y(n_78)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_39),
.Y(n_98)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_28),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_89),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_16),
.B1(n_41),
.B2(n_19),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_105)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_16),
.B1(n_35),
.B2(n_41),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_94),
.B1(n_17),
.B2(n_23),
.Y(n_116)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_33),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_33),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_30),
.Y(n_104)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_16),
.B1(n_32),
.B2(n_31),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_21),
.B1(n_38),
.B2(n_39),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_18),
.B1(n_30),
.B2(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_95),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_76),
.B1(n_82),
.B2(n_81),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_18),
.B1(n_20),
.B2(n_30),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_114),
.B1(n_122),
.B2(n_65),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_17),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_25),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_29),
.B(n_33),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_36),
.B(n_29),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_118),
.B1(n_102),
.B2(n_106),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_137),
.B(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_136),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_73),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_92),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_77),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_155),
.B1(n_118),
.B2(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_148),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_74),
.C(n_87),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_129),
.C(n_112),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_21),
.B(n_1),
.C(n_2),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_0),
.B(n_1),
.Y(n_188)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_158),
.B1(n_63),
.B2(n_67),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_69),
.B1(n_70),
.B2(n_82),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_22),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_160),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_126),
.C(n_107),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_104),
.B(n_128),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_162),
.A2(n_179),
.B(n_183),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_126),
.CI(n_114),
.CON(n_165),
.SN(n_165)
);

OAI211xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_15),
.B(n_14),
.C(n_12),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_105),
.B1(n_116),
.B2(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_175),
.B1(n_187),
.B2(n_190),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_171),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_112),
.C(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_178),
.B1(n_22),
.B2(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_145),
.B1(n_142),
.B2(n_137),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_120),
.B(n_121),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_120),
.C(n_124),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_109),
.B(n_115),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_60),
.B1(n_118),
.B2(n_109),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_0),
.B(n_2),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_133),
.A2(n_72),
.B1(n_67),
.B2(n_21),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_141),
.C(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_156),
.B1(n_144),
.B2(n_135),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_139),
.B(n_147),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_172),
.B(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_168),
.B1(n_177),
.B2(n_186),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_136),
.B1(n_154),
.B2(n_152),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_154),
.B1(n_140),
.B2(n_148),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_217),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_134),
.B1(n_158),
.B2(n_22),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_22),
.A3(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_210),
.B(n_165),
.CI(n_14),
.CON(n_235),
.SN(n_235)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_179),
.A2(n_183),
.B1(n_182),
.B2(n_159),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_215),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_174),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_221),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_162),
.B1(n_174),
.B2(n_181),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_2),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_191),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_160),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_203),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_171),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_234),
.B(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_193),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_180),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_184),
.C(n_165),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_238),
.C(n_241),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_184),
.C(n_11),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_11),
.C(n_10),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_11),
.C(n_4),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_241),
.C(n_215),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_196),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_195),
.C(n_203),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_256),
.C(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_217),
.C(n_194),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_194),
.C(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_243),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_240),
.A2(n_228),
.B1(n_231),
.B2(n_223),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_228),
.B1(n_200),
.B2(n_216),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_272),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_232),
.B(n_240),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_216),
.B(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_238),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_256),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_212),
.B1(n_246),
.B2(n_236),
.Y(n_291)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_201),
.C(n_236),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_201),
.Y(n_282)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_199),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_207),
.B1(n_252),
.B2(n_235),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_250),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_252),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_273),
.B(n_269),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_271),
.B1(n_281),
.B2(n_269),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_274),
.B1(n_268),
.B2(n_245),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_286),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_280),
.B(n_275),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_274),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_204),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_303),
.B1(n_304),
.B2(n_302),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_286),
.C(n_293),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_268),
.B1(n_198),
.B2(n_5),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_3),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_312),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_307),
.CI(n_311),
.CON(n_319),
.SN(n_319)
);

AOI211xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_305),
.B(n_314),
.C(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_305),
.C(n_319),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.C(n_309),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_303),
.B1(n_296),
.B2(n_5),
.Y(n_323)
);


endmodule