module fake_jpeg_9446_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_42),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_67),
.B1(n_68),
.B2(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_16),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_30),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_57),
.B1(n_17),
.B2(n_27),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_44),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_42),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_18),
.B(n_16),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_73),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_92),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_83),
.B1(n_58),
.B2(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_36),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_26),
.B(n_29),
.C(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_94),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_16),
.B1(n_37),
.B2(n_42),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_42),
.B1(n_33),
.B2(n_20),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_84),
.B1(n_87),
.B2(n_44),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_33),
.B1(n_20),
.B2(n_27),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_29),
.B1(n_26),
.B2(n_17),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_95),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_36),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_93),
.B(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_97),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_51),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_49),
.B1(n_60),
.B2(n_58),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_113),
.B1(n_88),
.B2(n_89),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_40),
.Y(n_112)
);

AO21x2_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_65),
.B(n_61),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_36),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_91),
.B(n_65),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_43),
.B1(n_36),
.B2(n_51),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_89),
.B1(n_76),
.B2(n_51),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_93),
.A3(n_91),
.B1(n_74),
.B2(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_123),
.A2(n_114),
.B(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_74),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_25),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_133),
.B1(n_115),
.B2(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_79),
.B1(n_88),
.B2(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_52),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_148),
.B1(n_82),
.B2(n_62),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_89),
.B1(n_102),
.B2(n_109),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_98),
.B(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_110),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_98),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_151),
.A2(n_166),
.B(n_173),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_162),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_170),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_118),
.B1(n_105),
.B2(n_116),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_103),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_118),
.B1(n_99),
.B2(n_114),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_167),
.B1(n_171),
.B2(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_165),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_118),
.B1(n_112),
.B2(n_76),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_139),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_54),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_174),
.C(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_148),
.B1(n_138),
.B2(n_131),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_97),
.B1(n_106),
.B2(n_96),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_54),
.C(n_62),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_176),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_145),
.C(n_129),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_197),
.C(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_180),
.B(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_190),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_134),
.B(n_129),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_185),
.B(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_199),
.B1(n_190),
.B2(n_194),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_124),
.C(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_217),
.C(n_220),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_150),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_222),
.B(n_176),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_215),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_154),
.B1(n_193),
.B2(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_216),
.B(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_158),
.C(n_174),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_183),
.B1(n_179),
.B2(n_82),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_151),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_235),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_191),
.C(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_197),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_214),
.B1(n_200),
.B2(n_209),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_205),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_82),
.C(n_54),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_240),
.C(n_213),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_21),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_61),
.C(n_43),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_21),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_61),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_241),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_246),
.C(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_214),
.C(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_210),
.B1(n_222),
.B2(n_204),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_254),
.B1(n_258),
.B2(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_240),
.C(n_225),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_239),
.C(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_32),
.C(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_32),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_1),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_271),
.Y(n_281)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_242),
.C(n_2),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_224),
.B1(n_43),
.B2(n_32),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_245),
.B1(n_251),
.B2(n_257),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_253),
.B(n_21),
.Y(n_275)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_272),
.C(n_256),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_9),
.C(n_3),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_280),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_256),
.B(n_21),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_272),
.B(n_267),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_9),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_265),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_264),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_291),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_261),
.A3(n_270),
.B1(n_7),
.B2(n_8),
.C1(n_12),
.C2(n_13),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_5),
.C(n_8),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_299),
.B(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_276),
.B(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_300),
.B(n_13),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_284),
.B(n_21),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_8),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_305),
.B(n_306),
.Y(n_307)
);

OAI211xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_14),
.B(n_15),
.C(n_1),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_14),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_308),
.B(n_304),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_15),
.Y(n_311)
);


endmodule