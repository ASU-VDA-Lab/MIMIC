module fake_jpeg_18690_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_23),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_29),
.B1(n_28),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_37),
.B1(n_28),
.B2(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_59),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_72),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_34),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_74),
.B1(n_76),
.B2(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_32),
.B1(n_21),
.B2(n_27),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_71),
.B1(n_84),
.B2(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_21),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_41),
.B1(n_36),
.B2(n_27),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_38),
.B(n_39),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_39),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_94),
.B1(n_98),
.B2(n_69),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_38),
.B1(n_25),
.B2(n_22),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_23),
.C(n_22),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_20),
.C(n_18),
.Y(n_127)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_20),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_17),
.B(n_1),
.C(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_0),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_115),
.B(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_125),
.Y(n_135)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_128),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_84),
.B(n_83),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_77),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_119),
.B(n_103),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_86),
.B1(n_99),
.B2(n_106),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_123),
.B1(n_92),
.B2(n_93),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_82),
.B(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_67),
.B1(n_63),
.B2(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_130),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_89),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_20),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_64),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_5),
.B(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_58),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_58),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_79),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_143),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_109),
.B1(n_93),
.B2(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_149),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_150),
.B(n_122),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_111),
.B1(n_130),
.B2(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_149),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_93),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_63),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_132),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_104),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_108),
.C(n_30),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_126),
.C(n_113),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_5),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_166),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_118),
.B(n_133),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_173),
.B(n_174),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_148),
.C(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_117),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_175),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_190),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_147),
.B1(n_154),
.B2(n_141),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_167),
.B1(n_158),
.B2(n_161),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_163),
.C(n_165),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_140),
.B(n_151),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_180),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_180),
.C(n_184),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_6),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_179),
.A2(n_167),
.B1(n_173),
.B2(n_166),
.Y(n_198)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_114),
.B1(n_178),
.B2(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_162),
.B1(n_155),
.B2(n_165),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_210),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_189),
.B(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_190),
.C(n_178),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_201),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_17),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_198),
.B1(n_210),
.B2(n_11),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_208),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_211),
.B(n_10),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_199),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_8),
.B(n_10),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_217),
.A3(n_220),
.B1(n_218),
.B2(n_16),
.C1(n_24),
.C2(n_30),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_12),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C1(n_24),
.C2(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_16),
.C(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_15),
.Y(n_230)
);


endmodule