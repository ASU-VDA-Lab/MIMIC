module real_jpeg_24756_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_64),
.C(n_86),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_78),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_58),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_4),
.A2(n_102),
.B1(n_171),
.B2(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_98),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_7),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_45),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_8),
.A2(n_45),
.B1(n_63),
.B2(n_64),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_8),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_28),
.C(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_11),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_75),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_19),
.B(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_81),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_20),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_59),
.B2(n_80),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_42),
.C(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_25),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_40),
.B1(n_98),
.B2(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_30),
.B(n_77),
.C(n_79),
.Y(n_76)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_30),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_29),
.B(n_49),
.C(n_53),
.Y(n_189)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_30),
.B(n_78),
.CON(n_188),
.SN(n_188)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_36),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_38),
.B(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_55),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_46),
.A2(n_51),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_56),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_47),
.A2(n_58),
.B1(n_188),
.B2(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_50),
.A2(n_52),
.B(n_187),
.C(n_189),
.Y(n_186)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_132),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_53),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_76),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_60),
.A2(n_61),
.B1(n_76),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_70),
.B2(n_74),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_62),
.B(n_105),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_62),
.A2(n_70),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_64),
.B1(n_86),
.B2(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_63),
.B(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_68),
.A2(n_73),
.B(n_119),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_71),
.A2(n_102),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_76),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_78),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_78),
.B(n_88),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_78),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_81),
.B(n_100),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_93),
.C(n_95),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_82),
.B(n_93),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B(n_90),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_122),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_83),
.A2(n_122),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_84),
.A2(n_88),
.B1(n_150),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_84),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_89),
.B(n_122),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_95),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_115),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_102),
.A2(n_104),
.B(n_118),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_133),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_125),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_120),
.B2(n_124),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_236),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_232),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_222),
.B(n_231),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_200),
.B(n_221),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_182),
.B(n_199),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_160),
.B(n_181),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_180),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_166),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_172),
.B(n_179),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_198),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_198),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_193),
.C(n_195),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_213),
.B2(n_214),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_216),
.C(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_209),
.C(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_230),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_227),
.C(n_228),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);


endmodule