module real_jpeg_12576_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_296, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_296;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_288;
wire n_292;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_131;
wire n_47;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_167;
wire n_213;
wire n_179;
wire n_128;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_31),
.B1(n_35),
.B2(n_98),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_6),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_6),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_31),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_41),
.B1(n_55),
.B2(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_26),
.B1(n_49),
.B2(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_10),
.A2(n_26),
.B1(n_31),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_10),
.A2(n_26),
.B1(n_55),
.B2(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_10),
.B(n_67),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_22),
.C(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_10),
.B(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_10),
.B(n_36),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_56),
.B(n_69),
.C(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_54),
.Y(n_191)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_275),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_119),
.B(n_273),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_16),
.B(n_99),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_59),
.C(n_76),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_17),
.A2(n_18),
.B1(n_59),
.B2(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_42),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_19),
.A2(n_20),
.B(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_20),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_20),
.A2(n_43),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_20),
.B(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_20),
.A2(n_27),
.B1(n_43),
.B2(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_25),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_21),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_21),
.B(n_25),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_21),
.A2(n_208),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

AO22x1_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_22),
.B(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_24),
.B(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_83),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_24),
.A2(n_82),
.B(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_26),
.A2(n_35),
.B(n_70),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_26),
.B(n_52),
.C(n_56),
.Y(n_206)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_37),
.B(n_39),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_28),
.A2(n_64),
.B(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_29),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_29),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_29),
.B(n_63),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_31),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_31),
.B(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_36),
.B(n_136),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_61),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_39),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_39),
.B(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_57),
.B(n_58),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_47),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_47),
.B(n_107),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_50),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_54),
.B(n_97),
.Y(n_214)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_57),
.A2(n_236),
.B(n_286),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_59),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_75),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_65),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_62),
.B(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_71),
.Y(n_65)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_67),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_67),
.B(n_91),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_67),
.A2(n_90),
.B(n_91),
.Y(n_237)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_74),
.Y(n_87)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_71),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_71),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_72),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_102),
.B1(n_103),
.B2(n_118),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_75),
.B(n_100),
.C(n_102),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_76),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.C(n_92),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_77),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_78),
.B(n_84),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_82),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_86),
.A2(n_92),
.B1(n_93),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_87),
.B(n_193),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_89),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_96),
.B(n_106),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_104),
.B(n_113),
.C(n_114),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_104),
.A2(n_105),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_112),
.A2(n_113),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_112),
.B(n_212),
.C(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_112),
.A2(n_113),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_267),
.B(n_272),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_254),
.B(n_266),
.Y(n_120)
);

AOI321xp33_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_220),
.A3(n_247),
.B1(n_252),
.B2(n_253),
.C(n_296),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_198),
.B(n_219),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_181),
.B(n_197),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_168),
.B(n_180),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_148),
.B(n_167),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_141),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_141),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_140),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_138),
.C(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_161),
.B(n_166),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_156),
.B(n_160),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_159),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_170),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_196),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_196),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B1(n_189),
.B2(n_195),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_203),
.C(n_210),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.CI(n_192),
.CON(n_189),
.SN(n_189)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_210),
.B2(n_211),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_209),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_241),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_241),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_229),
.C(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_227),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_225),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_256),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_263),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_293),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_287),
.B1(n_288),
.B2(n_292),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);


endmodule