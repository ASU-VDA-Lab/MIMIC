module fake_jpeg_8768_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx6_ASAP7_75t_SL g7 ( 
.A(n_3),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_2),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_13),
.B1(n_9),
.B2(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_25),
.B1(n_8),
.B2(n_18),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_6),
.B1(n_9),
.B2(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_14),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_22),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_11),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_22),
.C(n_19),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_27),
.B(n_11),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_27),
.B(n_19),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_34),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_28),
.Y(n_35)
);

AOI21x1_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_10),
.B(n_17),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_10),
.C(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_10),
.B1(n_4),
.B2(n_3),
.C(n_17),
.Y(n_40)
);


endmodule