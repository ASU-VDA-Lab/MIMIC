module fake_jpeg_15136_n_263 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_1),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_19),
.B1(n_30),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_50),
.B1(n_64),
.B2(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_19),
.B1(n_30),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_26),
.B1(n_17),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_19),
.B1(n_30),
.B2(n_20),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_33),
.B1(n_23),
.B2(n_32),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_37),
.B1(n_33),
.B2(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_66),
.A2(n_76),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_37),
.C(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_71),
.C(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_84),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_36),
.C(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_79),
.B1(n_88),
.B2(n_24),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_18),
.B(n_25),
.C(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_8),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_26),
.B1(n_36),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_86),
.B1(n_22),
.B2(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_78),
.B(n_91),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_80),
.Y(n_121)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_24),
.B1(n_22),
.B2(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_37),
.B1(n_41),
.B2(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_32),
.Y(n_89)
);

OR2x4_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_37),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_27),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_21),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_3),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_41),
.B(n_21),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_109),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_115),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_51),
.B1(n_41),
.B2(n_23),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_127),
.B1(n_125),
.B2(n_128),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_126),
.B(n_10),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_4),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_11),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_8),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_9),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_155),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_71),
.C(n_69),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_110),
.C(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_156),
.B1(n_127),
.B2(n_122),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_66),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_102),
.C(n_77),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_143),
.Y(n_164)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_98),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_110),
.B(n_12),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_88),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_150),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_72),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_100),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_10),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_126),
.B(n_114),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_105),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_141),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_176),
.B1(n_180),
.B2(n_179),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_165),
.B(n_174),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_178),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_106),
.B(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_143),
.B1(n_81),
.B2(n_82),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_145),
.B1(n_154),
.B2(n_151),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_181),
.C(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_147),
.Y(n_185)
);

AO32x1_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_146),
.A3(n_153),
.B1(n_147),
.B2(n_149),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_192),
.B(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_190),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_195),
.B1(n_163),
.B2(n_161),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_189),
.C(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_138),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_144),
.B(n_137),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_195),
.B(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_132),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_134),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_75),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_199),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_95),
.B1(n_121),
.B2(n_101),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_164),
.B1(n_178),
.B2(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_172),
.B(n_11),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_67),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_160),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_162),
.C(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.C(n_215),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_166),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_177),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_191),
.B(n_185),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_161),
.C(n_99),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_200),
.B1(n_81),
.B2(n_83),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_229),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_193),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_194),
.B(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_208),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_200),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_215),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_236),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_205),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_237),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_224),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_246),
.B(n_220),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_216),
.B(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_252),
.C(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_235),
.Y(n_252)
);

OAI321xp33_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_236),
.A3(n_202),
.B1(n_229),
.B2(n_232),
.C(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_212),
.B1(n_225),
.B2(n_67),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_225),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_12),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_256),
.C2(n_257),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_121),
.B1(n_99),
.B2(n_15),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.C(n_12),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_14),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);


endmodule