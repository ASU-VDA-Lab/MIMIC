module fake_jpeg_5084_n_39 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_19),
.B(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_0),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.C(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_1),
.C(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_10),
.B1(n_17),
.B2(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_20),
.B1(n_12),
.B2(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_22),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_24),
.B(n_22),
.C(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_27),
.B1(n_13),
.B2(n_5),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_25),
.B1(n_6),
.B2(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_3),
.B1(n_4),
.B2(n_29),
.Y(n_39)
);


endmodule