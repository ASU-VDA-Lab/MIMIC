module fake_jpeg_3079_n_468 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_468);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_468;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_50),
.B(n_72),
.Y(n_158)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_6),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_75),
.Y(n_160)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_SL g78 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_90),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_15),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_97),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_15),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_18),
.B(n_5),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_34),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_105),
.A2(n_107),
.B1(n_134),
.B2(n_148),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_117),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_76),
.B1(n_61),
.B2(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_110),
.B(n_142),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_47),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_44),
.B1(n_23),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_44),
.B1(n_45),
.B2(n_42),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_73),
.B(n_23),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_36),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_44),
.B1(n_22),
.B2(n_43),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_48),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_154),
.B1(n_27),
.B2(n_37),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_20),
.B1(n_36),
.B2(n_28),
.Y(n_154)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_168),
.Y(n_210)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_171),
.B(n_173),
.Y(n_237)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_86),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_SL g174 ( 
.A(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_175),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_179),
.Y(n_231)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_38),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_196),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_42),
.B1(n_14),
.B2(n_41),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_192),
.Y(n_234)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_108),
.B(n_81),
.C(n_95),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_133),
.C(n_160),
.Y(n_218)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_195),
.Y(n_212)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_79),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_194),
.A2(n_201),
.B1(n_27),
.B2(n_37),
.Y(n_236)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_28),
.Y(n_196)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_200),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_113),
.A2(n_14),
.B1(n_41),
.B2(n_39),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_214)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_112),
.B(n_38),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_115),
.B(n_39),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_27),
.Y(n_230)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

NOR2x1p5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_107),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_235),
.B(n_230),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_160),
.Y(n_252)
);

NAND2x1_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_130),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_242),
.B1(n_194),
.B2(n_204),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_167),
.A2(n_157),
.B(n_123),
.C(n_146),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_235),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_170),
.A2(n_105),
.B1(n_134),
.B2(n_119),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_246),
.B1(n_250),
.B2(n_262),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_197),
.B(n_206),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_188),
.C(n_166),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_208),
.B1(n_242),
.B2(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_165),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_254),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_255),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_201),
.B1(n_150),
.B2(n_157),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_187),
.B1(n_178),
.B2(n_161),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_260),
.B1(n_265),
.B2(n_213),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_266),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_214),
.B(n_234),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_264),
.Y(n_276)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_258),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_209),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_184),
.B1(n_195),
.B2(n_207),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_119),
.B1(n_190),
.B2(n_137),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_SL g264 ( 
.A(n_221),
.B(n_198),
.C(n_176),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_189),
.B1(n_164),
.B2(n_172),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_223),
.A2(n_109),
.B1(n_200),
.B2(n_202),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_133),
.B1(n_229),
.B2(n_224),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_220),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_211),
.B1(n_152),
.B2(n_224),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_205),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_222),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_217),
.B1(n_225),
.B2(n_210),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_280),
.B1(n_284),
.B2(n_295),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_244),
.A2(n_191),
.B1(n_169),
.B2(n_216),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_291),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_216),
.B1(n_219),
.B2(n_144),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_246),
.A2(n_219),
.B1(n_228),
.B2(n_227),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_265),
.B1(n_269),
.B2(n_251),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_212),
.B(n_220),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_238),
.B(n_258),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_233),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_248),
.B(n_211),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_249),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_257),
.A2(n_138),
.B1(n_141),
.B2(n_144),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_249),
.A2(n_152),
.B1(n_65),
.B2(n_80),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_262),
.B1(n_270),
.B2(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_247),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_298),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_308),
.B1(n_311),
.B2(n_277),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_304),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_302),
.A2(n_274),
.B1(n_297),
.B2(n_279),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_273),
.B(n_278),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_303),
.B(n_320),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_245),
.C(n_249),
.Y(n_304)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_307),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_260),
.B1(n_256),
.B2(n_255),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_278),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_312),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_250),
.B1(n_245),
.B2(n_271),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_252),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_264),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_266),
.C(n_127),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_316),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_155),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_238),
.C(n_116),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_287),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_276),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_267),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_287),
.B(n_290),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_279),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_274),
.Y(n_339)
);

OA22x2_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_272),
.B1(n_286),
.B2(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_342),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_280),
.B1(n_289),
.B2(n_311),
.Y(n_325)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_338),
.Y(n_361)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

AOI21xp33_ASAP7_75t_L g351 ( 
.A1(n_330),
.A2(n_306),
.B(n_313),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_332),
.A2(n_345),
.B1(n_306),
.B2(n_284),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_335),
.A2(n_122),
.B1(n_153),
.B2(n_163),
.Y(n_366)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_283),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_340),
.B(n_347),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_341),
.A2(n_109),
.B(n_58),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_282),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_300),
.A2(n_285),
.B1(n_295),
.B2(n_267),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_315),
.C(n_317),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_258),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_353),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_351),
.A2(n_336),
.B(n_342),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_308),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_331),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_360),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_359),
.B1(n_362),
.B2(n_363),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_338),
.C(n_326),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_336),
.C(n_324),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_301),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_323),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_348),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_300),
.B1(n_302),
.B2(n_285),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_296),
.B1(n_285),
.B2(n_59),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_332),
.B1(n_343),
.B2(n_365),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_83),
.B1(n_85),
.B2(n_84),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_345),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_380),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_355),
.B1(n_370),
.B2(n_364),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_376),
.A2(n_325),
.B1(n_324),
.B2(n_365),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_330),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_377),
.B(n_384),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_368),
.A2(n_341),
.B(n_325),
.C(n_337),
.Y(n_378)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_387),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_327),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_327),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_390),
.Y(n_408)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_371),
.B(n_389),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_325),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_392),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_352),
.B(n_325),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_401),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_14),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_374),
.C(n_380),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_399),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_364),
.C(n_370),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_371),
.B(n_383),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_403),
.A2(n_37),
.B1(n_5),
.B2(n_10),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_404),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_360),
.C(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_406),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_356),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_376),
.A2(n_363),
.B1(n_372),
.B2(n_324),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_11),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_369),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_410),
.B(n_375),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_394),
.A2(n_386),
.B(n_378),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_409),
.B(n_393),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_412),
.B(n_414),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_74),
.C(n_62),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_60),
.C(n_38),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_402),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_159),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_419),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_418),
.A2(n_420),
.B1(n_404),
.B2(n_405),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_11),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_401),
.B(n_13),
.CI(n_10),
.CON(n_420),
.SN(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_395),
.A2(n_100),
.B1(n_90),
.B2(n_39),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_424),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_407),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_429),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_399),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_433),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_400),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_416),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_400),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_434),
.A2(n_430),
.B(n_418),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_398),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_435),
.B(n_436),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_4),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_4),
.B(n_5),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_438),
.A2(n_420),
.B(n_422),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_446),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_414),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_445),
.B(n_437),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_413),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g452 ( 
.A1(n_444),
.A2(n_420),
.B(n_437),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_419),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_417),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_447),
.B(n_434),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_9),
.Y(n_454)
);

AO21x1_ASAP7_75t_L g457 ( 
.A1(n_450),
.A2(n_451),
.B(n_454),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_452),
.A2(n_456),
.B(n_40),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_40),
.B(n_9),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_455),
.A2(n_449),
.B(n_440),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_458),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_449),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_459),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_0),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_0),
.C(n_1),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_464),
.A2(n_465),
.B(n_463),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_457),
.C(n_40),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_466),
.A2(n_2),
.B(n_459),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_2),
.Y(n_468)
);


endmodule