module fake_jpeg_30819_n_85 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_42),
.B1(n_33),
.B2(n_35),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_35),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_34),
.B(n_30),
.C(n_32),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_4),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_6),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_4),
.B(n_5),
.Y(n_54)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_50),
.B(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_58),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_63),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_15),
.C(n_10),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_17),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND4xp25_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_72),
.C(n_62),
.D(n_48),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_13),
.C(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_16),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_27),
.C(n_68),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_66),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_74),
.B(n_77),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_78),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_65),
.B(n_67),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g85 ( 
.A(n_84),
.Y(n_85)
);


endmodule