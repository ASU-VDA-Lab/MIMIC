module fake_jpeg_15014_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_0),
.Y(n_86)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_65),
.B1(n_46),
.B2(n_49),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_92),
.B1(n_60),
.B2(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_3),
.Y(n_111)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_55),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_54),
.B1(n_63),
.B2(n_61),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_94)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_63),
.B1(n_54),
.B2(n_57),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_10),
.B1(n_14),
.B2(n_16),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_2),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_60),
.B1(n_50),
.B2(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_107),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_115),
.B1(n_117),
.B2(n_20),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_79),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_113),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_6),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_132)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_97),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_53),
.B1(n_52),
.B2(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_9),
.B1(n_10),
.B2(n_47),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_132),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_139),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_134),
.A2(n_120),
.B1(n_118),
.B2(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_112),
.B(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_97),
.C(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_133),
.C(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_119),
.B1(n_126),
.B2(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_119),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.Y(n_152)
);

AND2x4_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_138),
.B1(n_131),
.B2(n_122),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_152),
.C(n_153),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_151),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_155),
.B(n_27),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_26),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_124),
.C(n_101),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_28),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_29),
.B(n_31),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_102),
.C(n_35),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_33),
.B(n_36),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_105),
.C(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_173)
);


endmodule