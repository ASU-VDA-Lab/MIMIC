module real_jpeg_4948_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_1),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_1),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_1),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_110),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_1),
.B(n_372),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_2),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_2),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_2),
.B(n_325),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_3),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_3),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_3),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_3),
.B(n_232),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_3),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_3),
.B(n_62),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_3),
.B(n_123),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_5),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_5),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_5),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_6),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_6),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_6),
.B(n_232),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_6),
.B(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_8),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_9),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_9),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_66),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_10),
.Y(n_356)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_12),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_45),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_12),
.B(n_112),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_12),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_12),
.B(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_13),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_14),
.B(n_77),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_14),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_14),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_14),
.B(n_144),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_14),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_15),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_15),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_15),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_15),
.B(n_123),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_15),
.B(n_341),
.Y(n_340)
);

AND2x6_ASAP7_75t_SL g355 ( 
.A(n_15),
.B(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_16),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_17),
.B(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_200),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_199),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_156),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_22),
.B(n_156),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_22),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_101),
.CI(n_134),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_69),
.C(n_84),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_24),
.A2(n_25),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.C(n_52),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_26),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_33),
.C(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_33),
.B(n_104),
.C(n_109),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_33),
.A2(n_40),
.B1(n_109),
.B2(n_130),
.Y(n_155)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_35),
.Y(n_264)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_36),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_36),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_36),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_37),
.A2(n_41),
.B1(n_48),
.B2(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_39),
.Y(n_194)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_39),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_43),
.C(n_48),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_42),
.B(n_52),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_44),
.B(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_48),
.Y(n_183)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_54),
.B(n_59),
.C(n_65),
.Y(n_153)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_58),
.Y(n_180)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_63),
.Y(n_247)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_64),
.Y(n_295)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_68),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_84),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_74),
.C(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_78),
.B1(n_79),
.B2(n_83),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_78),
.A2(n_79),
.B1(n_98),
.B2(n_99),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_85),
.C(n_98),
.Y(n_84)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_82),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_82),
.Y(n_251)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_82),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_86),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.C(n_94),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_94),
.Y(n_166)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_90),
.B(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_124),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_113),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_149),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_148),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_143),
.B(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_154),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_163),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_184),
.C(n_186),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_181),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_165),
.B(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_167),
.A2(n_168),
.B1(n_181),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_177),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_169),
.B(n_177),
.Y(n_416)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_172),
.B(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_176),
.Y(n_308)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_181),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.C(n_196),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_193),
.Y(n_217)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_252),
.B(n_440),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_203),
.B(n_205),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_212),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_207),
.B(n_210),
.Y(n_436)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_212),
.B(n_436),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_236),
.C(n_239),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_214),
.B(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_226),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_215),
.A2(n_216),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_218),
.A2(n_219),
.B(n_221),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_218),
.B(n_226),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_234),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_384)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_234),
.B(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_324),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_239),
.Y(n_430)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_241),
.B(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_242),
.B(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_244),
.Y(n_397)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_248),
.B(n_249),
.Y(n_418)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_434),
.B(n_439),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_421),
.B(n_433),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_403),
.B(n_420),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_377),
.B(n_402),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_346),
.B(n_376),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_316),
.B(n_345),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_297),
.B(n_315),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_277),
.B(n_296),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_271),
.B(n_276),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_268),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.Y(n_278)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_279),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_288),
.C(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_314),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_314),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_303),
.C(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_302),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_335),
.C(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_319),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_333),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_334),
.C(n_337),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_323),
.C(n_326),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_329),
.B1(n_330),
.B2(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_342),
.C(n_343),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_340),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_342),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_375),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_375),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_359),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_358),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_358),
.C(n_401),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_357),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_355),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_391),
.C(n_392),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_366),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_368),
.C(n_373),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_363),
.C(n_364),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_373),
.B2(n_374),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_400),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_400),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_389),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_381),
.C(n_389),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_412),
.C(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_394),
.C(n_399),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_399),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_419),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_419),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_410),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_409),
.C(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_410),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_414),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_415),
.C(n_417),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_431),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_431),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_428),
.C(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_437),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_437),
.Y(n_439)
);


endmodule