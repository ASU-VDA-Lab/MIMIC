module fake_jpeg_14270_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx12f_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_23),
.Y(n_42)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_26),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_21),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_18),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_37),
.B1(n_24),
.B2(n_16),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_59),
.B1(n_46),
.B2(n_33),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_52),
.C(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_33),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_83),
.B(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_41),
.B1(n_45),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_59),
.B1(n_74),
.B2(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_63),
.B(n_33),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_2),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_57),
.B(n_60),
.C(n_65),
.D(n_13),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_33),
.B(n_20),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_53),
.B1(n_55),
.B2(n_64),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_13),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.C(n_96),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_63),
.C(n_67),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_79),
.B1(n_73),
.B2(n_71),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_18),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_79),
.B1(n_73),
.B2(n_82),
.C(n_6),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AO221x1_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_10),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_70),
.C(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_11),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_93),
.C(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_109),
.C(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_95),
.C(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_100),
.B1(n_99),
.B2(n_105),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_94),
.B1(n_89),
.B2(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_92),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_112),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_116),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_117),
.C(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_118),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_115),
.Y(n_128)
);

AOI31xp67_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_123),
.A3(n_4),
.B(n_5),
.Y(n_130)
);

OAI33xp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_128),
.A3(n_4),
.B1(n_3),
.B2(n_27),
.B3(n_13),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.Y(n_132)
);


endmodule