module fake_aes_10897_n_916 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_916);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_916;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_703;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g257 ( .A(n_161), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_89), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_137), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_251), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_189), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_74), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_172), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_250), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_224), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_76), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_43), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_184), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_168), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_21), .B(n_177), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_148), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_246), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_65), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_193), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_6), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_222), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_32), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_195), .B(n_206), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_145), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_121), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_51), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_2), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_219), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_124), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
BUFx2_ASAP7_75t_SL g288 ( .A(n_163), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_223), .Y(n_289) );
CKINVDCx14_ASAP7_75t_R g290 ( .A(n_55), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_255), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_6), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_95), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_160), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_185), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_111), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_125), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_60), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_92), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_210), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_227), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_256), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_8), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_201), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_105), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_233), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_180), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_169), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_247), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_213), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_133), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_38), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_229), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_166), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_248), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_178), .B(n_209), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_152), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_91), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_118), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_25), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_80), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_183), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_31), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_164), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_112), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_26), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_2), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_47), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_36), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_159), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_216), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_174), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_20), .Y(n_333) );
NOR2xp67_ASAP7_75t_L g334 ( .A(n_179), .B(n_167), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_241), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_103), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_249), .Y(n_337) );
CKINVDCx14_ASAP7_75t_R g338 ( .A(n_203), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_41), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_83), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_186), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_215), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_66), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_32), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_142), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_139), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_205), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_94), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_97), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_132), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_64), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_155), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_204), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_114), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_140), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_98), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_115), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_221), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_153), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_78), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_106), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_110), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_22), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_12), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_99), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_35), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_68), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_130), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_107), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_36), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_81), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_101), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_129), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_24), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_239), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_100), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_4), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_113), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_156), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_34), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_194), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_244), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_217), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_143), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_119), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_238), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_240), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_38), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_104), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_23), .Y(n_391) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_176), .B(n_181), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_225), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_109), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_120), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_182), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_207), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_9), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_9), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_50), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_131), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_56), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_108), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_87), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_88), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_245), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_307), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_271), .A2(n_45), .B(n_44), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_271), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_381), .B(n_0), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_353), .B(n_0), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_275), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_354), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_306), .B(n_1), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_296), .B(n_1), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_275), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_354), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_391), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_357), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_354), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_354), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_261), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g424 ( .A1(n_323), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_293), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_332), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_339), .A2(n_8), .B1(n_5), .B2(n_7), .Y(n_427) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_345), .B(n_46), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_387), .B(n_7), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_332), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_378), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_364), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_422), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_413), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_413), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_407), .B(n_263), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_413), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_419), .B(n_326), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_433), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
CKINVDCx6p67_ASAP7_75t_R g443 ( .A(n_432), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_433), .B(n_290), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_411), .A2(n_309), .B1(n_277), .B2(n_279), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_414), .B(n_290), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_430), .B(n_335), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_417), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AOI21x1_ASAP7_75t_L g452 ( .A1(n_408), .A2(n_348), .B(n_335), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_415), .Y(n_454) );
NAND2xp33_ASAP7_75t_SL g455 ( .A(n_410), .B(n_309), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g456 ( .A1(n_445), .A2(n_427), .B1(n_284), .B2(n_292), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_454), .B(n_418), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_452), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_441), .B(n_338), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_435), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_450), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_444), .B(n_262), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_446), .B(n_265), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_440), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_442), .B(n_428), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_453), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_447), .B(n_257), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_447), .B(n_258), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_451), .Y(n_470) );
BUFx6f_ASAP7_75t_SL g471 ( .A(n_443), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_455), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_455), .A2(n_424), .B1(n_371), .B2(n_375), .C(n_367), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_438), .A2(n_431), .B(n_416), .Y(n_474) );
INVxp33_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_434), .Y(n_476) );
BUFx6f_ASAP7_75t_SL g477 ( .A(n_437), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
NAND2xp33_ASAP7_75t_L g479 ( .A(n_437), .B(n_280), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_437), .B(n_259), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_437), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_436), .A2(n_294), .B1(n_300), .B2(n_286), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_439), .A2(n_412), .B1(n_423), .B2(n_416), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_449), .B(n_260), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_448), .B(n_266), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_449), .B(n_303), .Y(n_490) );
NAND3xp33_ASAP7_75t_SL g491 ( .A(n_449), .B(n_330), .C(n_389), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
AOI21x1_ASAP7_75t_L g493 ( .A1(n_459), .A2(n_392), .B(n_334), .Y(n_493) );
CKINVDCx10_ASAP7_75t_R g494 ( .A(n_471), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_457), .B(n_312), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_470), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_470), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_459), .A2(n_376), .B(n_344), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_492), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_460), .A2(n_270), .B(n_264), .Y(n_500) );
AOI21x1_ASAP7_75t_L g501 ( .A1(n_481), .A2(n_425), .B(n_423), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_475), .B(n_398), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_490), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_468), .A2(n_469), .B(n_463), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_472), .A2(n_425), .B1(n_431), .B2(n_426), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_468), .A2(n_281), .B(n_274), .Y(n_506) );
AO21x1_ASAP7_75t_L g507 ( .A1(n_466), .A2(n_285), .B(n_283), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_465), .B(n_399), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_469), .A2(n_479), .B(n_464), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_462), .A2(n_291), .B(n_287), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_462), .A2(n_302), .B(n_301), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_458), .B(n_365), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_467), .A2(n_313), .B(n_305), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_488), .A2(n_325), .B(n_322), .Y(n_516) );
INVx11_ASAP7_75t_L g517 ( .A(n_471), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_474), .B(n_320), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_456), .B(n_267), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_481), .A2(n_331), .B(n_328), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_466), .B(n_272), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_483), .B(n_269), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_486), .A2(n_341), .B(n_340), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_485), .A2(n_426), .B1(n_316), .B2(n_355), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_486), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_482), .A2(n_358), .B(n_351), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_476), .A2(n_360), .B(n_359), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_473), .B(n_327), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_480), .A2(n_366), .B(n_362), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_477), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_484), .B(n_370), .C(n_369), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_491), .B(n_329), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_500), .A2(n_510), .B(n_504), .C(n_509), .Y(n_535) );
AO21x1_ASAP7_75t_L g536 ( .A1(n_493), .A2(n_379), .B(n_374), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_498), .A2(n_487), .B(n_478), .Y(n_537) );
OAI21x1_ASAP7_75t_L g538 ( .A1(n_501), .A2(n_489), .B(n_487), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_528), .A2(n_352), .B(n_348), .Y(n_539) );
INVx3_ASAP7_75t_SL g540 ( .A(n_494), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_516), .A2(n_388), .B(n_395), .C(n_383), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_511), .A2(n_401), .B(n_402), .C(n_396), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_499), .B(n_333), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_522), .A2(n_406), .B(n_403), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_496), .A2(n_268), .B(n_352), .Y(n_545) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_528), .A2(n_372), .B(n_363), .Y(n_546) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_507), .A2(n_372), .B(n_363), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_497), .A2(n_380), .B(n_373), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_534), .A2(n_380), .B(n_382), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_503), .B(n_261), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_517), .Y(n_551) );
AO21x1_ASAP7_75t_L g552 ( .A1(n_525), .A2(n_288), .B(n_417), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_518), .A2(n_346), .B(n_276), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_514), .A2(n_346), .B(n_377), .C(n_417), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_513), .B(n_273), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_10), .Y(n_557) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_525), .A2(n_420), .A3(n_429), .B(n_421), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_533), .B(n_278), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_529), .B(n_282), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_531), .Y(n_561) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
AOI21xp33_ASAP7_75t_L g564 ( .A1(n_495), .A2(n_295), .B(n_289), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_519), .Y(n_565) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_512), .A2(n_377), .B(n_49), .Y(n_566) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_505), .A2(n_377), .B(n_420), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_512), .A2(n_298), .B(n_297), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_505), .A2(n_52), .B(n_48), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_527), .A2(n_524), .B(n_520), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_506), .A2(n_304), .B(n_299), .Y(n_571) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_530), .A2(n_421), .A3(n_429), .B(n_420), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_521), .Y(n_573) );
AO21x1_ASAP7_75t_L g574 ( .A1(n_523), .A2(n_421), .B(n_420), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_532), .Y(n_575) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_532), .A2(n_54), .B(n_53), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_504), .A2(n_310), .B(n_308), .Y(n_577) );
AND3x1_ASAP7_75t_SL g578 ( .A(n_494), .B(n_11), .C(n_12), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_508), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_499), .B(n_13), .Y(n_580) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_538), .A2(n_429), .B(n_421), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_561), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_580), .B(n_13), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_535), .A2(n_429), .B(n_314), .Y(n_584) );
AND2x4_ASAP7_75t_SL g585 ( .A(n_580), .B(n_14), .Y(n_585) );
OA21x2_ASAP7_75t_L g586 ( .A1(n_539), .A2(n_315), .B(n_311), .Y(n_586) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_546), .A2(n_566), .B(n_567), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_561), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_563), .B(n_14), .Y(n_590) );
OR2x6_ASAP7_75t_L g591 ( .A(n_540), .B(n_15), .Y(n_591) );
AO31x2_ASAP7_75t_L g592 ( .A1(n_552), .A2(n_18), .A3(n_16), .B(n_17), .Y(n_592) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
BUFx3_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_570), .A2(n_318), .B(n_317), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_565), .B(n_17), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_558), .Y(n_598) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_547), .A2(n_576), .B(n_537), .Y(n_599) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_555), .A2(n_321), .B(n_319), .Y(n_600) );
BUFx24_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
AO21x2_ASAP7_75t_L g602 ( .A1(n_544), .A2(n_536), .B(n_574), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
OAI21x1_ASAP7_75t_L g604 ( .A1(n_548), .A2(n_58), .B(n_57), .Y(n_604) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_542), .A2(n_336), .B(n_324), .Y(n_605) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_545), .A2(n_61), .B(n_59), .Y(n_606) );
OAI21x1_ASAP7_75t_L g607 ( .A1(n_554), .A2(n_63), .B(n_62), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_562), .B(n_337), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_541), .A2(n_343), .B(n_342), .Y(n_609) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_564), .A2(n_349), .B(n_350), .C(n_347), .Y(n_610) );
AO21x2_ASAP7_75t_L g611 ( .A1(n_549), .A2(n_69), .B(n_67), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_573), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_71), .B(n_70), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_572), .Y(n_614) );
BUFx5_ASAP7_75t_L g615 ( .A(n_557), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_575), .B(n_559), .Y(n_616) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_568), .A2(n_73), .B(n_72), .Y(n_617) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_571), .A2(n_77), .B(n_75), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_572), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_556), .A2(n_361), .B(n_356), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_578), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_540), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_540), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_579), .B(n_19), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_553), .Y(n_628) );
NOR2x1_ASAP7_75t_SL g629 ( .A(n_575), .B(n_79), .Y(n_629) );
BUFx10_ASAP7_75t_L g630 ( .A(n_551), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_535), .B(n_405), .C(n_368), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_553), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_603), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_598), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_628), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_601), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_598), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_594), .B(n_19), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_628), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_632), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_632), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_590), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_589), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_593), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_585), .B(n_20), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_589), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_583), .Y(n_648) );
OAI21x1_ASAP7_75t_L g649 ( .A1(n_581), .A2(n_84), .B(n_82), .Y(n_649) );
BUFx12f_ASAP7_75t_L g650 ( .A(n_625), .Y(n_650) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_589), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_614), .Y(n_652) );
BUFx3_ASAP7_75t_L g653 ( .A(n_582), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_592), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_623), .A2(n_404), .B1(n_400), .B2(n_397), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_623), .A2(n_394), .B1(n_393), .B2(n_390), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_619), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_592), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_592), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_619), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_612), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_623), .A2(n_386), .B1(n_385), .B2(n_384), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_622), .Y(n_663) );
CKINVDCx11_ASAP7_75t_R g664 ( .A(n_630), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_627), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_622), .Y(n_666) );
OAI21x1_ASAP7_75t_L g667 ( .A1(n_599), .A2(n_86), .B(n_85), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_620), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_596), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_597), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_586), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_626), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_604), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_605), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_591), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_616), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_607), .Y(n_678) );
BUFx3_ASAP7_75t_L g679 ( .A(n_616), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_629), .B(n_29), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_605), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_615), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_615), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_608), .B(n_30), .Y(n_684) );
AO21x2_ASAP7_75t_L g685 ( .A1(n_602), .A2(n_33), .B(n_34), .Y(n_685) );
OR2x6_ASAP7_75t_L g686 ( .A(n_617), .B(n_37), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_618), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_611), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_600), .Y(n_689) );
BUFx2_ASAP7_75t_R g690 ( .A(n_606), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_613), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_584), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_595), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_587), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_609), .A2(n_39), .B1(n_40), .B2(n_41), .C1(n_42), .C2(n_90), .Y(n_695) );
INVx3_ASAP7_75t_L g696 ( .A(n_621), .Y(n_696) );
NAND2x1_ASAP7_75t_L g697 ( .A(n_631), .B(n_93), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_610), .B(n_39), .Y(n_698) );
BUFx4f_ASAP7_75t_SL g699 ( .A(n_624), .Y(n_699) );
BUFx2_ASAP7_75t_SL g700 ( .A(n_637), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_634), .B(n_40), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_636), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g704 ( .A(n_645), .B(n_42), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_641), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_642), .B(n_96), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_661), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_657), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_657), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_646), .B(n_684), .Y(n_710) );
OR2x2_ASAP7_75t_SL g711 ( .A(n_668), .B(n_102), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_660), .Y(n_712) );
AO31x2_ASAP7_75t_L g713 ( .A1(n_654), .A2(n_658), .A3(n_659), .B(n_688), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_660), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_635), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_666), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_638), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_643), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_679), .B(n_116), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_665), .B(n_117), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_663), .B(n_122), .Y(n_721) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_685), .B(n_123), .Y(n_722) );
CKINVDCx9p33_ASAP7_75t_R g723 ( .A(n_699), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_696), .B(n_126), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_677), .B(n_127), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_695), .B(n_128), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_652), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_633), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_648), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_669), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_675), .B(n_134), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_666), .B(n_254), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_673), .B(n_135), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_670), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_683), .B(n_136), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_670), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_639), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_698), .B(n_138), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_676), .A2(n_141), .B(n_144), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_685), .Y(n_740) );
INVxp33_ASAP7_75t_L g741 ( .A(n_664), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_693), .A2(n_146), .B1(n_147), .B2(n_149), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g743 ( .A1(n_680), .A2(n_150), .B(n_151), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_653), .B(n_154), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_653), .B(n_157), .Y(n_745) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_644), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_675), .B(n_158), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_681), .Y(n_748) );
BUFx4f_ASAP7_75t_SL g749 ( .A(n_650), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_647), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_655), .B(n_253), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_647), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_682), .B(n_162), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_644), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_689), .B(n_165), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_689), .B(n_671), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_692), .A2(n_170), .B1(n_171), .B2(n_173), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_655), .B(n_175), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_656), .B(n_187), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_644), .B(n_252), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_672), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_651), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_686), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_694), .B(n_651), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_651), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_656), .B(n_188), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_662), .B(n_190), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_686), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_667), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_687), .B(n_191), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_649), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_707), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_702), .B(n_691), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_703), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_705), .Y(n_775) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_700), .B(n_697), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_712), .B(n_674), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_710), .B(n_678), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_729), .B(n_690), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_727), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_730), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_714), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_728), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_763), .B(n_768), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_726), .A2(n_662), .B1(n_192), .B2(n_196), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_718), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_734), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_708), .B(n_197), .Y(n_788) );
INVx1_ASAP7_75t_SL g789 ( .A(n_750), .Y(n_789) );
NOR2xp67_ASAP7_75t_L g790 ( .A(n_739), .B(n_198), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_709), .Y(n_791) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_715), .Y(n_792) );
BUFx2_ASAP7_75t_L g793 ( .A(n_723), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_717), .B(n_200), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_716), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_752), .B(n_202), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_736), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_761), .Y(n_798) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_756), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_701), .B(n_211), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_748), .B(n_212), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_738), .B(n_214), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_737), .B(n_220), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_762), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_765), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_733), .B(n_228), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_764), .B(n_746), .Y(n_807) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_764), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_706), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_758), .A2(n_230), .B1(n_231), .B2(n_232), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_711), .B(n_234), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_740), .B(n_235), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_749), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_706), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_770), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_735), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_741), .B(n_236), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_731), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_754), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_731), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_747), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_747), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_755), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_755), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_704), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_773), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_781), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_772), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_778), .B(n_713), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_780), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_808), .B(n_713), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_782), .B(n_724), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_784), .B(n_722), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_784), .B(n_722), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_799), .B(n_769), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_799), .B(n_754), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_807), .B(n_787), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_789), .B(n_745), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_774), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_783), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_792), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_797), .B(n_719), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_795), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_775), .B(n_720), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_786), .B(n_725), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_798), .B(n_732), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_818), .B(n_771), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_791), .B(n_744), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_804), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_805), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_777), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_820), .B(n_771), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_821), .B(n_753), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_809), .B(n_753), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_822), .B(n_743), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_823), .B(n_760), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_824), .B(n_721), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_814), .B(n_767), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_827), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_828), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_841), .B(n_815), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_839), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_849), .B(n_779), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_829), .B(n_816), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_826), .B(n_819), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_843), .B(n_793), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_837), .B(n_825), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_851), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_830), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_850), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_831), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_836), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_840), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_840), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_861), .Y(n_875) );
NAND4xp75_ASAP7_75t_SL g876 ( .A(n_866), .B(n_790), .C(n_817), .D(n_855), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_859), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_860), .Y(n_878) );
INVxp67_ASAP7_75t_L g879 ( .A(n_870), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_867), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_871), .B(n_835), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_862), .Y(n_882) );
OAI21xp33_ASAP7_75t_L g883 ( .A1(n_863), .A2(n_855), .B(n_845), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_872), .A2(n_811), .B1(n_848), .B2(n_838), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_864), .B(n_831), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_877), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_878), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_884), .A2(n_857), .B1(n_858), .B2(n_844), .Y(n_888) );
AO22x1_ASAP7_75t_L g889 ( .A1(n_879), .A2(n_842), .B1(n_833), .B2(n_834), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_880), .A2(n_865), .B1(n_842), .B2(n_868), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_875), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_883), .A2(n_833), .B1(n_834), .B2(n_847), .Y(n_892) );
OAI32xp33_ASAP7_75t_L g893 ( .A1(n_881), .A2(n_813), .A3(n_806), .B1(n_846), .B2(n_854), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_891), .B(n_882), .Y(n_894) );
OAI211xp5_ASAP7_75t_L g895 ( .A1(n_893), .A2(n_785), .B(n_776), .C(n_885), .Y(n_895) );
AO22x1_ASAP7_75t_L g896 ( .A1(n_890), .A2(n_887), .B1(n_886), .B2(n_889), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_888), .A2(n_853), .B1(n_852), .B2(n_856), .Y(n_897) );
NAND3xp33_ASAP7_75t_SL g898 ( .A(n_895), .B(n_892), .C(n_810), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_894), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_897), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_896), .A2(n_803), .B(n_832), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_899), .Y(n_902) );
NOR2x1_ASAP7_75t_L g903 ( .A(n_898), .B(n_876), .Y(n_903) );
NOR3xp33_ASAP7_75t_L g904 ( .A(n_903), .B(n_900), .C(n_901), .Y(n_904) );
XNOR2x1_ASAP7_75t_L g905 ( .A(n_902), .B(n_802), .Y(n_905) );
NOR2x1p5_ASAP7_75t_L g906 ( .A(n_905), .B(n_800), .Y(n_906) );
NAND4xp75_ASAP7_75t_L g907 ( .A(n_904), .B(n_759), .C(n_766), .D(n_751), .Y(n_907) );
NOR2xp33_ASAP7_75t_R g908 ( .A(n_907), .B(n_237), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_908), .B(n_906), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_909), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_910), .B(n_874), .Y(n_911) );
OA22x2_ASAP7_75t_L g912 ( .A1(n_911), .A2(n_796), .B1(n_801), .B2(n_788), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_912), .A2(n_742), .B(n_757), .Y(n_913) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_913), .A2(n_812), .B(n_794), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_914), .A2(n_873), .B(n_869), .Y(n_915) );
AOI21xp33_ASAP7_75t_SL g916 ( .A1(n_915), .A2(n_242), .B(n_243), .Y(n_916) );
endmodule