module fake_netlist_1_12533_n_759 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_759);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_759;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_22), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_75), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_57), .B(n_85), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_94), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_102), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_60), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_88), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_35), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_64), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_83), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_15), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_10), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_25), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_27), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_11), .Y(n_131) );
INVxp33_ASAP7_75t_SL g132 ( .A(n_87), .Y(n_132) );
INVx4_ASAP7_75t_R g133 ( .A(n_24), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_30), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_22), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_21), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_38), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_19), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_66), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_40), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_73), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_58), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_47), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_10), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_37), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_15), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_29), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_147), .B(n_0), .Y(n_150) );
CKINVDCx11_ASAP7_75t_R g151 ( .A(n_129), .Y(n_151) );
INVx1_ASAP7_75t_SL g152 ( .A(n_148), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_107), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_116), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_136), .B(n_1), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
NOR2x1_ASAP7_75t_L g160 ( .A(n_136), .B(n_26), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_112), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_112), .Y(n_162) );
OR2x6_ASAP7_75t_L g163 ( .A(n_110), .B(n_2), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
CKINVDCx11_ASAP7_75t_R g166 ( .A(n_129), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_118), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_110), .B(n_3), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_155), .Y(n_170) );
BUFx10_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_158), .A2(n_107), .B1(n_108), .B2(n_146), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_158), .A2(n_131), .B1(n_111), .B2(n_146), .Y(n_173) );
BUFx8_ASAP7_75t_SL g174 ( .A(n_163), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_159), .B(n_130), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_169), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g181 ( .A(n_153), .B(n_131), .C(n_111), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_159), .B(n_147), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_161), .B(n_115), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_161), .B(n_117), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_162), .B(n_167), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
AND3x2_ASAP7_75t_L g196 ( .A(n_151), .B(n_114), .C(n_134), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_162), .B(n_144), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_167), .B(n_119), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_184), .B(n_152), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_184), .B(n_168), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_186), .B(n_168), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_174), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_184), .B(n_150), .Y(n_205) );
BUFx6f_ASAP7_75t_SL g206 ( .A(n_186), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_188), .B(n_163), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_188), .B(n_163), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_188), .B(n_125), .Y(n_210) );
INVx5_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_170), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_175), .B(n_137), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_186), .B(n_108), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_186), .B(n_127), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_175), .B(n_141), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_127), .B1(n_135), .B2(n_128), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_190), .A2(n_166), .B1(n_132), .B2(n_128), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_193), .B(n_145), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_190), .A2(n_135), .B1(n_139), .B2(n_160), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_193), .B(n_165), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_174), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_190), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_198), .B(n_165), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_176), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_190), .B(n_176), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_179), .B(n_143), .Y(n_229) );
AND2x6_ASAP7_75t_SL g230 ( .A(n_196), .B(n_139), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
OR2x4_ASAP7_75t_L g233 ( .A(n_196), .B(n_119), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_190), .B(n_164), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_198), .B(n_164), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_198), .B(n_120), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_176), .A2(n_138), .B1(n_149), .B2(n_123), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_179), .B(n_182), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_198), .B(n_120), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_225), .B(n_179), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_201), .A2(n_181), .B(n_178), .C(n_185), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_211), .B(n_176), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_203), .A2(n_180), .B(n_176), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_208), .B(n_198), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_214), .A2(n_180), .B1(n_178), .B2(n_185), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_204), .B(n_199), .C(n_183), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_211), .B(n_180), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
AO32x2_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_180), .A3(n_155), .B1(n_189), .B2(n_198), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_200), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_236), .A2(n_149), .B(n_122), .C(n_123), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_181), .B(n_189), .C(n_183), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_203), .A2(n_180), .B(n_189), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_217), .B(n_172), .C(n_173), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_223), .Y(n_259) );
INVx5_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_211), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_208), .B(n_189), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_189), .B(n_177), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_223), .B(n_172), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_240), .A2(n_173), .B(n_195), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_205), .B(n_171), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_222), .A2(n_170), .B(n_191), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_210), .B(n_171), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_215), .A2(n_197), .B1(n_195), .B2(n_192), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_239), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_235), .Y(n_273) );
CKINVDCx6p67_ASAP7_75t_R g274 ( .A(n_206), .Y(n_274) );
NOR2xp33_ASAP7_75t_R g275 ( .A(n_206), .B(n_194), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AO31x2_ASAP7_75t_L g277 ( .A1(n_249), .A2(n_232), .A3(n_170), .B(n_191), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_271), .A2(n_228), .B1(n_237), .B2(n_206), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_270), .A2(n_219), .B(n_229), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_220), .B(n_187), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_SL g282 ( .A1(n_245), .A2(n_221), .B(n_197), .C(n_192), .Y(n_282) );
AOI221xp5_ASAP7_75t_SL g283 ( .A1(n_242), .A2(n_234), .B1(n_194), .B2(n_216), .C(n_213), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_256), .A2(n_234), .B(n_228), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_228), .B(n_212), .Y(n_285) );
O2A1O1Ixp5_ASAP7_75t_L g286 ( .A1(n_245), .A2(n_224), .B(n_170), .C(n_177), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_269), .A2(n_212), .B(n_177), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_265), .A2(n_227), .B1(n_231), .B2(n_202), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_254), .B(n_218), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
INVx3_ASAP7_75t_SL g292 ( .A(n_274), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_272), .Y(n_293) );
O2A1O1Ixp5_ASAP7_75t_SL g294 ( .A1(n_251), .A2(n_124), .B(n_126), .C(n_138), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_259), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_255), .A2(n_194), .B(n_227), .C(n_202), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_270), .A2(n_202), .B(n_231), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_268), .A2(n_231), .B(n_194), .C(n_211), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_248), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_300), .B(n_250), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_299), .B(n_260), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_300), .B(n_243), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_299), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_299), .B(n_263), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_279), .A2(n_268), .B(n_246), .C(n_257), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_299), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_292), .A2(n_233), .B1(n_247), .B2(n_252), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_292), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_264), .B(n_187), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_289), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_277), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_277), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_287), .A2(n_285), .B(n_294), .Y(n_318) );
INVx4_ASAP7_75t_SL g319 ( .A(n_292), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_266), .B(n_251), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_290), .B(n_273), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_288), .B(n_241), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_305), .B(n_283), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_310), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_322), .A2(n_262), .B1(n_284), .B2(n_278), .C(n_296), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_318), .A2(n_284), .B(n_287), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_310), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_307), .B(n_253), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_319), .B(n_275), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_303), .B(n_281), .Y(n_334) );
OAI211xp5_ASAP7_75t_L g335 ( .A1(n_301), .A2(n_275), .B(n_113), .C(n_244), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_306), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_309), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_309), .B(n_289), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_316), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_318), .A2(n_286), .B(n_276), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_322), .A2(n_233), .B1(n_295), .B2(n_260), .Y(n_348) );
AOI21xp5_ASAP7_75t_SL g349 ( .A1(n_317), .A2(n_289), .B(n_291), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_307), .B(n_253), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_346), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_325), .B(n_321), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_336), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_325), .B(n_321), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_326), .B(n_320), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_336), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_346), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_329), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_338), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_338), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_341), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_333), .B(n_320), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_320), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_333), .B(n_320), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_340), .B(n_314), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_341), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_340), .B(n_314), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
OR2x2_ASAP7_75t_SL g384 ( .A(n_334), .B(n_319), .Y(n_384) );
NOR2x1_ASAP7_75t_SL g385 ( .A(n_339), .B(n_309), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_352), .B(n_314), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_314), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_307), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_328), .B(n_253), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_324), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_328), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_324), .B(n_323), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_328), .B(n_253), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_331), .B(n_307), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_350), .B(n_281), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_328), .B(n_122), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_350), .B(n_327), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_337), .B(n_230), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_385), .A2(n_349), .B(n_332), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_355), .B(n_344), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_382), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_355), .B(n_344), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_399), .B(n_344), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_355), .B(n_345), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_399), .B(n_345), .Y(n_412) );
AND2x4_ASAP7_75t_SL g413 ( .A(n_382), .B(n_337), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_357), .B(n_345), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_382), .B(n_337), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_354), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_363), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_371), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_357), .B(n_351), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_357), .B(n_327), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_384), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_356), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_366), .B(n_319), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_356), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_348), .B1(n_311), .B2(n_335), .C(n_142), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_371), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_401), .B(n_351), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_389), .B(n_351), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_359), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_359), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_359), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_369), .B(n_319), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_360), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_389), .B(n_342), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
INVx5_ASAP7_75t_L g442 ( .A(n_382), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_389), .B(n_342), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_401), .B(n_319), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_384), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_374), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_396), .B(n_342), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_402), .B(n_335), .Y(n_448) );
NAND5xp2_ASAP7_75t_SL g449 ( .A(n_385), .B(n_312), .C(n_308), .D(n_5), .E(n_6), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_381), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_402), .B(n_124), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_396), .B(n_342), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_366), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_381), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_376), .B(n_349), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_365), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_369), .B(n_144), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_396), .B(n_126), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_358), .B(n_140), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_364), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_365), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_383), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_358), .B(n_140), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_366), .Y(n_464) );
INVx6_ASAP7_75t_L g465 ( .A(n_366), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_364), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_358), .B(n_142), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_383), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_375), .B(n_281), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_376), .B(n_302), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_379), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_390), .B(n_302), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_388), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_375), .B(n_3), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_365), .Y(n_475) );
NAND2x1_ASAP7_75t_L g476 ( .A(n_369), .B(n_289), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_390), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_417), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_413), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_460), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_406), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_473), .B(n_398), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_440), .B(n_375), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_440), .B(n_378), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_413), .Y(n_485) );
AND3x2_ASAP7_75t_L g486 ( .A(n_438), .B(n_373), .C(n_403), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_448), .B(n_388), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_443), .B(n_378), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_406), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_416), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_470), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_458), .B(n_393), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_458), .B(n_393), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_444), .A2(n_373), .B1(n_398), .B2(n_369), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_416), .Y(n_497) );
OR2x6_ASAP7_75t_L g498 ( .A(n_405), .B(n_366), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_470), .B(n_379), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_459), .B(n_400), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_459), .B(n_463), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_433), .B(n_367), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_404), .B(n_367), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_426), .B(n_367), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_451), .B(n_366), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_466), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_418), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_429), .B(n_366), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_418), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_420), .B(n_368), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_463), .B(n_400), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_407), .B(n_391), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_407), .B(n_391), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_467), .B(n_378), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_421), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_420), .B(n_368), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_421), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_471), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_467), .B(n_380), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_409), .B(n_394), .Y(n_520) );
NOR2xp33_ASAP7_75t_SL g521 ( .A(n_427), .B(n_302), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_439), .B(n_368), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_428), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_409), .B(n_394), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_474), .B(n_380), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_411), .B(n_380), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_430), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_425), .B(n_377), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_445), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_474), .B(n_386), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_419), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_442), .B(n_370), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_410), .B(n_370), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_430), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_422), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_443), .B(n_386), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_447), .B(n_386), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_447), .B(n_387), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_452), .B(n_387), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_410), .B(n_370), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_452), .B(n_387), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_422), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_434), .B(n_392), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_442), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_434), .B(n_392), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_411), .B(n_397), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_477), .B(n_377), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_412), .B(n_372), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_412), .B(n_372), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_415), .B(n_397), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_477), .B(n_372), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_423), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_415), .B(n_392), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_419), .A2(n_395), .B1(n_276), .B2(n_293), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_423), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_442), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_432), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_395), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_414), .B(n_395), .Y(n_559) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_438), .B(n_395), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_432), .Y(n_561) );
INVxp33_ASAP7_75t_L g562 ( .A(n_419), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_431), .B(n_294), .C(n_5), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_435), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_441), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_441), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_480), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_483), .B(n_462), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_528), .B(n_462), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g570 ( .A1(n_505), .A2(n_457), .B(n_468), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_480), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_529), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_544), .B(n_442), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_484), .B(n_424), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_484), .B(n_468), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_455), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_528), .B(n_457), .C(n_455), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_505), .A2(n_457), .B(n_472), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_487), .B(n_408), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_487), .B(n_446), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_488), .B(n_446), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_536), .B(n_450), .Y(n_585) );
INVx6_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_536), .B(n_424), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_481), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_499), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_537), .B(n_450), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_537), .B(n_424), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_538), .B(n_454), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_560), .B(n_442), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_538), .B(n_454), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_493), .B(n_472), .C(n_408), .D(n_438), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_539), .B(n_408), .Y(n_598) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_562), .A2(n_476), .B(n_449), .C(n_453), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_489), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_539), .B(n_469), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_541), .B(n_453), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_479), .B(n_465), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_544), .B(n_465), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_485), .B(n_464), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_541), .B(n_435), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_546), .B(n_436), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_510), .Y(n_609) );
NAND2xp33_ASAP7_75t_L g610 ( .A(n_562), .B(n_449), .Y(n_610) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_498), .A2(n_464), .B(n_476), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_496), .A2(n_465), .B1(n_475), .B2(n_461), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g613 ( .A(n_556), .B(n_436), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_497), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_501), .B(n_465), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_482), .B(n_437), .Y(n_616) );
NOR2x1p5_ASAP7_75t_L g617 ( .A(n_525), .B(n_437), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_516), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_507), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_556), .B(n_456), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_503), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_491), .B(n_456), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_495), .A2(n_461), .B1(n_475), .B2(n_395), .C1(n_194), .C2(n_9), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_550), .B(n_395), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_498), .A2(n_395), .B1(n_177), .B2(n_187), .C(n_191), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_526), .B(n_4), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_509), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_515), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_517), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_535), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_530), .B(n_4), .Y(n_631) );
AOI31xp33_ASAP7_75t_L g632 ( .A1(n_508), .A2(n_282), .A3(n_244), .B(n_280), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_542), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_552), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_555), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_504), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_512), .B(n_6), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_532), .A2(n_293), .B(n_280), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_557), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_502), .B(n_7), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_561), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_565), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_SL g643 ( .A1(n_496), .A2(n_7), .B(n_8), .C(n_11), .Y(n_643) );
NOR4xp25_ASAP7_75t_L g644 ( .A(n_532), .B(n_8), .C(n_12), .D(n_13), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_601), .B(n_543), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_569), .B(n_486), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_596), .A2(n_498), .B(n_524), .Y(n_647) );
XNOR2x1_ASAP7_75t_L g648 ( .A(n_626), .B(n_486), .Y(n_648) );
OAI321xp33_ASAP7_75t_L g649 ( .A1(n_596), .A2(n_547), .A3(n_519), .B1(n_514), .B2(n_500), .C(n_511), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_567), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_571), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_576), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_610), .A2(n_521), .B(n_554), .C(n_563), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_573), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_644), .A2(n_558), .B1(n_566), .B2(n_545), .C(n_543), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_568), .Y(n_657) );
OAI311xp33_ASAP7_75t_L g658 ( .A1(n_623), .A2(n_522), .A3(n_559), .B1(n_551), .C1(n_533), .Y(n_658) );
OAI322xp33_ASAP7_75t_L g659 ( .A1(n_640), .A2(n_549), .A3(n_548), .B1(n_540), .B2(n_558), .C1(n_513), .C2(n_520), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_584), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_620), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_620), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_572), .B(n_545), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_578), .A2(n_574), .B1(n_586), .B2(n_617), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_594), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_623), .B(n_494), .C(n_478), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_612), .B(n_553), .C(n_564), .D(n_534), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_644), .A2(n_564), .B(n_534), .C(n_527), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_582), .B(n_478), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_613), .A2(n_527), .B(n_523), .C(n_494), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_588), .Y(n_671) );
OAI21xp33_ASAP7_75t_SL g672 ( .A1(n_593), .A2(n_523), .B(n_492), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_600), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_631), .A2(n_492), .B1(n_191), .B2(n_187), .C1(n_133), .C2(n_18), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_608), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_643), .A2(n_298), .B(n_133), .C(n_16), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_575), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_602), .B(n_12), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_580), .B(n_289), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_637), .Y(n_680) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_632), .A2(n_261), .B(n_241), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_583), .B(n_14), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_587), .B(n_14), .Y(n_683) );
NOR3xp33_ASAP7_75t_SL g684 ( .A(n_599), .B(n_16), .C(n_17), .Y(n_684) );
AOI33xp33_ASAP7_75t_L g685 ( .A1(n_609), .A2(n_17), .A3(n_19), .B1(n_20), .B2(n_21), .B3(n_23), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_581), .A2(n_276), .B1(n_293), .B2(n_280), .Y(n_686) );
AOI21xp33_ASAP7_75t_SL g687 ( .A1(n_597), .A2(n_20), .B(n_23), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_591), .B(n_24), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_586), .A2(n_291), .B1(n_261), .B2(n_260), .Y(n_689) );
OAI33xp33_ASAP7_75t_L g690 ( .A1(n_585), .A2(n_592), .A3(n_590), .B1(n_639), .B2(n_641), .B3(n_614), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_609), .B(n_28), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g693 ( .A1(n_618), .A2(n_291), .B1(n_224), .B2(n_272), .C1(n_42), .C2(n_43), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_619), .Y(n_694) );
NOR4xp25_ASAP7_75t_L g695 ( .A(n_658), .B(n_625), .C(n_570), .D(n_605), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_692), .B(n_598), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_687), .A2(n_632), .B(n_570), .C(n_579), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_649), .A2(n_604), .B1(n_577), .B2(n_579), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_690), .A2(n_615), .B1(n_627), .B2(n_629), .C(n_635), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_646), .A2(n_656), .B1(n_667), .B2(n_690), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_647), .A2(n_603), .B(n_611), .C(n_642), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_659), .A2(n_634), .B1(n_633), .B2(n_630), .C(n_628), .Y(n_702) );
OAI31xp33_ASAP7_75t_SL g703 ( .A1(n_664), .A2(n_611), .A3(n_616), .B(n_589), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_656), .A2(n_622), .B(n_606), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_672), .A2(n_636), .B(n_621), .C(n_607), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_684), .A2(n_624), .B(n_638), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_648), .A2(n_291), .B1(n_297), .B2(n_272), .Y(n_707) );
AOI32xp33_ASAP7_75t_L g708 ( .A1(n_654), .A2(n_291), .A3(n_36), .B1(n_41), .B2(n_44), .Y(n_708) );
O2A1O1Ixp5_ASAP7_75t_L g709 ( .A1(n_668), .A2(n_32), .B(n_45), .C(n_46), .Y(n_709) );
NOR2x1_ASAP7_75t_SL g710 ( .A(n_668), .B(n_291), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_684), .A2(n_48), .B(n_49), .C(n_50), .Y(n_711) );
OAI211xp5_ASAP7_75t_SL g712 ( .A1(n_685), .A2(n_53), .B(n_54), .C(n_55), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_655), .A2(n_56), .B(n_59), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_645), .B(n_61), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_669), .B(n_62), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_680), .A2(n_272), .B1(n_65), .B2(n_67), .C(n_68), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_660), .Y(n_717) );
OAI31xp33_ASAP7_75t_L g718 ( .A1(n_670), .A2(n_63), .A3(n_69), .B(n_70), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_674), .A2(n_71), .B(n_72), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_676), .A2(n_74), .B(n_76), .C(n_77), .Y(n_720) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_681), .A2(n_239), .B(n_209), .C(n_81), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_695), .A2(n_680), .B1(n_655), .B2(n_666), .C(n_682), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g723 ( .A1(n_703), .A2(n_693), .B(n_676), .C(n_650), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_704), .B(n_677), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_717), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_705), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_700), .B(n_691), .C(n_678), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_698), .A2(n_651), .B1(n_694), .B2(n_671), .C(n_673), .Y(n_728) );
NOR2xp33_ASAP7_75t_R g729 ( .A(n_714), .B(n_688), .Y(n_729) );
AOI321xp33_ASAP7_75t_L g730 ( .A1(n_701), .A2(n_683), .A3(n_665), .B1(n_689), .B2(n_657), .C(n_653), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_696), .B(n_662), .Y(n_731) );
AOI211x1_ASAP7_75t_SL g732 ( .A1(n_712), .A2(n_661), .B(n_679), .C(n_675), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g733 ( .A1(n_702), .A2(n_652), .B1(n_663), .B2(n_686), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g734 ( .A1(n_697), .A2(n_78), .B(n_80), .Y(n_734) );
NAND5xp2_ASAP7_75t_L g735 ( .A(n_708), .B(n_82), .C(n_84), .D(n_86), .E(n_90), .Y(n_735) );
NOR2x1p5_ASAP7_75t_L g736 ( .A(n_727), .B(n_715), .Y(n_736) );
NAND3xp33_ASAP7_75t_SL g737 ( .A(n_732), .B(n_711), .C(n_721), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_730), .A2(n_707), .B1(n_706), .B2(n_699), .C(n_719), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_734), .B(n_712), .C(n_709), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_723), .B(n_709), .C(n_720), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_722), .A2(n_718), .B1(n_716), .B2(n_713), .C(n_710), .Y(n_741) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_726), .B(n_91), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_742), .B(n_731), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_740), .B(n_728), .Y(n_744) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_737), .B(n_735), .C(n_724), .D(n_725), .Y(n_745) );
OAI211xp5_ASAP7_75t_SL g746 ( .A1(n_738), .A2(n_733), .B(n_729), .C(n_731), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_744), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_746), .Y(n_748) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_745), .B(n_736), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_747), .Y(n_750) );
XNOR2xp5_ASAP7_75t_L g751 ( .A(n_749), .B(n_743), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_750), .Y(n_752) );
AOI22xp5_ASAP7_75t_SL g753 ( .A1(n_751), .A2(n_749), .B1(n_748), .B2(n_739), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_752), .A2(n_741), .B1(n_239), .B2(n_209), .Y(n_754) );
OAI222xp33_ASAP7_75t_L g755 ( .A1(n_753), .A2(n_93), .B1(n_95), .B2(n_96), .C1(n_97), .C2(n_98), .Y(n_755) );
OAI21x1_ASAP7_75t_SL g756 ( .A1(n_754), .A2(n_99), .B(n_100), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_755), .B(n_209), .C(n_239), .Y(n_757) );
AO221x2_ASAP7_75t_SL g758 ( .A1(n_756), .A2(n_101), .B1(n_103), .B2(n_104), .C(n_105), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_758), .A2(n_757), .B1(n_209), .B2(n_106), .Y(n_759) );
endmodule