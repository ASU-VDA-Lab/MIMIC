module real_jpeg_16112_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_19),
.Y(n_18)
);

AND2x4_ASAP7_75t_SL g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_0),
.B(n_48),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_0),
.B(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_62),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_6),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_6),
.B(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_102),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_100),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_64),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_64),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_35),
.C(n_49),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_14),
.B(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_26),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_16),
.A2(n_27),
.B(n_34),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_16),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

NOR2x1_ASAP7_75t_R g16 ( 
.A(n_17),
.B(n_22),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_17),
.A2(n_18),
.B1(n_96),
.B2(n_99),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_30),
.B(n_32),
.Y(n_29)
);

NAND2x1p5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_30),
.Y(n_32)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_21),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_22),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_22),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_27),
.A2(n_124),
.B(n_127),
.C(n_133),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_27),
.B(n_124),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_27),
.A2(n_33),
.B1(n_124),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_30),
.A2(n_113),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_30),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_35),
.A2(n_49),
.B1(n_50),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.C(n_45),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_36),
.A2(n_37),
.B1(n_45),
.B2(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_40),
.A2(n_41),
.B1(n_84),
.B2(n_89),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_40),
.A2(n_41),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_45),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_57),
.C(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_82),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_81),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_74),
.B1(n_75),
.B2(n_80),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_85),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_140),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_96),
.Y(n_99)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_112),
.B(n_113),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_121),
.B(n_148),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_107),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_117),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_117),
.B1(n_118),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_137),
.B(n_147),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_134),
.Y(n_147)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_128),
.Y(n_131)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_143),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B(n_146),
.Y(n_137)
);


endmodule