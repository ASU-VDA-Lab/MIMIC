module fake_jpeg_22236_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_39),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_53),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_19),
.B1(n_20),
.B2(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_28),
.B1(n_27),
.B2(n_17),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_68),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_56),
.B1(n_52),
.B2(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_89),
.Y(n_93)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_75),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_15),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_33),
.B1(n_18),
.B2(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_74),
.B1(n_88),
.B2(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_24),
.B1(n_26),
.B2(n_56),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_52),
.B1(n_56),
.B2(n_21),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_76),
.B1(n_83),
.B2(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_60),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_53),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_22),
.B1(n_35),
.B2(n_15),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_11),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_68),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_123),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

OAI211xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_74),
.B(n_59),
.C(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_127),
.B1(n_65),
.B2(n_112),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_72),
.C(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_130),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_64),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_97),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_62),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_61),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_61),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_116),
.C(n_93),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_116),
.C(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_67),
.B(n_80),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_111),
.B(n_115),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_99),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_151),
.Y(n_168)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_136),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_159),
.B1(n_164),
.B2(n_126),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_114),
.C(n_108),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_114),
.C(n_115),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_98),
.B(n_3),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_104),
.B(n_3),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_2),
.B(n_4),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_2),
.B(n_4),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_174),
.C(n_146),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_134),
.A3(n_118),
.B1(n_126),
.B2(n_127),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_118),
.B1(n_123),
.B2(n_137),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_131),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_179),
.A2(n_120),
.B(n_164),
.C(n_8),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_129),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_174),
.C(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_138),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_145),
.A3(n_157),
.B1(n_156),
.B2(n_158),
.C1(n_129),
.C2(n_154),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_168),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_149),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_172),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_178),
.B(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_192),
.C(n_194),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_173),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_151),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_5),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_156),
.C(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_202),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_10),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_200),
.B(n_201),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_183),
.B(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_184),
.C(n_186),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.B(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_204),
.B1(n_187),
.B2(n_8),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_147),
.B1(n_14),
.B2(n_13),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_189),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_212),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_187),
.C(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_9),
.B1(n_10),
.B2(n_208),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_201),
.B(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_6),
.C(n_9),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_223),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_225),
.C(n_217),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_229),
.CI(n_223),
.CON(n_230),
.SN(n_230)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_215),
.C(n_225),
.Y(n_229)
);


endmodule