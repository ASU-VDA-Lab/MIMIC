module fake_jpeg_16541_n_386 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_47),
.Y(n_88)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_14),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_67),
.B(n_79),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_25),
.B(n_31),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_81),
.B(n_35),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_90),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_34),
.B1(n_26),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_76),
.A2(n_103),
.B1(n_105),
.B2(n_1),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_26),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_84),
.A2(n_85),
.B1(n_9),
.B2(n_10),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_18),
.B1(n_30),
.B2(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_102),
.Y(n_130)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_45),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_51),
.A2(n_20),
.B1(n_19),
.B2(n_24),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_20),
.B1(n_24),
.B2(n_31),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_30),
.Y(n_108)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_39),
.B(n_30),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_111),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_18),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_123),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_62),
.B1(n_13),
.B2(n_22),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_118),
.A2(n_126),
.B(n_127),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_119),
.B(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_32),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_124),
.B(n_131),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_32),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_129),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_68),
.A2(n_35),
.B1(n_22),
.B2(n_4),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_68),
.A2(n_35),
.B1(n_22),
.B2(n_5),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_96),
.B1(n_98),
.B2(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_133),
.B1(n_136),
.B2(n_149),
.Y(n_175)
);

NAND2x1_ASAP7_75t_SL g131 ( 
.A(n_86),
.B(n_32),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_21),
.C(n_58),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_140),
.C(n_144),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_58),
.B1(n_54),
.B2(n_21),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_21),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_167),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_76),
.B1(n_70),
.B2(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_142),
.B1(n_107),
.B2(n_66),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_21),
.C(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_113),
.B1(n_101),
.B2(n_72),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_2),
.C(n_8),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_92),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_84),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_77),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_12),
.B1(n_71),
.B2(n_136),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_106),
.B(n_11),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_168),
.C(n_71),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_114),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_115),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_77),
.A2(n_11),
.B1(n_12),
.B2(n_107),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_11),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_66),
.B(n_115),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_171),
.B(n_179),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_185),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_173),
.A2(n_176),
.B1(n_188),
.B2(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_180),
.B(n_190),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_124),
.A2(n_106),
.B(n_85),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_158),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_133),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_125),
.A2(n_159),
.B1(n_123),
.B2(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_78),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_198),
.Y(n_237)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_12),
.C(n_134),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_215),
.C(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_200),
.Y(n_249)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_201),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_148),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_202),
.B(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_121),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_214),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_12),
.B1(n_140),
.B2(n_147),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_211),
.A2(n_181),
.B1(n_205),
.B2(n_197),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_137),
.B(n_159),
.C(n_162),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_162),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_SL g291 ( 
.A(n_217),
.B(n_243),
.C(n_232),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_218),
.A2(n_230),
.B(n_234),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_254),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_SL g223 ( 
.A(n_188),
.B(n_147),
.C(n_151),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_223),
.B(n_251),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_187),
.B(n_178),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_256),
.B(n_234),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_182),
.C(n_207),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_228),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_144),
.C(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_170),
.A2(n_146),
.B1(n_151),
.B2(n_161),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_257),
.B1(n_206),
.B2(n_213),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_243),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_170),
.A2(n_154),
.B(n_181),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_154),
.C(n_199),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_242),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_178),
.B(n_173),
.C(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_208),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_175),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_169),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_245),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_174),
.C(n_177),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_189),
.B(n_200),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_176),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_263),
.B1(n_288),
.B2(n_276),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_206),
.B1(n_213),
.B2(n_201),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_214),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_269),
.Y(n_293)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_184),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_225),
.C(n_228),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_184),
.C(n_236),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_256),
.C(n_246),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_247),
.B(n_267),
.Y(n_314)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_278),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_221),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_286),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_222),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_281),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_218),
.B(n_248),
.C(n_242),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_287),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_238),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_257),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_230),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_220),
.C(n_229),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_220),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_233),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_306),
.Y(n_320)
);

NAND4xp25_ASAP7_75t_SL g300 ( 
.A(n_265),
.B(n_252),
.C(n_249),
.D(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_292),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_314),
.B(n_285),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_237),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_311),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_238),
.C(n_250),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_290),
.A2(n_247),
.B1(n_250),
.B2(n_289),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_313),
.A2(n_316),
.B1(n_273),
.B2(n_266),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_309),
.B1(n_301),
.B2(n_318),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_282),
.B1(n_281),
.B2(n_262),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_278),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_321),
.B(n_322),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_297),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_270),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_323),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_263),
.B1(n_261),
.B2(n_285),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_325),
.A2(n_337),
.B1(n_303),
.B2(n_312),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_304),
.Y(n_326)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_305),
.B(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_269),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_329),
.A2(n_338),
.B1(n_293),
.B2(n_314),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_298),
.B(n_293),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_338),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_335),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_295),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_340),
.C(n_294),
.Y(n_341)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_316),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_334),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_344),
.A2(n_350),
.B1(n_351),
.B2(n_354),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_311),
.C(n_299),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_352),
.C(n_334),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_332),
.A2(n_298),
.B1(n_306),
.B2(n_313),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_301),
.C(n_312),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_348),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_333),
.B1(n_329),
.B2(n_337),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_326),
.B1(n_335),
.B2(n_340),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_358),
.A2(n_361),
.B1(n_368),
.B2(n_352),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_320),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_362),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_366),
.B(n_367),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_326),
.B1(n_336),
.B2(n_320),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_349),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_355),
.C(n_354),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_357),
.B1(n_342),
.B2(n_350),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_346),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_372),
.B(n_362),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_357),
.B1(n_342),
.B2(n_356),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_347),
.C(n_366),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_347),
.B(n_346),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_374),
.A2(n_358),
.B(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_375),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_377),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_380),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_381),
.A2(n_379),
.B(n_371),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_370),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_378),
.Y(n_384)
);

OAI211xp5_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_374),
.B(n_369),
.C(n_360),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_363),
.Y(n_386)
);


endmodule