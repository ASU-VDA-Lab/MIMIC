module fake_netlist_1_7027_n_697 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_27), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_19), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_39), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_29), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_75), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_9), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_34), .Y(n_84) );
NOR2xp67_ASAP7_75t_L g85 ( .A(n_54), .B(n_67), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_26), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_49), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_40), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_0), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_63), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_66), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_10), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_5), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_47), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_48), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_0), .B(n_36), .Y(n_100) );
INVx4_ASAP7_75t_R g101 ( .A(n_52), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_20), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_25), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_11), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_42), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_64), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_59), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_11), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_57), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_33), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_32), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_2), .Y(n_119) );
CKINVDCx14_ASAP7_75t_R g120 ( .A(n_3), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_7), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_38), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_16), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_116), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
NOR2x1_ASAP7_75t_L g128 ( .A(n_104), .B(n_1), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_106), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_104), .B(n_2), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_82), .B(n_3), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_118), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_120), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_86), .B(n_4), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_91), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_118), .B(n_8), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_90), .B(n_9), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_95), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_95), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_94), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_94), .B(n_12), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_77), .B(n_50), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_96), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_86), .B(n_13), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_78), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_79), .Y(n_159) );
NOR2x1_ASAP7_75t_L g160 ( .A(n_84), .B(n_107), .Y(n_160) );
NAND2xp33_ASAP7_75t_SL g161 ( .A(n_96), .B(n_14), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_97), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_102), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_114), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_114), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_137), .A2(n_121), .B1(n_124), .B2(n_108), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_146), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_153), .B(n_109), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_153), .B(n_121), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_165), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_139), .B(n_153), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_139), .B(n_79), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_125), .Y(n_181) );
NOR2x1p5_ASAP7_75t_L g182 ( .A(n_126), .B(n_111), .Y(n_182) );
NAND3xp33_ASAP7_75t_L g183 ( .A(n_132), .B(n_154), .C(n_156), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_134), .B(n_80), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_159), .B(n_80), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_125), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
NAND2xp33_ASAP7_75t_L g188 ( .A(n_155), .B(n_81), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_134), .B(n_81), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_145), .B(n_105), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_125), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_125), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_131), .A2(n_115), .B1(n_119), .B2(n_100), .Y(n_195) );
NAND3x1_ASAP7_75t_L g196 ( .A(n_137), .B(n_122), .C(n_103), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_134), .B(n_110), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_145), .B(n_88), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_129), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_163), .B(n_110), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_151), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_131), .B(n_92), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_129), .Y(n_209) );
INVxp33_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_127), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_129), .Y(n_213) );
INVxp33_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_128), .B(n_117), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_166), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_163), .B(n_92), .Y(n_219) );
AND2x6_ASAP7_75t_L g220 ( .A(n_128), .B(n_101), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_135), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_136), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_149), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_140), .B(n_88), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_141), .B(n_123), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_149), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_212), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_223), .B(n_141), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_177), .B(n_160), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_211), .B(n_136), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_172), .B(n_160), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_227), .B(n_147), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_172), .B(n_148), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_175), .B(n_172), .Y(n_238) );
AO21x1_ASAP7_75t_L g239 ( .A1(n_188), .A2(n_215), .B(n_211), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_204), .B(n_147), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_225), .A2(n_161), .B1(n_148), .B2(n_138), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_222), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_222), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_219), .B(n_127), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_170), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_188), .A2(n_127), .B(n_162), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_183), .B(n_164), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_200), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_180), .B(n_164), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_216), .A2(n_144), .B1(n_150), .B2(n_158), .Y(n_251) );
NOR2x1_ASAP7_75t_L g252 ( .A(n_182), .B(n_152), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_201), .Y(n_254) );
NOR2xp33_ASAP7_75t_R g255 ( .A(n_221), .B(n_155), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_199), .B(n_158), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_199), .B(n_208), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_211), .B(n_162), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_169), .A2(n_150), .B1(n_162), .B2(n_149), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_187), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_174), .A2(n_130), .B1(n_144), .B2(n_113), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_178), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_208), .B(n_144), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_210), .A2(n_130), .B1(n_144), .B2(n_85), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_192), .B(n_185), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_205), .A2(n_15), .B1(n_17), .B2(n_18), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_195), .B(n_15), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_184), .B(n_17), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_189), .B(n_22), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_23), .B1(n_28), .B2(n_30), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_193), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_198), .B(n_31), .Y(n_278) );
NOR2xp33_ASAP7_75t_SL g279 ( .A(n_215), .B(n_35), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_228), .B(n_41), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_215), .B(n_43), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_200), .B(n_44), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_197), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_206), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_220), .B(n_46), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_220), .B(n_53), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_207), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_209), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_220), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_202), .B(n_55), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_229), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_214), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_220), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_235), .B(n_220), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_246), .A2(n_190), .B(n_202), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_294), .Y(n_299) );
AO32x1_ASAP7_75t_L g300 ( .A1(n_265), .A2(n_194), .A3(n_173), .B1(n_181), .B2(n_186), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_271), .B(n_196), .Y(n_301) );
CKINVDCx8_ASAP7_75t_R g302 ( .A(n_271), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_241), .A2(n_214), .B1(n_176), .B2(n_168), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_248), .Y(n_305) );
AOI222xp33_ASAP7_75t_L g306 ( .A1(n_237), .A2(n_176), .B1(n_170), .B2(n_217), .C1(n_221), .C2(n_216), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_232), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_294), .Y(n_310) );
AOI21x1_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_190), .B(n_226), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_243), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_238), .A2(n_240), .B(n_236), .C(n_231), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_266), .B(n_220), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_238), .A2(n_229), .B(n_226), .C(n_213), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_233), .B(n_217), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_248), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_235), .B(n_216), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_253), .B(n_216), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_263), .A2(n_196), .B(n_173), .C(n_181), .Y(n_324) );
HAxp5_ASAP7_75t_L g325 ( .A(n_237), .B(n_216), .CON(n_325), .SN(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_254), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_255), .B(n_203), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_249), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_245), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_248), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_252), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_233), .A2(n_216), .B1(n_203), .B2(n_202), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_247), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_250), .B(n_203), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_264), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_244), .A2(n_203), .B(n_202), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_250), .A2(n_194), .B(n_186), .C(n_171), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_247), .B(n_171), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_255), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_257), .B(n_191), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_256), .A2(n_56), .B(n_58), .C(n_60), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_234), .A2(n_191), .B1(n_62), .B2(n_65), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_302), .B(n_286), .Y(n_348) );
CKINVDCx11_ASAP7_75t_R g349 ( .A(n_338), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_301), .A2(n_251), .B1(n_262), .B2(n_286), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_311), .A2(n_281), .B(n_291), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_337), .A2(n_291), .B(n_278), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_301), .A2(n_251), .B1(n_262), .B2(n_284), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_SL g355 ( .A1(n_339), .A2(n_282), .B(n_274), .C(n_272), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_304), .B(n_295), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_301), .A2(n_249), .B1(n_290), .B2(n_270), .Y(n_357) );
AO31x2_ASAP7_75t_L g358 ( .A1(n_343), .A2(n_239), .A3(n_274), .B(n_287), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_306), .A2(n_242), .B1(n_259), .B2(n_269), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_296), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_344), .A2(n_275), .B(n_280), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_259), .B(n_269), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_268), .B(n_230), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_332), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_296), .Y(n_370) );
OAI21x1_ASAP7_75t_SL g371 ( .A1(n_324), .A2(n_261), .B(n_293), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_298), .A2(n_258), .B(n_289), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_299), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_297), .B(n_292), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_298), .A2(n_288), .B(n_273), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_348), .A2(n_306), .B1(n_334), .B2(n_318), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
OR2x6_ASAP7_75t_L g380 ( .A(n_361), .B(n_322), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_317), .B1(n_315), .B2(n_303), .Y(n_381) );
AO221x2_ASAP7_75t_L g382 ( .A1(n_369), .A2(n_372), .B1(n_363), .B2(n_364), .C(n_359), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_369), .B(n_314), .Y(n_383) );
AOI21x1_ASAP7_75t_L g384 ( .A1(n_366), .A2(n_323), .B(n_300), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_308), .B1(n_310), .B2(n_335), .Y(n_385) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_366), .A2(n_323), .B(n_300), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_316), .B(n_345), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_351), .A2(n_310), .B1(n_329), .B2(n_341), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_359), .A2(n_331), .B1(n_297), .B2(n_322), .C(n_336), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_325), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_328), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
OR2x6_ASAP7_75t_L g394 ( .A(n_361), .B(n_307), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_300), .B(n_279), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_335), .B1(n_333), .B2(n_312), .C(n_326), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_364), .B(n_313), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_348), .A2(n_305), .B1(n_327), .B2(n_319), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_354), .B(n_305), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_392), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_390), .B(n_347), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_391), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_390), .B(n_347), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_398), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_378), .B(n_377), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_392), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_399), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_383), .B(n_358), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx4_ASAP7_75t_R g415 ( .A(n_379), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_347), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_399), .B(n_367), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_383), .B(n_358), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_382), .B(n_347), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
INVx5_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_398), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_399), .B(n_370), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_395), .Y(n_434) );
CKINVDCx10_ASAP7_75t_R g435 ( .A(n_394), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_402), .B(n_370), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_402), .B(n_370), .Y(n_437) );
AND2x4_ASAP7_75t_SL g438 ( .A(n_398), .B(n_370), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_385), .B(n_367), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_413), .A2(n_396), .B(n_384), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_404), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_407), .B(n_385), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_436), .B(n_403), .Y(n_446) );
AOI322xp5_ASAP7_75t_L g447 ( .A1(n_421), .A2(n_388), .A3(n_381), .B1(n_360), .B2(n_356), .C1(n_357), .C2(n_389), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_416), .B(n_403), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_427), .B(n_398), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_436), .B(n_395), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_437), .B(n_395), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_414), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_437), .B(n_403), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_429), .B(n_394), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_427), .B(n_374), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_428), .B(n_374), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_394), .B1(n_380), .B2(n_397), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_414), .B(n_386), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_412), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_429), .B(n_386), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_410), .A2(n_397), .B1(n_368), .B2(n_375), .C(n_371), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_405), .A2(n_375), .B1(n_380), .B2(n_401), .Y(n_466) );
INVx5_ASAP7_75t_SL g467 ( .A(n_418), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_424), .A2(n_380), .B1(n_375), .B2(n_394), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_423), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_415), .Y(n_472) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_413), .A2(n_384), .B(n_371), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_430), .B(n_394), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_415), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_380), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_419), .A2(n_375), .B1(n_376), .B2(n_191), .C(n_350), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
AOI31xp33_ASAP7_75t_L g479 ( .A1(n_422), .A2(n_349), .A3(n_376), .B(n_350), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_412), .Y(n_480) );
NOR2xp67_ASAP7_75t_L g481 ( .A(n_425), .B(n_433), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_409), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g483 ( .A(n_425), .B(n_433), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_424), .B(n_386), .Y(n_485) );
INVx2_ASAP7_75t_R g486 ( .A(n_425), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx5_ASAP7_75t_L g489 ( .A(n_418), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_431), .B(n_386), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_380), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_471), .B(n_405), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_454), .B(n_408), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_489), .B(n_420), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_460), .A2(n_417), .B1(n_420), .B2(n_439), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_440), .B(n_408), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_440), .B(n_417), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_446), .B(n_439), .Y(n_498) );
NAND2xp33_ASAP7_75t_SL g499 ( .A(n_472), .B(n_435), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_451), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_451), .B(n_418), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_447), .B(n_432), .C(n_191), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_448), .B(n_434), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_445), .B(n_418), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_446), .B(n_434), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_452), .B(n_434), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_445), .B(n_432), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_468), .B(n_425), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_426), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_468), .B(n_433), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_479), .B(n_433), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_448), .B(n_409), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_465), .B(n_425), .C(n_433), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_476), .A2(n_433), .B1(n_438), .B2(n_409), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_453), .B(n_409), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_444), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_453), .B(n_409), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_485), .B(n_438), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_485), .B(n_438), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_444), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_458), .B(n_435), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_456), .B(n_409), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_459), .B(n_358), .Y(n_529) );
NAND2x1_ASAP7_75t_L g530 ( .A(n_472), .B(n_350), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_476), .B(n_358), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_463), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
OR2x4_ASAP7_75t_L g535 ( .A(n_475), .B(n_358), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_457), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_456), .B(n_358), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_489), .B(n_387), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_461), .B(n_365), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_489), .B(n_330), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_461), .B(n_365), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_469), .A2(n_362), .B1(n_387), .B2(n_353), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_352), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_464), .B(n_487), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_449), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_464), .B(n_352), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_489), .B(n_330), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_488), .B(n_352), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_541), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_498), .B(n_473), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_532), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_510), .B(n_474), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_498), .B(n_473), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_507), .B(n_491), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_547), .B(n_473), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_547), .B(n_488), .Y(n_560) );
NAND2x1_ASAP7_75t_L g561 ( .A(n_532), .B(n_484), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_494), .B(n_481), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_537), .B(n_490), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_533), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_515), .A2(n_467), .B1(n_483), .B2(n_466), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_537), .B(n_490), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_536), .B(n_450), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_508), .B(n_470), .Y(n_568) );
NAND2xp67_ASAP7_75t_L g569 ( .A(n_499), .B(n_470), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_496), .B(n_449), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_493), .B(n_455), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_529), .B(n_455), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_534), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_467), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_538), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_532), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_462), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_492), .B(n_462), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_509), .B(n_497), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_506), .B(n_491), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_521), .B(n_443), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_505), .A2(n_484), .B(n_477), .C(n_482), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_494), .B(n_484), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_500), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_521), .B(n_443), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_506), .B(n_467), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_499), .A2(n_515), .B(n_518), .C(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_504), .B(n_467), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_443), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_539), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_535), .B(n_482), .Y(n_591) );
AND5x1_ASAP7_75t_L g592 ( .A(n_535), .B(n_486), .C(n_68), .D(n_69), .E(n_70), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_531), .B(n_486), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_531), .B(n_362), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_517), .B(n_362), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_523), .B(n_61), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_520), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_528), .B(n_71), .Y(n_598) );
OR2x6_ASAP7_75t_L g599 ( .A(n_494), .B(n_319), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_500), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_501), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_528), .B(n_72), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_74), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_562), .B(n_519), .Y(n_604) );
AO22x1_ASAP7_75t_L g605 ( .A1(n_562), .A2(n_511), .B1(n_513), .B2(n_540), .Y(n_605) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_591), .A2(n_530), .B(n_546), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_576), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_564), .A2(n_495), .B1(n_524), .B2(n_525), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_553), .B(n_546), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_554), .A2(n_540), .B1(n_512), .B2(n_549), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_587), .A2(n_516), .B1(n_540), .B2(n_550), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_587), .A2(n_516), .B1(n_550), .B2(n_543), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_554), .A2(n_549), .B1(n_542), .B2(n_544), .Y(n_613) );
NAND2x1_ASAP7_75t_L g614 ( .A(n_562), .B(n_522), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_552), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_563), .B(n_522), .Y(n_616) );
BUFx2_ASAP7_75t_SL g617 ( .A(n_576), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_557), .A2(n_545), .B(n_551), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_551), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
AOI221x1_ASAP7_75t_SL g621 ( .A1(n_565), .A2(n_514), .B1(n_548), .B2(n_526), .C(n_501), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_566), .B(n_514), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_555), .A2(n_526), .B1(n_548), .B2(n_502), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_575), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_561), .A2(n_550), .B(n_543), .Y(n_626) );
NOR2xp67_ASAP7_75t_L g627 ( .A(n_583), .B(n_502), .Y(n_627) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_591), .A2(n_330), .B(n_248), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g629 ( .A1(n_593), .A2(n_276), .B(n_603), .C(n_588), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_579), .B(n_276), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_583), .A2(n_276), .B(n_582), .C(n_603), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_590), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_581), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_597), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_557), .B(n_276), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_560), .Y(n_636) );
NOR2xp67_ASAP7_75t_SL g637 ( .A(n_569), .B(n_602), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_558), .Y(n_638) );
OAI222xp33_ASAP7_75t_L g639 ( .A1(n_586), .A2(n_599), .B1(n_583), .B2(n_574), .C1(n_556), .C2(n_559), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_613), .B(n_585), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_611), .A2(n_599), .B(n_571), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_615), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_609), .B(n_589), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_607), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_614), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_633), .B(n_589), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_622), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_625), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_632), .Y(n_650) );
AOI21xp5_ASAP7_75t_SL g651 ( .A1(n_631), .A2(n_599), .B(n_596), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_616), .Y(n_652) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_604), .B(n_602), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_624), .B(n_601), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
OAI21xp33_ASAP7_75t_L g656 ( .A1(n_618), .A2(n_585), .B(n_581), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_612), .A2(n_599), .B(n_578), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
XOR2x2_ASAP7_75t_L g659 ( .A(n_605), .B(n_592), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_636), .B(n_568), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_620), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_639), .A2(n_596), .B(n_598), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_642), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_656), .A2(n_621), .B1(n_633), .B2(n_639), .C(n_638), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_644), .A2(n_620), .B(n_629), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_644), .A2(n_637), .B(n_608), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_662), .A2(n_653), .B1(n_659), .B2(n_640), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_653), .A2(n_654), .B1(n_657), .B2(n_641), .C(n_646), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_648), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_654), .A2(n_606), .B(n_608), .C(n_628), .Y(n_670) );
NOR2x1_ASAP7_75t_SL g671 ( .A(n_661), .B(n_598), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_651), .A2(n_610), .B1(n_627), .B2(n_624), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_659), .A2(n_626), .B(n_619), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_570), .B(n_572), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_658), .B(n_568), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_663), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_669), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_675), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_674), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_665), .Y(n_680) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_667), .A2(n_661), .A3(n_650), .B1(n_655), .B2(n_649), .C1(n_652), .C2(n_643), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_668), .A2(n_647), .B1(n_660), .B2(n_567), .Y(n_682) );
AOI22xp5_ASAP7_75t_SL g683 ( .A1(n_672), .A2(n_577), .B1(n_635), .B2(n_594), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_680), .A2(n_673), .B1(n_664), .B2(n_666), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_679), .Y(n_685) );
OAI222xp33_ASAP7_75t_R g686 ( .A1(n_682), .A2(n_670), .B1(n_671), .B2(n_584), .C1(n_600), .C2(n_601), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_678), .B(n_580), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_685), .B(n_683), .C(n_677), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_687), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_684), .B(n_676), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_689), .Y(n_691) );
NOR4xp25_ASAP7_75t_SL g692 ( .A(n_690), .B(n_686), .C(n_681), .D(n_677), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_688), .B1(n_677), .B2(n_630), .Y(n_693) );
BUFx3_ASAP7_75t_L g694 ( .A(n_693), .Y(n_694) );
AOI32xp33_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_691), .A3(n_577), .B1(n_595), .B2(n_600), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_694), .B(n_584), .Y(n_697) );
endmodule