module fake_jpeg_12195_n_480 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_480);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_480;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_58),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_59),
.B(n_64),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

BUFx2_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_94),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_25),
.B(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_77),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_73),
.B(n_75),
.Y(n_176)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_12),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_80),
.Y(n_195)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_12),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_93),
.Y(n_137)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_88),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_40),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_11),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_100),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_33),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_111),
.Y(n_153)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_34),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_109),
.B(n_114),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_34),
.B(n_8),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_19),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_44),
.B(n_8),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_119),
.Y(n_160)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_52),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_21),
.B1(n_51),
.B2(n_54),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_123),
.A2(n_126),
.B1(n_135),
.B2(n_148),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_42),
.B(n_56),
.C(n_31),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_124),
.A2(n_170),
.B(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_48),
.B1(n_55),
.B2(n_51),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_125),
.A2(n_128),
.B1(n_48),
.B2(n_55),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_21),
.B1(n_54),
.B2(n_57),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_48),
.B1(n_55),
.B2(n_24),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_128),
.A2(n_168),
.B1(n_187),
.B2(n_192),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_57),
.B1(n_24),
.B2(n_36),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_36),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_159),
.C(n_172),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_36),
.B1(n_24),
.B2(n_39),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_48),
.B1(n_55),
.B2(n_47),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_151),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_31),
.B1(n_47),
.B2(n_42),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_154),
.A2(n_186),
.B1(n_190),
.B2(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_56),
.C(n_44),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_52),
.B1(n_30),
.B2(n_37),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_165),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_68),
.A2(n_37),
.B(n_30),
.C(n_3),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_0),
.B(n_2),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_86),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_80),
.A2(n_7),
.B(n_120),
.C(n_112),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_98),
.A2(n_95),
.B1(n_83),
.B2(n_81),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_178),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_91),
.B(n_101),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_92),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_172),
.C(n_180),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_58),
.A2(n_28),
.B1(n_21),
.B2(n_46),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_58),
.A2(n_28),
.B1(n_21),
.B2(n_46),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_69),
.A2(n_28),
.B1(n_21),
.B2(n_46),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_69),
.A2(n_67),
.B1(n_84),
.B2(n_105),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_96),
.A2(n_67),
.B1(n_92),
.B2(n_104),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_93),
.A2(n_82),
.B(n_75),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_93),
.B(n_94),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_139),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_204),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_248),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_125),
.A2(n_141),
.B1(n_144),
.B2(n_175),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_199),
.A2(n_231),
.B1(n_238),
.B2(n_249),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_200),
.Y(n_298)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_202),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_124),
.Y(n_204)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_SL g210 ( 
.A(n_137),
.B(n_159),
.C(n_160),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_210),
.B(n_223),
.Y(n_294)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_212),
.B(n_215),
.Y(n_265)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_133),
.B(n_153),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_137),
.B(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_217),
.B(n_228),
.Y(n_287)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_232),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_147),
.Y(n_220)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g221 ( 
.A(n_143),
.Y(n_221)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_222),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_129),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_142),
.B(n_127),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_225),
.B(n_234),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_239),
.C(n_203),
.Y(n_285)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_129),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_141),
.A2(n_144),
.B1(n_161),
.B2(n_175),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_169),
.C(n_157),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_176),
.B(n_149),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_236),
.B(n_237),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_131),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_134),
.C(n_166),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_134),
.B(n_156),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_241),
.B(n_246),
.Y(n_299)
);

OR2x2_ASAP7_75t_SL g242 ( 
.A(n_157),
.B(n_169),
.Y(n_242)
);

OR2x2_ASAP7_75t_SL g295 ( 
.A(n_242),
.B(n_223),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_260),
.B1(n_171),
.B2(n_150),
.Y(n_263)
);

INVx4_ASAP7_75t_SL g244 ( 
.A(n_162),
.Y(n_244)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_122),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_162),
.Y(n_247)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_122),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_168),
.A2(n_187),
.B1(n_138),
.B2(n_152),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_154),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_152),
.B(n_163),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_140),
.B(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_242),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_121),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_258),
.Y(n_289)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_121),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_163),
.B(n_140),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_207),
.A2(n_150),
.B(n_171),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_208),
.B(n_300),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_275),
.B1(n_260),
.B2(n_209),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_210),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_277),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_243),
.B1(n_228),
.B2(n_204),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_301),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_217),
.B(n_197),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_226),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_232),
.B(n_229),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_293),
.B(n_296),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_244),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_205),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_303),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_205),
.B(n_258),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_211),
.B(n_216),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_196),
.B(n_220),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_200),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_306),
.B(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_308),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_238),
.B1(n_254),
.B2(n_233),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_310),
.B(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_247),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_317),
.C(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_245),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_318),
.A2(n_283),
.B(n_299),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_263),
.A2(n_206),
.B1(n_218),
.B2(n_222),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_333),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_202),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_268),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_328),
.Y(n_372)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_213),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_331),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_227),
.B1(n_202),
.B2(n_235),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_330),
.A2(n_332),
.B1(n_276),
.B2(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_202),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_287),
.A2(n_221),
.B1(n_266),
.B2(n_269),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_221),
.B1(n_288),
.B2(n_271),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_267),
.B(n_281),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_336),
.B(n_337),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_270),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_341),
.Y(n_367)
);

OAI22x1_ASAP7_75t_L g340 ( 
.A1(n_274),
.A2(n_295),
.B1(n_278),
.B2(n_271),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_340),
.A2(n_272),
.B(n_297),
.C(n_302),
.Y(n_365)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_343),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_R g391 ( 
.A(n_346),
.B(n_320),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_306),
.B(n_318),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_333),
.A2(n_266),
.B(n_278),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_364),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_313),
.B1(n_312),
.B2(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_319),
.A2(n_307),
.B1(n_308),
.B2(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_276),
.C(n_304),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_362),
.C(n_335),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_304),
.C(n_302),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_311),
.A2(n_269),
.B(n_297),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_365),
.A2(n_366),
.B(n_334),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_298),
.B(n_272),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_273),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_355),
.Y(n_381)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_378),
.C(n_386),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_340),
.C(n_315),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_366),
.B(n_356),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_361),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_383),
.Y(n_401)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_348),
.Y(n_382)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_361),
.B(n_314),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_384),
.B(n_391),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_387),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_360),
.C(n_352),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_341),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_388),
.Y(n_397)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_392),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_339),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_324),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_394),
.C(n_346),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_362),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_309),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_395),
.A2(n_344),
.B(n_358),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_359),
.B(n_342),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_372),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_402),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_372),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_404),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_359),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_364),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_414),
.C(n_417),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_409),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_353),
.B(n_365),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_415),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_365),
.C(n_353),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_369),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_371),
.Y(n_418)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

A2O1A1O1Ixp25_ASAP7_75t_L g420 ( 
.A1(n_400),
.A2(n_374),
.B(n_381),
.C(n_390),
.D(n_391),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_404),
.Y(n_442)
);

BUFx4f_ASAP7_75t_SL g422 ( 
.A(n_415),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_424),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_416),
.Y(n_424)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_427),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_412),
.A2(n_390),
.B1(n_347),
.B2(n_382),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_411),
.B1(n_408),
.B2(n_405),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_396),
.C(n_390),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_431),
.C(n_403),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_401),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_432),
.B1(n_410),
.B2(n_409),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_395),
.C(n_385),
.Y(n_431)
);

AO22x1_ASAP7_75t_SL g432 ( 
.A1(n_412),
.A2(n_379),
.B1(n_365),
.B2(n_387),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_417),
.B(n_371),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_433),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_406),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_435),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_397),
.B1(n_413),
.B2(n_414),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_413),
.B1(n_398),
.B2(n_408),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_441),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_446),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_421),
.C(n_426),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_428),
.A2(n_351),
.B1(n_405),
.B2(n_388),
.Y(n_444)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_423),
.A2(n_392),
.B1(n_351),
.B2(n_402),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_395),
.B(n_432),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_450),
.B(n_422),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_441),
.A2(n_420),
.B(n_432),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_454),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_SL g454 ( 
.A(n_440),
.B(n_365),
.C(n_429),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_431),
.C(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_419),
.C(n_442),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_449),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_461),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_434),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_463),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_460),
.B(n_462),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_419),
.C(n_437),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_452),
.B(n_446),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_427),
.Y(n_464)
);

NOR4xp25_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_454),
.C(n_422),
.D(n_455),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_458),
.A2(n_453),
.B1(n_447),
.B2(n_450),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_467),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_455),
.C(n_451),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g471 ( 
.A1(n_468),
.A2(n_469),
.A3(n_465),
.B1(n_445),
.B2(n_464),
.C1(n_470),
.C2(n_467),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_472),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_459),
.C(n_383),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_343),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_473),
.B(n_325),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_475),
.B(n_474),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_478),
.C(n_370),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_476),
.A2(n_370),
.B(n_363),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_357),
.Y(n_480)
);


endmodule