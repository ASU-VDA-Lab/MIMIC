module fake_jpeg_30260_n_544 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_544);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_58),
.Y(n_115)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_60),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_17),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_24),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_94),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_0),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_102),
.Y(n_151)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_96),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_99),
.Y(n_137)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_22),
.Y(n_158)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_158),
.Y(n_173)
);

BUFx12f_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_121),
.Y(n_178)
);

CKINVDCx9p33_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_122),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_40),
.B1(n_26),
.B2(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_129),
.A2(n_100),
.B1(n_88),
.B2(n_67),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_22),
.B(n_39),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_135),
.B(n_154),
.C(n_25),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_150),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_144),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_70),
.B(n_27),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_44),
.B(n_52),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_152),
.B(n_164),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_99),
.A2(n_22),
.B(n_52),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_101),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_93),
.B(n_24),
.Y(n_164)
);

BUFx16f_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_68),
.B1(n_54),
.B2(n_65),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_129),
.B1(n_160),
.B2(n_165),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_174),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_119),
.A2(n_97),
.B1(n_86),
.B2(n_104),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_210),
.B1(n_221),
.B2(n_226),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_186),
.Y(n_264)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_49),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_196),
.Y(n_232)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_74),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_143),
.C(n_132),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_116),
.B(n_47),
.Y(n_196)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_47),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_204),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_49),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_46),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_207),
.B(n_208),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_46),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_119),
.A2(n_69),
.B1(n_56),
.B2(n_82),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_149),
.A2(n_105),
.B1(n_66),
.B2(n_71),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_213),
.A2(n_161),
.B1(n_156),
.B2(n_136),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_37),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_214),
.B(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_124),
.B(n_37),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_118),
.B(n_30),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_30),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_223),
.Y(n_250)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_225),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_224),
.B1(n_73),
.B2(n_72),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_137),
.B(n_44),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_149),
.A2(n_85),
.B1(n_81),
.B2(n_75),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_28),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_178),
.A2(n_163),
.B1(n_159),
.B2(n_145),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_236),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_178),
.A2(n_159),
.B1(n_112),
.B2(n_165),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_238),
.A2(n_241),
.B1(n_248),
.B2(n_254),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_175),
.A2(n_112),
.B1(n_155),
.B2(n_131),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_266),
.B1(n_221),
.B2(n_233),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_131),
.B1(n_140),
.B2(n_160),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_192),
.A2(n_140),
.B1(n_50),
.B2(n_45),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_26),
.A3(n_51),
.B1(n_40),
.B2(n_25),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_271),
.B1(n_182),
.B2(n_190),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_193),
.A2(n_167),
.B1(n_132),
.B2(n_156),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_266),
.A2(n_269),
.B1(n_171),
.B2(n_197),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_170),
.A2(n_51),
.B1(n_167),
.B2(n_50),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_172),
.A2(n_173),
.B1(n_170),
.B2(n_195),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_184),
.A2(n_45),
.B1(n_161),
.B2(n_36),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_217),
.B1(n_176),
.B2(n_197),
.Y(n_298)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_276),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_195),
.B(n_209),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_283),
.B(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_168),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_280),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_206),
.Y(n_280)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_179),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_292),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_198),
.B(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_286),
.A2(n_298),
.B1(n_272),
.B2(n_268),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_289),
.B1(n_305),
.B2(n_262),
.Y(n_318)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_246),
.A2(n_185),
.B1(n_213),
.B2(n_212),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_237),
.A2(n_225),
.B(n_198),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_290),
.B(n_272),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_217),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_259),
.B(n_36),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_299),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_36),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_232),
.B(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_301),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_144),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_251),
.B(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_308),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_247),
.B(n_169),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_SL g346 ( 
.A(n_303),
.B(n_153),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_230),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_304),
.B(n_310),
.Y(n_339)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_205),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_311),
.B(n_315),
.Y(n_352)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.Y(n_321)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

BUFx16f_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_316),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_199),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_176),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_171),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_318),
.A2(n_322),
.B1(n_323),
.B2(n_334),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_269),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_320),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_233),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_233),
.B1(n_243),
.B2(n_235),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_228),
.B1(n_245),
.B2(n_264),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_267),
.C(n_245),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_332),
.C(n_336),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_278),
.C(n_277),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_305),
.A2(n_228),
.B1(n_263),
.B2(n_234),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_268),
.C(n_263),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_337),
.A2(n_302),
.B(n_290),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_338),
.A2(n_341),
.B1(n_344),
.B2(n_347),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_242),
.B1(n_258),
.B2(n_253),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_282),
.B(n_153),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_284),
.C(n_293),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_286),
.A2(n_301),
.B1(n_283),
.B2(n_275),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_292),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_242),
.B1(n_258),
.B2(n_253),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_153),
.C(n_239),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_317),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_291),
.A2(n_239),
.B1(n_234),
.B2(n_260),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_313),
.B1(n_307),
.B2(n_265),
.Y(n_385)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_308),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_359),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_360),
.A2(n_367),
.B(n_323),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_340),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_316),
.B(n_312),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_345),
.B(n_300),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_368),
.B(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_315),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_374),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_353),
.A2(n_288),
.B1(n_285),
.B2(n_304),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_375),
.A2(n_351),
.B1(n_354),
.B2(n_325),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_376),
.B(n_378),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_318),
.A2(n_289),
.B1(n_295),
.B2(n_309),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_337),
.B1(n_320),
.B2(n_343),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_345),
.B(n_294),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_265),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_379),
.B(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_329),
.B(n_331),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_311),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_310),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_388),
.C(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_386),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_389),
.B1(n_334),
.B2(n_351),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_329),
.B(n_314),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_314),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_390),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_314),
.C(n_281),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_319),
.A2(n_281),
.B1(n_276),
.B2(n_306),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g390 ( 
.A(n_324),
.B(n_306),
.CI(n_276),
.CON(n_390),
.SN(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_1),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_400),
.B1(n_410),
.B2(n_421),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_403),
.C(n_418),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_364),
.A2(n_346),
.B1(n_322),
.B2(n_337),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_333),
.C(n_335),
.Y(n_403)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_326),
.C(n_333),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_404),
.B(n_411),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_372),
.B1(n_364),
.B2(n_377),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_350),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_417),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_365),
.B(n_325),
.CI(n_321),
.CON(n_411),
.SN(n_411)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_365),
.A2(n_340),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_413)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_1),
.Y(n_416)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_416),
.Y(n_430)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_53),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_53),
.C(n_43),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_1),
.Y(n_420)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_372),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_390),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_446),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_400),
.B1(n_405),
.B2(n_406),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_388),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_438),
.Y(n_454)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_418),
.Y(n_452)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_436),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_390),
.C(n_360),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_440),
.C(n_442),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_389),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_384),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_439),
.B(n_441),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_380),
.C(n_373),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_393),
.B(n_358),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_385),
.C(n_391),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_371),
.C(n_362),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_445),
.C(n_394),
.Y(n_455)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_422),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_362),
.C(n_53),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_412),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_53),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_411),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_455),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_453),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_456),
.B(n_465),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_423),
.C(n_396),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_460),
.C(n_464),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_431),
.B(n_408),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_458),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_412),
.C(n_396),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_461),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_425),
.A2(n_449),
.B1(n_430),
.B2(n_429),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_466),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_394),
.C(n_398),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_413),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_448),
.A2(n_421),
.B1(n_398),
.B2(n_407),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_407),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_469),
.C(n_471),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_53),
.C(n_43),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_5),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_470),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_43),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_448),
.B1(n_437),
.B2(n_445),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_475),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_433),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_460),
.A2(n_424),
.B(n_444),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_485),
.B(n_491),
.Y(n_504)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_487),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_435),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_479),
.B(n_12),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_426),
.C(n_450),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_454),
.C(n_468),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_456),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_10),
.B(n_11),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_464),
.A2(n_10),
.B(n_11),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_475),
.A2(n_455),
.B(n_451),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_490),
.B(n_480),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_457),
.Y(n_493)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_502),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_497),
.B(n_482),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_469),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_501),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_454),
.C(n_471),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_500),
.C(n_503),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_43),
.C(n_13),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_475),
.B(n_12),
.CI(n_13),
.CON(n_502),
.SN(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_43),
.C(n_13),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_12),
.C(n_13),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_491),
.C(n_478),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_14),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_506),
.A2(n_485),
.B(n_481),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g507 ( 
.A(n_481),
.B(n_15),
.CI(n_487),
.CON(n_507),
.SN(n_507)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_15),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_497),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_517),
.C(n_494),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_510),
.B(n_512),
.Y(n_529)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_513),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_480),
.C(n_484),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_486),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_518),
.B(n_505),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_500),
.B(n_15),
.Y(n_519)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_519),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_502),
.Y(n_523)
);

OA21x2_ASAP7_75t_SL g521 ( 
.A1(n_516),
.A2(n_499),
.B(n_507),
.Y(n_521)
);

CKINVDCx14_ASAP7_75t_R g533 ( 
.A(n_521),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_522),
.B(n_524),
.Y(n_534)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_523),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_509),
.A2(n_504),
.B(n_496),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_522),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_529),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_531),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_525),
.B(n_527),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_537),
.B(n_508),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_SL g540 ( 
.A(n_538),
.B(n_539),
.Y(n_540)
);

AOI322xp5_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_532),
.A3(n_533),
.B1(n_524),
.B2(n_515),
.C1(n_528),
.C2(n_517),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_504),
.B(n_523),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_511),
.B(n_512),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_507),
.B(n_502),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_543),
.A2(n_520),
.B(n_15),
.Y(n_544)
);


endmodule