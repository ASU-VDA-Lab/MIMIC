module real_jpeg_12798_n_17 (n_5, n_4, n_8, n_0, n_12, n_274, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_274;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx10_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_39),
.B1(n_63),
.B2(n_65),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_31),
.B1(n_34),
.B2(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_57),
.B1(n_63),
.B2(n_65),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_49),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_31),
.B1(n_34),
.B2(n_49),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_6),
.A2(n_49),
.B1(n_63),
.B2(n_65),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_70),
.Y(n_110)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_140),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_10),
.A2(n_33),
.B(n_34),
.C(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_10),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_10),
.B(n_45),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_154),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_10),
.B(n_63),
.C(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_10),
.B(n_35),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_10),
.A2(n_66),
.B(n_200),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_31),
.B1(n_34),
.B2(n_154),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_31),
.B1(n_34),
.B2(n_81),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_31),
.B1(n_34),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_12),
.B(n_31),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_13),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_31),
.B1(n_34),
.B2(n_100),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_100),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_13),
.A2(n_63),
.B1(n_65),
.B2(n_100),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_62),
.Y(n_90)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_16),
.A2(n_31),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_16),
.A2(n_42),
.B1(n_63),
.B2(n_65),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_104),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_21),
.B(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_84),
.C(n_92),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_22),
.A2(n_23),
.B1(n_84),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_83),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_43),
.C(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_27),
.A2(n_40),
.B1(n_41),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_27),
.A2(n_40),
.B1(n_136),
.B2(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_27),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_27),
.A2(n_167),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_30),
.A2(n_36),
.B(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_34),
.A2(n_46),
.A3(n_52),
.B1(n_164),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_35),
.B(n_103),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_37),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_37),
.B(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_38),
.A2(n_40),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_40),
.A2(n_102),
.B(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B(n_54),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_44),
.A2(n_50),
.B1(n_51),
.B2(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_46),
.A2(n_50),
.B(n_154),
.C(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_51),
.A2(n_99),
.B(n_121),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_55),
.B(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_72),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_59),
.A2(n_72),
.B1(n_73),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_59),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_65),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_66),
.A2(n_71),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_66),
.A2(n_71),
.B1(n_144),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_66),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_68),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_67),
.A2(n_68),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_68),
.B(n_157),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_143),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_71),
.A2(n_156),
.B(n_205),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_71),
.B(n_154),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_80),
.B1(n_82),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_75),
.B(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_75),
.A2(n_82),
.B1(n_147),
.B2(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_90),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_79),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_79),
.A2(n_170),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_79),
.B(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_84),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_86),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_91),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_92),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.C(n_101),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_93),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_94),
.B(n_96),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_95),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_97),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_98),
.B(n_101),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_126),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_114),
.B2(n_115),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_113),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_111),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_109),
.A2(n_148),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_267),
.B(n_272),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_241),
.A3(n_260),
.B1(n_265),
.B2(n_266),
.C(n_274),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_181),
.B(n_240),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_158),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_132),
.B(n_158),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_145),
.C(n_150),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_133),
.A2(n_134),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_138),
.C(n_142),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_145),
.A2(n_150),
.B1(n_151),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_152),
.B(n_155),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_172),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_159),
.B(n_173),
.C(n_174),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_165),
.B2(n_171),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_160),
.B(n_166),
.C(n_168),
.Y(n_252)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_179),
.Y(n_250)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_233),
.B(n_239),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_220),
.B(n_232),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_201),
.B(n_219),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_196),
.C(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_199),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_209),
.B(n_218),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_207),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_213),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_228),
.C(n_231),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_253),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_253),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.C(n_252),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_244),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_252),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.C(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_271),
.Y(n_272)
);


endmodule