module real_jpeg_1793_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_295;
wire n_213;
wire n_128;
wire n_179;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_0),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_0),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_35),
.B1(n_37),
.B2(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_2),
.A2(n_45),
.B1(n_49),
.B2(n_60),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_3),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_94),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_94),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_94),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_131),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_131),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_45),
.B1(n_49),
.B2(n_131),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_6),
.B(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_6),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_6),
.A2(n_26),
.B(n_166),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_63),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_37),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_45),
.C(n_48),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_202),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_6),
.B(n_85),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_6),
.B(n_43),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_28),
.B1(n_52),
.B2(n_53),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_28),
.B1(n_45),
.B2(n_49),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_176),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_176),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_45),
.B1(n_49),
.B2(n_176),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_156),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_156),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_14),
.A2(n_45),
.B1(n_49),
.B2(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_16),
.A2(n_35),
.B1(n_37),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_16),
.A2(n_45),
.B1(n_49),
.B2(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_95),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_21),
.B(n_95),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_78),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_22),
.A2(n_71),
.B1(n_72),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_22),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_23),
.A2(n_24),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_42),
.C(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_25),
.A2(n_29),
.B1(n_34),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_33),
.A3(n_37),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_29),
.A2(n_34),
.B1(n_93),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_29),
.A2(n_34),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_29),
.A2(n_34),
.B1(n_175),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_30),
.A2(n_130),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_32),
.B(n_35),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_34),
.Y(n_157)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_35),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_37),
.A2(n_53),
.A3(n_64),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_70),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_50),
.B(n_55),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_50),
.B1(n_55),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_50),
.B1(n_77),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_43),
.A2(n_50),
.B1(n_90),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_43),
.A2(n_50),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_43),
.A2(n_50),
.B1(n_198),
.B2(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_43),
.A2(n_50),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_43),
.A2(n_50),
.B1(n_225),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_44),
.A2(n_124),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_44),
.A2(n_149),
.B1(n_197),
.B2(n_237),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_45),
.B(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_50),
.Y(n_149)
);

AO22x2_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_52),
.B(n_65),
.Y(n_203)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_53),
.B(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_67),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_63),
.B1(n_127),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_68),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_62),
.A2(n_75),
.B1(n_102),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_62),
.A2(n_102),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_62),
.A2(n_102),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_62),
.A2(n_102),
.B1(n_172),
.B2(n_188),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_62),
.A2(n_102),
.B1(n_187),
.B2(n_234),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_78),
.B(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_91),
.B(n_92),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_79),
.A2(n_80),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_91),
.B1(n_92),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_86),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_84),
.B1(n_120),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_82),
.A2(n_84),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_82),
.A2(n_84),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_83),
.A2(n_85),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_83),
.A2(n_85),
.B1(n_169),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_83),
.A2(n_85),
.B1(n_206),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_83),
.A2(n_85),
.B1(n_202),
.B2(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_83),
.A2(n_85),
.B1(n_255),
.B2(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_292),
.B(n_297),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_158),
.B(n_291),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_140),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_140),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_132),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_114),
.B(n_134),
.C(n_139),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.C(n_128),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_116),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_139),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_145),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.C(n_154),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_147),
.B(n_150),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_154),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_181),
.B(n_290),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_179),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_160),
.B(n_179),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_178),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_161),
.B(n_178),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_163),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.C(n_174),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_164),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_171),
.B(n_174),
.Y(n_281)
);

AOI31xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_275),
.A3(n_284),
.B(n_287),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_220),
.B(n_274),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_208),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_184),
.B(n_208),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.C(n_199),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_190),
.C(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_195),
.B(n_199),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_208),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_208),
.B(n_285),
.Y(n_288)
);

FAx1_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.CI(n_211),
.CON(n_208),
.SN(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_215),
.C(n_219),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_269),
.B(n_273),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_238),
.B(n_268),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_230),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_227),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_233),
.C(n_236),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_249),
.B(n_267),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_261),
.B(n_266),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_260),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_258),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_272),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_296),
.Y(n_297)
);


endmodule