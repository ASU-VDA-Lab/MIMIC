module real_jpeg_17090_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_2),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_2),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_3),
.B(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_3),
.B(n_29),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_3),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_3),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_126),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_4),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_4),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_4),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_5),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_5),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_5),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_5),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_5),
.B(n_135),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_8),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_8),
.B(n_105),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_8),
.B(n_181),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_8),
.B(n_257),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_10),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_10),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_10),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_10),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_10),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_11),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_11),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_11),
.B(n_316),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_12),
.Y(n_321)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_13),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_15),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_68),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_15),
.B(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_16),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_111),
.B(n_343),
.C(n_410),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_24),
.A2(n_25),
.B1(n_62),
.B2(n_70),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.C(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_26),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_56),
.C(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_26),
.A2(n_49),
.B1(n_58),
.B2(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_26),
.B(n_189),
.C(n_194),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_26),
.A2(n_49),
.B1(n_189),
.B2(n_190),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_27),
.B(n_130),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_27),
.B(n_146),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_27),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_30),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_67),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_31),
.B(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_32),
.A2(n_33),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_33),
.B(n_168),
.C(n_171),
.Y(n_207)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_36),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

XNOR2x1_ASAP7_75t_SL g358 ( 
.A(n_37),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_71),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_43),
.B(n_71),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_61),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.C(n_55),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_46),
.B(n_194),
.C(n_362),
.Y(n_373)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g74 ( 
.A(n_55),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_101),
.C(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_58),
.B(n_162),
.C(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_58),
.A2(n_101),
.B1(n_110),
.B2(n_311),
.Y(n_371)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_63),
.A2(n_64),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_77),
.C(n_83),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_64),
.B(n_69),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_67),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_67),
.B(n_186),
.C(n_218),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.C(n_96),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_72),
.B(n_75),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.C(n_92),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_98),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_78),
.B(n_83),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_82),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_83),
.A2(n_84),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_83),
.B(n_199),
.C(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_93),
.A2(n_99),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_93),
.A2(n_99),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_95),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_96),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_108),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_97),
.B(n_368),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_99),
.B(n_209),
.C(n_212),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_99),
.B(n_343),
.C(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_100),
.B(n_108),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_101),
.B(n_251),
.C(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_101),
.A2(n_251),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_101),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_101),
.A2(n_217),
.B1(n_218),
.B2(n_311),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_SL g372 ( 
.A(n_101),
.B(n_218),
.C(n_350),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_104),
.B(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_110),
.B(n_278),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_364),
.B(n_404),
.C(n_409),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_270),
.B(n_325),
.C(n_326),
.D(n_363),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_237),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_115),
.B(n_237),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_175),
.Y(n_115)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_116),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_152),
.C(n_166),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_118),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_131),
.C(n_141),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_119),
.B(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_125),
.C(n_129),
.Y(n_168)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_122),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_131),
.A2(n_132),
.B1(n_141),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_132),
.A2(n_133),
.B(n_138),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_141),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.C(n_147),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_142),
.B(n_143),
.Y(n_245)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_147),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_152),
.A2(n_166),
.B1(n_167),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_152),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_161),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_153),
.B(n_157),
.Y(n_262)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_161),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_162),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_164),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_214),
.B1(n_235),
.B2(n_236),
.Y(n_175)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_205),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_177),
.B(n_206),
.C(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.C(n_198),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_188),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_185),
.B(n_186),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_184),
.A2(n_185),
.B1(n_248),
.B2(n_249),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_186),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_187),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_193),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_194),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_194),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_194),
.A2(n_266),
.B1(n_360),
.B2(n_362),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2x1_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_269),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_213),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_213),
.Y(n_334)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_214),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_215),
.B(n_220),
.C(n_223),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_229),
.B1(n_233),
.B2(n_234),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_229),
.B(n_234),
.C(n_278),
.Y(n_357)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.C(n_267),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_238),
.A2(n_239),
.B1(n_268),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_261),
.C(n_263),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.C(n_250),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_244),
.B(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_254),
.Y(n_361)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_256),
.B(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_296),
.B(n_324),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_293),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.C(n_290),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_280)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.C(n_307),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.C(n_313),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.C(n_322),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_332),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.C(n_331),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_R g386 ( 
.A(n_333),
.B(n_336),
.C(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_347),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_339),
.C(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_343),
.Y(n_346)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_356),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_357),
.C(n_358),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_385),
.C(n_399),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_365),
.A2(n_405),
.B(n_408),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_383),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_383),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.C(n_374),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_369),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_373),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.C(n_381),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_386),
.B(n_388),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_397),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_393),
.B2(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_393),
.C(n_397),
.Y(n_403)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_400),
.A2(n_406),
.B(n_407),
.Y(n_405)
);

NOR2x1_ASAP7_75t_R g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_403),
.Y(n_407)
);


endmodule