module fake_netlist_6_2107_n_149 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_149);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_149;

wire n_52;
wire n_119;
wire n_91;
wire n_46;
wire n_146;
wire n_147;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_48),
.Y(n_55)
);

OR2x6_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_5),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_9),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_13),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_42),
.B(n_40),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_50),
.B(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_40),
.B1(n_18),
.B2(n_20),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_14),
.B(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_69),
.B(n_70),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_70),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_67),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_59),
.B(n_74),
.C(n_65),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_58),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_61),
.B(n_56),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_74),
.B1(n_56),
.B2(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_68),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_61),
.B(n_56),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_67),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

AO21x2_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_76),
.B(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AO21x2_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_92),
.B(n_95),
.Y(n_105)
);

NAND4xp25_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_75),
.C(n_86),
.D(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_94),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_73),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_98),
.C(n_93),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_73),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_110),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_103),
.B(n_115),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_118),
.Y(n_126)
);

NOR2x1_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_117),
.B1(n_118),
.B2(n_61),
.C(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_91),
.B1(n_104),
.B2(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_64),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_64),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_64),
.Y(n_141)
);

AND2x4_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_64),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_140),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_146),
.B1(n_141),
.B2(n_142),
.C(n_143),
.Y(n_149)
);


endmodule