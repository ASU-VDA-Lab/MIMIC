module fake_jpeg_27256_n_296 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_36),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_58),
.B1(n_62),
.B2(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_34),
.B1(n_36),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_26),
.B1(n_25),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_34),
.B1(n_26),
.B2(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_35),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_63),
.A2(n_93),
.B1(n_101),
.B2(n_21),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_68),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_76),
.B(n_78),
.C(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_18),
.B(n_33),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_88),
.B(n_0),
.Y(n_108)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_29),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_85),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_81),
.Y(n_125)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_28),
.B1(n_45),
.B2(n_24),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_84),
.B1(n_98),
.B2(n_17),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_22),
.B(n_38),
.C(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_94),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

OR2x4_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_19),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_32),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_92),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_21),
.C(n_24),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_25),
.B1(n_27),
.B2(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_27),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_27),
.B1(n_17),
.B2(n_19),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_116),
.B1(n_84),
.B2(n_78),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_127),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_114),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_21),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_31),
.B1(n_29),
.B2(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_75),
.B1(n_103),
.B2(n_88),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_0),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_132),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_1),
.B(n_2),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_126),
.B(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_79),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_93),
.C(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_149),
.C(n_124),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_124),
.B1(n_109),
.B2(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_74),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_148),
.B1(n_158),
.B2(n_113),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_76),
.B1(n_78),
.B2(n_73),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_87),
.C(n_76),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_86),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_114),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_82),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_89),
.B1(n_85),
.B2(n_83),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_R g159 ( 
.A(n_112),
.B(n_132),
.Y(n_159)
);

XOR2x1_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_127),
.Y(n_165)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_167),
.B1(n_187),
.B2(n_190),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_122),
.B(n_129),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_129),
.B(n_132),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_175),
.B(n_180),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_184),
.C(n_160),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_118),
.B(n_117),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_133),
.C(n_131),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_104),
.B(n_106),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_104),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_156),
.B1(n_91),
.B2(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_106),
.B(n_120),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_148),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_211),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_149),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_186),
.B(n_178),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_138),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_200),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_202),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_203),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_130),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_171),
.B1(n_8),
.B2(n_10),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_213),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_179),
.C(n_175),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_140),
.A3(n_147),
.B1(n_97),
.B2(n_91),
.C1(n_81),
.C2(n_86),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_215),
.B1(n_178),
.B2(n_173),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_201),
.B1(n_162),
.B2(n_192),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_219),
.B1(n_222),
.B2(n_205),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_206),
.A2(n_184),
.B1(n_168),
.B2(n_185),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_224),
.C(n_232),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_188),
.B1(n_172),
.B2(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_182),
.C(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_214),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_228),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_215),
.B1(n_209),
.B2(n_196),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_6),
.C(n_10),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_16),
.C(n_11),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_238),
.A2(n_242),
.B1(n_221),
.B2(n_212),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_207),
.B(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_248),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_247),
.B1(n_225),
.B2(n_199),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_245),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_207),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_252),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_203),
.B1(n_212),
.B2(n_196),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_219),
.C(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_235),
.B1(n_231),
.B2(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_222),
.C(n_193),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_225),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_238),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_273),
.B(n_258),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_252),
.B(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_260),
.C(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_261),
.Y(n_281)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_274),
.Y(n_285)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_251),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_289),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_283),
.B(n_282),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_284),
.B(n_286),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_291),
.B(n_284),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_278),
.B(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_294),
.B(n_256),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_256),
.Y(n_296)
);


endmodule