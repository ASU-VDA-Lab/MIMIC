module fake_jpeg_22685_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_24),
.B1(n_19),
.B2(n_32),
.Y(n_54)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_35),
.B1(n_41),
.B2(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_62),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_85),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_84),
.B1(n_80),
.B2(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_82),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_40),
.B1(n_41),
.B2(n_19),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_39),
.B1(n_37),
.B2(n_53),
.Y(n_107)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_75),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_37),
.B1(n_19),
.B2(n_33),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_79),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_38),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_84),
.B(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_40),
.B(n_39),
.C(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_103),
.B1(n_107),
.B2(n_77),
.Y(n_123)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_39),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_53),
.B(n_58),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_38),
.C(n_33),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_46),
.C(n_69),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_39),
.B1(n_33),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_77),
.B1(n_26),
.B2(n_23),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_68),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_104),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_74),
.B(n_70),
.C(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_23),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_132),
.B(n_88),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_115),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_69),
.B1(n_81),
.B2(n_58),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_123),
.B1(n_127),
.B2(n_104),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_120),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_16),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_118),
.C(n_126),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_83),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_105),
.Y(n_136)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_133),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_46),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_134),
.C(n_98),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_31),
.B(n_30),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_1),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_142),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_107),
.B(n_103),
.C(n_87),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_150),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_155),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_93),
.B(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_92),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

AO221x1_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_142),
.B1(n_156),
.B2(n_149),
.C(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_132),
.B1(n_114),
.B2(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_91),
.B1(n_21),
.B2(n_27),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_118),
.B1(n_134),
.B2(n_127),
.C(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_110),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_1),
.B(n_2),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_97),
.C(n_110),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_163),
.C(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_162),
.B1(n_144),
.B2(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_91),
.B1(n_100),
.B2(n_31),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_30),
.C(n_28),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_22),
.B(n_18),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_152),
.B(n_145),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_174),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_135),
.B1(n_145),
.B2(n_4),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_13),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_175),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_22),
.B(n_18),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_176),
.B(n_152),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_28),
.B(n_2),
.C(n_3),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_13),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_168),
.B1(n_163),
.B2(n_174),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_186),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_182),
.B(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_188),
.B(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_162),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_189),
.B1(n_5),
.B2(n_6),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_2),
.B(n_3),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_3),
.C(n_4),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_171),
.C(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_199),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_169),
.B(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_198),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_159),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_197),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_168),
.B1(n_165),
.B2(n_176),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_188),
.B1(n_6),
.B2(n_7),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_181),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_179),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_200),
.A3(n_196),
.B1(n_193),
.B2(n_197),
.C1(n_198),
.C2(n_8),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_5),
.B(n_8),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_184),
.B1(n_183),
.B2(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

AOI31xp33_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_210),
.A3(n_209),
.B(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_5),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_204),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_212),
.B1(n_213),
.B2(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_9),
.B1(n_207),
.B2(n_217),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_216),
.B(n_207),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_222),
.C(n_9),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_224),
.Y(n_229)
);


endmodule