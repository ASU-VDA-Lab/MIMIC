module fake_jpeg_22231_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_22),
.Y(n_67)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_34),
.C(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_35),
.B1(n_24),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_85),
.B1(n_9),
.B2(n_16),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_61),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_37),
.B1(n_35),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_36),
.B1(n_34),
.B2(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_37),
.B1(n_20),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_71),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_37),
.B1(n_29),
.B2(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_36),
.B1(n_23),
.B2(n_29),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_36),
.B1(n_28),
.B2(n_27),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_36),
.B1(n_28),
.B2(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_33),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_25),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_36),
.B1(n_18),
.B2(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_89),
.A2(n_97),
.B1(n_115),
.B2(n_117),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_39),
.B1(n_10),
.B2(n_3),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_104),
.B1(n_108),
.B2(n_54),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_39),
.B(n_2),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_6),
.C(n_7),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_81),
.B(n_80),
.Y(n_132)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_106),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_8),
.B1(n_15),
.B2(n_3),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_17),
.B1(n_9),
.B2(n_4),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_82),
.Y(n_129)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_67),
.B(n_71),
.C(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_145),
.B1(n_106),
.B2(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_134),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_50),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_139),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_118),
.B(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_51),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_52),
.B(n_76),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_150),
.B(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_57),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_53),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_112),
.C(n_95),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_62),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_115),
.B1(n_99),
.B2(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_148),
.B1(n_152),
.B2(n_132),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_53),
.B1(n_52),
.B2(n_65),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_86),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_100),
.B(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_118),
.B1(n_110),
.B2(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_119),
.B(n_115),
.C(n_105),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_159),
.B(n_124),
.Y(n_187)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_157),
.B(n_123),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_170),
.B(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_113),
.B(n_116),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_109),
.B1(n_94),
.B2(n_79),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_94),
.B1(n_88),
.B2(n_112),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_140),
.C(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_112),
.B1(n_95),
.B2(n_13),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_121),
.B1(n_125),
.B2(n_126),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_95),
.B1(n_12),
.B2(n_14),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_11),
.B(n_14),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_184),
.B(n_197),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_188),
.C(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_194),
.B(n_204),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_129),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_170),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_138),
.C(n_142),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_202),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_128),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_203),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_140),
.B(n_150),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_140),
.C(n_143),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_127),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_123),
.B(n_136),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_206),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_137),
.B(n_141),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_187),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_216),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_176),
.B1(n_174),
.B2(n_179),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_224),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_154),
.B1(n_182),
.B2(n_165),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_163),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_185),
.C(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_169),
.Y(n_241)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_193),
.A3(n_198),
.B1(n_207),
.B2(n_205),
.C(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

AOI321xp33_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_194),
.A3(n_190),
.B1(n_199),
.B2(n_193),
.C(n_181),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_219),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_190),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_243),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_184),
.B(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_236),
.B1(n_216),
.B2(n_155),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_155),
.B(n_161),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_200),
.C(n_203),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_242),
.C(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_200),
.C(n_161),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_178),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_221),
.B1(n_208),
.B2(n_226),
.C(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_256),
.C(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_255),
.Y(n_264)
);

OAI322xp33_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_217),
.A3(n_214),
.B1(n_220),
.B2(n_209),
.C1(n_224),
.C2(n_222),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_236),
.C(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_209),
.C(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_253),
.C(n_242),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_225),
.C(n_210),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_160),
.B(n_178),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_178),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_178),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_177),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_156),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_237),
.C(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_244),
.C(n_257),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_253),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_264),
.B(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_254),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_244),
.C(n_254),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_255),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_229),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_265),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_278),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_274),
.C(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_169),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.C(n_166),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_145),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_282),
.B(n_229),
.CI(n_166),
.CON(n_284),
.SN(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_133),
.C(n_135),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_284),
.C(n_121),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_135),
.Y(n_289)
);


endmodule