module fake_jpeg_22803_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_20),
.C(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_52),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_49),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_26),
.B1(n_14),
.B2(n_23),
.Y(n_45)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_2),
.B(n_3),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_26),
.B(n_15),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_21),
.B(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_27),
.B1(n_15),
.B2(n_28),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_22),
.B1(n_15),
.B2(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_20),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_63),
.B1(n_45),
.B2(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_28),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_67),
.B(n_68),
.Y(n_71)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_43),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_21),
.C(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_9),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_9),
.B(n_4),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_48),
.C(n_44),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_59),
.C(n_69),
.Y(n_87)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_76),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_77),
.B(n_60),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_47),
.B1(n_41),
.B2(n_45),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_82),
.B1(n_61),
.B2(n_40),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_45),
.B1(n_51),
.B2(n_40),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_68),
.C(n_59),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_87),
.C(n_91),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_89),
.B(n_93),
.Y(n_103)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_71),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_39),
.C(n_58),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_63),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_97),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_55),
.B(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_40),
.B1(n_51),
.B2(n_80),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_77),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_104),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_73),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_106),
.C(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_90),
.B1(n_84),
.B2(n_75),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_111),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.C(n_98),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_83),
.B(n_75),
.C(n_95),
.D(n_3),
.Y(n_115)
);

OAI21x1_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_83),
.B(n_3),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_5),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_124),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_117),
.C(n_112),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_129),
.C(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_120),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_5),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_125),
.C(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.C(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_5),
.Y(n_138)
);


endmodule