module real_jpeg_30963_n_19 (n_17, n_8, n_0, n_157, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_6, n_159, n_153, n_151, n_11, n_14, n_160, n_7, n_18, n_3, n_5, n_4, n_150, n_1, n_158, n_16, n_15, n_13, n_155, n_19);

input n_17;
input n_8;
input n_0;
input n_157;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_6;
input n_159;
input n_153;
input n_151;
input n_11;
input n_14;
input n_160;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_0),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_139),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_11),
.B1(n_86),
.B2(n_90),
.C(n_94),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_5),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_9),
.B(n_70),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_11),
.B(n_86),
.C(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_52),
.A3(n_54),
.B1(n_62),
.B2(n_128),
.C1(n_130),
.C2(n_160),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_118),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_14),
.B(n_64),
.Y(n_126)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_34),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_145),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_136),
.B(n_142),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_31),
.B(n_134),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_24),
.B(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_29),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_40),
.B(n_133),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI31xp67_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_75),
.A3(n_116),
.B(n_123),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_61),
.C(n_69),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_43),
.A2(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_45),
.B(n_69),
.C(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_151),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

OA21x2_ASAP7_75t_SL g124 ( 
.A1(n_61),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_106),
.C(n_107),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_98),
.B(n_105),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B1(n_96),
.B2(n_97),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_156),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_150),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_152),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_153),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_154),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_155),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_157),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_158),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_159),
.Y(n_119)
);


endmodule