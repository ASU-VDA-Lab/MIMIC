module fake_jpeg_25986_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_23),
.B1(n_17),
.B2(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_17),
.B(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_10),
.B1(n_15),
.B2(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_27),
.B1(n_20),
.B2(n_16),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_21),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_38),
.B1(n_27),
.B2(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_23),
.B1(n_22),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_30),
.B2(n_38),
.Y(n_49)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_34),
.Y(n_52)
);

AOI32xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_31),
.A3(n_46),
.B1(n_42),
.B2(n_39),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_40),
.B(n_9),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_36),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_45),
.CI(n_46),
.CON(n_55),
.SN(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_50),
.C(n_42),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_60),
.B(n_51),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_44),
.C(n_55),
.Y(n_67)
);

AO221x1_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.C(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_59),
.B1(n_54),
.B2(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_63),
.A3(n_14),
.B1(n_7),
.B2(n_5),
.C1(n_6),
.C2(n_13),
.Y(n_68)
);

NAND4xp25_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_0),
.C(n_2),
.D(n_3),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_0),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_70),
.B2(n_3),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_19),
.C(n_2),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_19),
.Y(n_75)
);


endmodule