module fake_jpeg_20785_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_26),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_27),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_57),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_16),
.B1(n_21),
.B2(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_52),
.B1(n_48),
.B2(n_17),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_21),
.B1(n_16),
.B2(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_26),
.Y(n_54)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_59),
.B(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_19),
.B1(n_20),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_78),
.B1(n_45),
.B2(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_25),
.C(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_29),
.B1(n_31),
.B2(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_102),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_84),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_46),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_100),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_37),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_101),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_40),
.B1(n_36),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_40),
.B1(n_27),
.B2(n_22),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_36),
.B1(n_42),
.B2(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_24),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_103),
.B(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_43),
.B1(n_32),
.B2(n_18),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_53),
.B1(n_72),
.B2(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_54),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_28),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_82),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_128),
.B1(n_131),
.B2(n_117),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_115),
.B1(n_85),
.B2(n_117),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_50),
.B(n_37),
.C(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_109),
.C(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_133),
.C(n_142),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_77),
.B1(n_60),
.B2(n_50),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_71),
.B(n_99),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_41),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_41),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_146),
.B(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_41),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_28),
.B(n_7),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_157),
.B(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_97),
.B1(n_96),
.B2(n_84),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_163),
.B1(n_164),
.B2(n_168),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_144),
.C(n_127),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_141),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_171),
.C(n_174),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_116),
.B(n_42),
.Y(n_159)
);

OR2x4_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_81),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_165),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_106),
.B1(n_83),
.B2(n_93),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_106),
.B1(n_64),
.B2(n_94),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_106),
.B1(n_83),
.B2(n_64),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_140),
.B1(n_127),
.B2(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_104),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_60),
.B1(n_68),
.B2(n_65),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_123),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_131),
.B1(n_133),
.B2(n_124),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_173),
.B1(n_125),
.B2(n_119),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_41),
.C(n_39),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_41),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_42),
.B1(n_46),
.B2(n_67),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_41),
.C(n_39),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_126),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_176),
.B(n_181),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_46),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_67),
.B1(n_46),
.B2(n_32),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_179),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_114),
.B(n_1),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_182),
.A2(n_189),
.B1(n_205),
.B2(n_211),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_191),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_148),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_141),
.B(n_81),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_209),
.B(n_172),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_111),
.B(n_82),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_46),
.C(n_125),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_198),
.C(n_201),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_46),
.C(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_32),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_171),
.C(n_168),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_8),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_181),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_8),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_151),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_159),
.B1(n_175),
.B2(n_152),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_236),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_217),
.B(n_194),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_163),
.B1(n_157),
.B2(n_175),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_157),
.B1(n_159),
.B2(n_178),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_172),
.B(n_166),
.C(n_173),
.D(n_177),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_232),
.B(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_0),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_227),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_10),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_0),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_111),
.B1(n_82),
.B2(n_2),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_237),
.B1(n_202),
.B2(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_0),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_233),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_10),
.B(n_15),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_190),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_111),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_257),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_245),
.B1(n_248),
.B2(n_253),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_206),
.B1(n_193),
.B2(n_187),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_195),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_212),
.B1(n_202),
.B2(n_184),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_184),
.C(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_261),
.C(n_215),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_212),
.B1(n_213),
.B2(n_4),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_7),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_226),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_215),
.B(n_6),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_6),
.C(n_13),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_214),
.C(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_274),
.C(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_246),
.A2(n_217),
.B1(n_222),
.B2(n_232),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_225),
.B1(n_237),
.B2(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_234),
.B1(n_11),
.B2(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_248),
.C(n_246),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_249),
.B(n_261),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_220),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_228),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_249),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_252),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_274),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_243),
.B1(n_245),
.B2(n_240),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_297)
);

NAND4xp25_ASAP7_75t_SL g290 ( 
.A(n_262),
.B(n_242),
.C(n_234),
.D(n_253),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_263),
.B1(n_277),
.B2(n_278),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_302),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_296),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_304),
.B1(n_292),
.B2(n_281),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_269),
.C(n_12),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_293),
.C(n_282),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_284),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_312),
.Y(n_317)
);

XOR2x2_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_292),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_298),
.C(n_296),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_311),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_315),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_303),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_309),
.B(n_307),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_319),
.B1(n_314),
.B2(n_313),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_308),
.B(n_312),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_288),
.C(n_284),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.C(n_13),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_14),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_4),
.C(n_1),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_1),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_3),
.B(n_255),
.Y(n_327)
);


endmodule