module fake_jpeg_29395_n_362 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_362);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_362;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_50),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_54),
.B(n_0),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR4xp25_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_6),
.C(n_12),
.D(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_67),
.B(n_47),
.Y(n_129)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_13),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_73),
.Y(n_109)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_12),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_77),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_24),
.B1(n_38),
.B2(n_26),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_102),
.B1(n_107),
.B2(n_113),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_39),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_114),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_74),
.A2(n_38),
.B1(n_26),
.B2(n_24),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_39),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_57),
.A2(n_16),
.B1(n_11),
.B2(n_10),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_121),
.B1(n_122),
.B2(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_118),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_4),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_44),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_1),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_3),
.B1(n_73),
.B2(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_78),
.B1(n_68),
.B2(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_65),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_112),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_43),
.B1(n_42),
.B2(n_36),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_54),
.B(n_56),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_114),
.Y(n_164)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_132),
.CON(n_133),
.SN(n_133)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_133),
.A2(n_165),
.B(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_141),
.Y(n_194)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_149),
.Y(n_205)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_171),
.Y(n_191)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_160),
.Y(n_184)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_124),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_104),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_96),
.A2(n_95),
.B1(n_123),
.B2(n_91),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_106),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_87),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_172),
.Y(n_200)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2x1_ASAP7_75t_SL g170 ( 
.A(n_87),
.B(n_116),
.Y(n_170)
);

OR2x4_ASAP7_75t_L g171 ( 
.A(n_90),
.B(n_104),
.Y(n_171)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_90),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_174),
.Y(n_208)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_100),
.B1(n_119),
.B2(n_143),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_90),
.C(n_86),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_160),
.Y(n_221)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_97),
.B1(n_115),
.B2(n_131),
.Y(n_186)
);

AO22x1_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_197),
.B1(n_176),
.B2(n_191),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_135),
.A2(n_124),
.B(n_131),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_207),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_86),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_153),
.B1(n_152),
.B2(n_142),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_156),
.B1(n_155),
.B2(n_154),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_140),
.B(n_119),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_175),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_135),
.A2(n_170),
.B(n_173),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_135),
.B(n_158),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_142),
.A2(n_171),
.B1(n_133),
.B2(n_138),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_210),
.A2(n_144),
.B1(n_157),
.B2(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_213),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_151),
.B1(n_145),
.B2(n_150),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_237),
.B(n_202),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_229),
.B(n_240),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_225),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_185),
.Y(n_258)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_231),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_172),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_232),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_174),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_137),
.B1(n_136),
.B2(n_139),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_195),
.B1(n_199),
.B2(n_187),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_194),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_236),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_143),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_143),
.B(n_159),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_204),
.B(n_203),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_241),
.A2(n_196),
.B(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_248),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_202),
.B(n_186),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_186),
.B1(n_177),
.B2(n_179),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_251),
.B1(n_264),
.B2(n_218),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_239),
.A2(n_216),
.B1(n_227),
.B2(n_214),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_186),
.B(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_237),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_221),
.A2(n_204),
.B(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_189),
.C(n_180),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_237),
.C(n_238),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_267),
.B(n_287),
.CI(n_187),
.CON(n_305),
.SN(n_305)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_272),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_224),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_271),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_234),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_242),
.C(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_232),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_283),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_244),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_262),
.B1(n_254),
.B2(n_248),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_245),
.A2(n_252),
.B1(n_263),
.B2(n_251),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_285),
.B1(n_264),
.B2(n_215),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_215),
.B1(n_217),
.B2(n_241),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_230),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_247),
.B1(n_225),
.B2(n_223),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_265),
.B1(n_180),
.B2(n_231),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_306),
.Y(n_309)
);

OAI31xp33_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_253),
.A3(n_242),
.B(n_243),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_236),
.B(n_199),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_277),
.C(n_280),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_276),
.B(n_282),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_297),
.A2(n_293),
.B(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_303),
.B1(n_287),
.B2(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_281),
.A2(n_274),
.B1(n_267),
.B2(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_265),
.B1(n_211),
.B2(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_305),
.B(n_268),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_260),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_297),
.B1(n_295),
.B2(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_268),
.C(n_288),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_319),
.C(n_290),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_320),
.B(n_305),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_321),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_183),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_292),
.B(n_266),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_330),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_289),
.B1(n_302),
.B2(n_300),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_315),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_329),
.A2(n_331),
.B(n_308),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_291),
.B(n_306),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_291),
.B1(n_212),
.B2(n_222),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_315),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_316),
.B(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_337),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_342),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_347),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_337),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_333),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_330),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_351),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_344),
.A2(n_346),
.B(n_345),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_349),
.B(n_314),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_352),
.B(n_354),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_327),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_341),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_325),
.C(n_331),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_343),
.B(n_335),
.Y(n_358)
);

AOI321xp33_ASAP7_75t_L g360 ( 
.A1(n_358),
.A2(n_359),
.A3(n_356),
.B1(n_328),
.B2(n_307),
.C(n_319),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_309),
.C(n_212),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_190),
.Y(n_362)
);


endmodule