module fake_jpeg_31743_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_15),
.A2(n_2),
.B(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_26),
.C(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_74),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_22),
.B1(n_32),
.B2(n_18),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_18),
.B1(n_23),
.B2(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_4),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_21),
.B1(n_17),
.B2(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_48),
.C(n_28),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_52),
.C(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_54),
.B1(n_59),
.B2(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_98),
.B1(n_75),
.B2(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_10),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_14),
.B(n_7),
.C(n_9),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_11),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_104),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_73),
.B1(n_64),
.B2(n_71),
.Y(n_103)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_98),
.B1(n_90),
.B2(n_5),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_80),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_71),
.CI(n_6),
.CON(n_106),
.SN(n_106)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_60),
.C(n_71),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_111),
.C(n_113),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_60),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_71),
.C(n_12),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_5),
.B(n_14),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_87),
.C(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_91),
.B1(n_84),
.B2(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_132),
.B1(n_99),
.B2(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_106),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_97),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_103),
.B1(n_102),
.B2(n_107),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_100),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_120),
.C(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_100),
.B(n_103),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_132),
.B1(n_108),
.B2(n_5),
.C(n_117),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_120),
.C(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_104),
.C(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_114),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_132),
.B1(n_127),
.B2(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_144),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_141),
.B1(n_133),
.B2(n_138),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_108),
.B1(n_139),
.B2(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_153),
.B1(n_148),
.B2(n_138),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_134),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.C(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_145),
.C(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_167),
.C(n_154),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_162),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_155),
.B1(n_161),
.B2(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);


endmodule