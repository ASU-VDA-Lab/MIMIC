module fake_jpeg_7756_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_53),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_58),
.Y(n_66)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_1),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_36),
.B1(n_47),
.B2(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_43),
.B1(n_35),
.B2(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_75),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_2),
.B1(n_10),
.B2(n_11),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_15),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_14),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.C(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_80),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_78),
.C(n_89),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_87),
.B(n_82),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_87),
.C(n_84),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_82),
.B(n_79),
.C(n_84),
.D(n_25),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_16),
.B(n_18),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_23),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_26),
.B(n_27),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_29),
.CON(n_104),
.SN(n_104)
);


endmodule