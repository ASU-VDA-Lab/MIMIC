module fake_jpeg_23157_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_41),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_48),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_54),
.Y(n_89)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_30),
.C(n_34),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_72),
.C(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_81),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_83),
.B1(n_23),
.B2(n_25),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_21),
.B1(n_33),
.B2(n_27),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_78),
.B(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_34),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_20),
.B1(n_26),
.B2(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_18),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_33),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_98),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_87),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_90),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_91),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_92),
.B(n_99),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_14),
.B(n_15),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_103),
.B(n_15),
.Y(n_147)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_42),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_105),
.C(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_41),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_26),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_111),
.B1(n_117),
.B2(n_58),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_55),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_73),
.B1(n_45),
.B2(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_59),
.B1(n_33),
.B2(n_45),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_37),
.C(n_52),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_122),
.B1(n_18),
.B2(n_23),
.Y(n_131)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_25),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_25),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_127),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_121),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_0),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_147),
.B(n_104),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_135),
.B1(n_111),
.B2(n_120),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_58),
.B1(n_76),
.B2(n_17),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_23),
.B(n_32),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_142),
.B(n_105),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_76),
.B1(n_32),
.B2(n_40),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_35),
.B(n_2),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_85),
.A2(n_40),
.B1(n_35),
.B2(n_3),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_149),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_154),
.B(n_155),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_112),
.B1(n_94),
.B2(n_92),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_163),
.B1(n_174),
.B2(n_187),
.Y(n_204)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_94),
.C(n_113),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_160),
.C(n_172),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_84),
.C(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_162),
.A2(n_178),
.B(n_7),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_112),
.B1(n_97),
.B2(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_171),
.Y(n_205)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_86),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_118),
.B1(n_116),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_134),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_114),
.B(n_119),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_181),
.B(n_152),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_93),
.B1(n_107),
.B2(n_117),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_122),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_93),
.B1(n_95),
.B2(n_110),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_102),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_185),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_93),
.B1(n_91),
.B2(n_87),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_99),
.B(n_120),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_14),
.C(n_13),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_88),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_130),
.Y(n_197)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_129),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_203),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_139),
.B1(n_151),
.B2(n_147),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_209),
.B1(n_213),
.B2(n_164),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_139),
.B1(n_136),
.B2(n_151),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_151),
.B1(n_140),
.B2(n_134),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_200),
.B1(n_211),
.B2(n_218),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_125),
.B1(n_130),
.B2(n_152),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_222),
.B1(n_155),
.B2(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_214),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_185),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_198),
.A2(n_207),
.B(n_217),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_146),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_156),
.B(n_6),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_221),
.C(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_6),
.B(n_7),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_12),
.C(n_9),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_194),
.B1(n_198),
.B2(n_209),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_246),
.B(n_250),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_154),
.C(n_161),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_240),
.C(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_165),
.B1(n_169),
.B2(n_179),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_237),
.B1(n_244),
.B2(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_176),
.Y(n_238)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_167),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_174),
.C(n_169),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_162),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_241),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_249),
.B1(n_241),
.B2(n_226),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_181),
.B1(n_185),
.B2(n_158),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_181),
.C(n_166),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_10),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_223),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_212),
.B1(n_216),
.B2(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_190),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_215),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_242),
.B1(n_234),
.B2(n_246),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_221),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_267),
.C(n_273),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_195),
.B1(n_207),
.B2(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_227),
.A2(n_201),
.B1(n_197),
.B2(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_10),
.B1(n_11),
.B2(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_10),
.C(n_11),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_256),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_10),
.B(n_11),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_247),
.B(n_239),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_11),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_275),
.B(n_258),
.Y(n_307)
);

XNOR2x2_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_224),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_279),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_229),
.Y(n_279)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_238),
.C(n_235),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.C(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_228),
.C(n_227),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_262),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_223),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_231),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_292),
.B1(n_258),
.B2(n_269),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_257),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_233),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.Y(n_310)
);

AO221x1_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_250),
.B1(n_230),
.B2(n_264),
.C(n_255),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_286),
.C(n_287),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_272),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_263),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_306),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_274),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_309),
.C(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_284),
.B(n_274),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_316),
.B(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_276),
.C(n_280),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_285),
.B1(n_277),
.B2(n_284),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_276),
.C(n_279),
.Y(n_316)
);

OAI221xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_275),
.B1(n_303),
.B2(n_297),
.C(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_301),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_323),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_308),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_298),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_329),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_311),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_336),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_281),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_335),
.B(n_271),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_307),
.B(n_304),
.Y(n_335)
);

NOR5xp2_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_268),
.C(n_315),
.D(n_293),
.E(n_316),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_340),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_334),
.B(n_325),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_312),
.B(n_338),
.Y(n_343)
);

OAI221xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_342),
.B1(n_251),
.B2(n_293),
.C(n_261),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_267),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_273),
.Y(n_347)
);


endmodule