module fake_aes_2091_n_724 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_724);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_724;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_43), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_69), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_22), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_42), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_41), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_37), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_47), .Y(n_87) );
INVx3_ASAP7_75t_L g88 ( .A(n_3), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_79), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_0), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_65), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_55), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_68), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_54), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_56), .Y(n_96) );
BUFx2_ASAP7_75t_L g97 ( .A(n_16), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_51), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_12), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_73), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_50), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_12), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_11), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_2), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_9), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_45), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_25), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_35), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_48), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_31), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_7), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_77), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_59), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_1), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_17), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_97), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_90), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_88), .B(n_4), .Y(n_135) );
OR2x6_ASAP7_75t_L g136 ( .A(n_88), .B(n_4), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_118), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_82), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_87), .B(n_5), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_125), .B(n_5), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_110), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_111), .B(n_80), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_110), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_81), .B(n_34), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_105), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_105), .B(n_6), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_125), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_124), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
CKINVDCx11_ASAP7_75t_R g161 ( .A(n_107), .Y(n_161) );
OAI22x1_ASAP7_75t_R g162 ( .A1(n_112), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_91), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_92), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_96), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_99), .A2(n_130), .B(n_116), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_103), .Y(n_169) );
BUFx12f_ASAP7_75t_L g170 ( .A(n_81), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_112), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_121), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_109), .A2(n_38), .B(n_75), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_114), .Y(n_175) );
INVx4_ASAP7_75t_SL g176 ( .A(n_136), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_149), .B(n_106), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_133), .B(n_113), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_158), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_170), .Y(n_183) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_136), .A2(n_123), .B1(n_113), .B2(n_127), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_133), .B(n_123), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_135), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_132), .Y(n_192) );
XNOR2xp5_ASAP7_75t_L g193 ( .A(n_139), .B(n_101), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
BUFx10_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_137), .B(n_129), .C(n_128), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_133), .B(n_93), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_141), .B(n_128), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_136), .A2(n_83), .B1(n_119), .B2(n_84), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_175), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_141), .B(n_108), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_170), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_150), .B(n_120), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_166), .B(n_120), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_136), .A2(n_83), .B1(n_84), .B2(n_106), .Y(n_217) );
BUFx10_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_150), .B(n_119), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_149), .B(n_85), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_136), .Y(n_224) );
NAND2xp33_ASAP7_75t_L g225 ( .A(n_166), .B(n_85), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_155), .B(n_104), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_155), .B(n_100), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_115), .B1(n_102), .B2(n_14), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_137), .B(n_10), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_166), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_157), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_166), .B(n_36), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_165), .B(n_13), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_165), .B(n_13), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_154), .B(n_14), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_160), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_167), .B(n_40), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_160), .Y(n_241) );
INVx5_ASAP7_75t_L g242 ( .A(n_166), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_179), .B(n_173), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_203), .B(n_142), .Y(n_245) );
NOR2x2_ASAP7_75t_L g246 ( .A(n_193), .B(n_159), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_185), .B(n_173), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_212), .B(n_142), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_220), .B(n_156), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_229), .B(n_156), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_176), .B(n_172), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
AO22x1_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_134), .B1(n_162), .B2(n_161), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_202), .B(n_172), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_176), .B(n_167), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_153), .B1(n_134), .B2(n_164), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_206), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_215), .B(n_164), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_202), .B(n_164), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_231), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_188), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_202), .B(n_168), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_238), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_176), .B(n_169), .Y(n_266) );
NOR2xp33_ASAP7_75t_SL g267 ( .A(n_224), .B(n_163), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_227), .A2(n_223), .B1(n_177), .B2(n_224), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_218), .B(n_147), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_226), .B(n_168), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_183), .B(n_174), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_199), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_182), .A2(n_168), .B(n_174), .Y(n_275) );
BUFx12f_ASAP7_75t_L g276 ( .A(n_218), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_177), .A2(n_169), .B1(n_147), .B2(n_140), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_238), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_192), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_223), .A2(n_184), .B1(n_207), .B2(n_217), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_190), .A2(n_174), .B(n_163), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_194), .Y(n_282) );
AOI22xp33_ASAP7_75t_SL g283 ( .A1(n_187), .A2(n_162), .B1(n_147), .B2(n_144), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_178), .Y(n_284) );
AND2x6_ASAP7_75t_SL g285 ( .A(n_193), .B(n_15), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_176), .B(n_169), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_188), .A2(n_163), .B1(n_147), .B2(n_140), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_188), .A2(n_204), .B1(n_178), .B2(n_186), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_178), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_186), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_186), .Y(n_292) );
NOR2x2_ASAP7_75t_L g293 ( .A(n_211), .B(n_15), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_204), .B(n_140), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_201), .A2(n_140), .B1(n_144), .B2(n_169), .Y(n_295) );
AND2x6_ASAP7_75t_L g296 ( .A(n_204), .B(n_169), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_200), .B(n_144), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_SL g298 ( .A1(n_240), .A2(n_144), .B(n_131), .C(n_151), .Y(n_298) );
INVx8_ASAP7_75t_L g299 ( .A(n_211), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_234), .B(n_169), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_199), .B(n_174), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_199), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_237), .B(n_151), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_209), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_214), .A2(n_174), .B1(n_151), .B2(n_148), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_222), .B(n_148), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_233), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_239), .B(n_148), .Y(n_311) );
AND2x6_ASAP7_75t_SL g312 ( .A(n_241), .B(n_18), .Y(n_312) );
AND2x6_ASAP7_75t_SL g313 ( .A(n_230), .B(n_20), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_260), .B(n_225), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_302), .A2(n_213), .B(n_225), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_265), .A2(n_213), .B(n_235), .C(n_208), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_278), .B(n_235), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_264), .A2(n_232), .B(n_228), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_253), .B(n_208), .C(n_219), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_274), .B(n_242), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
O2A1O1Ixp5_ASAP7_75t_L g322 ( .A1(n_307), .A2(n_232), .B(n_228), .C(n_198), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_270), .A2(n_197), .B(n_221), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_244), .A2(n_242), .B1(n_221), .B2(n_219), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_262), .A2(n_242), .B1(n_205), .B2(n_198), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_274), .B(n_242), .Y(n_326) );
NOR3xp33_ASAP7_75t_SL g327 ( .A(n_269), .B(n_21), .C(n_23), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_280), .A2(n_205), .B1(n_197), .B2(n_242), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_274), .B(n_196), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_290), .B(n_196), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_303), .B(n_196), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_252), .A2(n_131), .B1(n_145), .B2(n_146), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_250), .B(n_131), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_263), .Y(n_334) );
NOR2xp33_ASAP7_75t_R g335 ( .A(n_299), .B(n_24), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_256), .A2(n_181), .B1(n_189), .B2(n_191), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_275), .A2(n_181), .B(n_189), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_251), .B(n_26), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_245), .B(n_146), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_303), .B(n_196), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_248), .A2(n_146), .B(n_145), .C(n_191), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_258), .B(n_28), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_303), .B(n_195), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_243), .B(n_145), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_299), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_247), .B(n_195), .Y(n_347) );
AOI21x1_ASAP7_75t_L g348 ( .A1(n_281), .A2(n_195), .B(n_180), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_263), .Y(n_349) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_304), .B(n_195), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_283), .B(n_195), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_263), .B(n_180), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_249), .B(n_254), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_294), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_305), .A2(n_180), .B(n_30), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_251), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_279), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_267), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_282), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_261), .B(n_29), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_284), .A2(n_180), .B(n_39), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_289), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_267), .B(n_180), .C(n_49), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_291), .A2(n_33), .B(n_52), .C(n_53), .Y(n_364) );
INVxp33_ASAP7_75t_SL g365 ( .A(n_246), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_268), .B(n_57), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_292), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_356), .B(n_255), .Y(n_369) );
OAI21x1_ASAP7_75t_SL g370 ( .A1(n_368), .A2(n_297), .B(n_277), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_353), .A2(n_288), .B1(n_310), .B2(n_287), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_SL g372 ( .A1(n_364), .A2(n_298), .B(n_301), .C(n_286), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_345), .Y(n_373) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_315), .A2(n_308), .A3(n_272), .B(n_300), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_318), .A2(n_271), .B(n_257), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_346), .B(n_295), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_353), .A2(n_259), .B(n_311), .C(n_266), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_319), .A2(n_296), .B1(n_273), .B2(n_313), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_358), .A2(n_273), .B(n_309), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_321), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_358), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_339), .A2(n_313), .B(n_293), .C(n_312), .Y(n_382) );
OAI22x1_ASAP7_75t_L g383 ( .A1(n_365), .A2(n_285), .B1(n_312), .B2(n_296), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_357), .Y(n_384) );
CKINVDCx8_ASAP7_75t_R g385 ( .A(n_349), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_342), .A2(n_296), .B1(n_285), .B2(n_63), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_348), .A2(n_296), .B(n_62), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_317), .A2(n_58), .B(n_64), .C(n_70), .Y(n_388) );
CKINVDCx9p33_ASAP7_75t_R g389 ( .A(n_335), .Y(n_389) );
AO32x2_ASAP7_75t_L g390 ( .A1(n_332), .A2(n_74), .A3(n_78), .B1(n_322), .B2(n_325), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_356), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
OAI21xp33_ASAP7_75t_SL g393 ( .A1(n_328), .A2(n_367), .B(n_330), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_354), .B(n_317), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_351), .B(n_338), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_338), .B(n_319), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g398 ( .A1(n_366), .A2(n_347), .B(n_343), .C(n_340), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_334), .Y(n_399) );
BUFx10_ASAP7_75t_L g400 ( .A(n_330), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_334), .B(n_350), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_360), .A2(n_333), .B1(n_314), .B2(n_344), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_397), .A2(n_327), .B1(n_341), .B2(n_336), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_395), .A2(n_327), .B1(n_363), .B2(n_355), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_387), .A2(n_322), .B(n_337), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_402), .A2(n_316), .B(n_323), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_398), .A2(n_329), .B(n_331), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_384), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_395), .A2(n_324), .B1(n_320), .B2(n_326), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_375), .A2(n_361), .B(n_324), .Y(n_411) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_399), .Y(n_412) );
AOI21x1_ASAP7_75t_L g413 ( .A1(n_379), .A2(n_352), .B(n_370), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
OR2x6_ASAP7_75t_L g415 ( .A(n_382), .B(n_383), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_371), .A2(n_393), .B1(n_386), .B2(n_394), .C(n_373), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_372), .A2(n_393), .B(n_377), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_378), .B(n_376), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_373), .B(n_385), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_391), .B(n_380), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_378), .A2(n_381), .B(n_388), .Y(n_422) );
AO31x2_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_374), .A3(n_400), .B(n_401), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_401), .B(n_369), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_390), .A2(n_374), .B(n_400), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_369), .A2(n_397), .B1(n_395), .B2(n_378), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_358), .B(n_402), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_393), .A2(n_382), .B(n_397), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_380), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_382), .A2(n_393), .B(n_353), .C(n_280), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_424), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_407), .B(n_414), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_428), .A2(n_417), .B(n_422), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_419), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_409), .B(n_431), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_423), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_418), .B(n_429), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_418), .B(n_429), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_423), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_426), .B(n_415), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_426), .B(n_415), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_430), .B(n_412), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_415), .A2(n_416), .B1(n_427), .B2(n_420), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_423), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_425), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_406), .A2(n_408), .B(n_403), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_403), .B1(n_410), .B2(n_421), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_410), .B(n_404), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_411), .Y(n_453) );
OR2x6_ASAP7_75t_L g454 ( .A(n_411), .B(n_426), .Y(n_454) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_428), .A2(n_417), .B(n_422), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_428), .A2(n_417), .B(n_405), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
OR2x6_ASAP7_75t_L g459 ( .A(n_426), .B(n_415), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
OR2x6_ASAP7_75t_L g462 ( .A(n_426), .B(n_415), .Y(n_462) );
OR2x6_ASAP7_75t_L g463 ( .A(n_426), .B(n_415), .Y(n_463) );
INVx4_ASAP7_75t_SL g464 ( .A(n_415), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_431), .A2(n_393), .B(n_382), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_424), .B(n_395), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_446), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_446), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_438), .B(n_439), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_446), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_438), .B(n_439), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_452), .B(n_433), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_436), .B(n_452), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_465), .A2(n_462), .B1(n_443), .B2(n_459), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_458), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_433), .B(n_460), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_451), .B(n_447), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_460), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_441), .B(n_463), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_461), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_461), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_459), .B(n_463), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_459), .B(n_463), .Y(n_487) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_450), .A2(n_442), .B(n_453), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_459), .B(n_463), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_456), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_463), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_443), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_445), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_443), .B(n_462), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_462), .B(n_432), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_462), .B(n_464), .Y(n_500) );
NOR2xp67_ASAP7_75t_L g501 ( .A(n_437), .B(n_448), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_467), .B(n_432), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_454), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_440), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_432), .B(n_454), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_454), .B(n_448), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_440), .B(n_434), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_449), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_442), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_446), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_434), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_454), .B(n_434), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_455), .B(n_466), .Y(n_513) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_455), .A2(n_457), .B(n_466), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_464), .B(n_455), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_457), .B(n_464), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_472), .B(n_457), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_495), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_473), .B(n_464), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_472), .B(n_457), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_500), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_470), .B(n_466), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_473), .B(n_466), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_494), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_480), .B(n_444), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_494), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_475), .B(n_480), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_477), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_475), .B(n_481), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_506), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_500), .B(n_515), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_477), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_502), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_506), .B(n_511), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_479), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_498), .B(n_490), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_502), .B(n_481), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVx5_ASAP7_75t_L g541 ( .A(n_468), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_479), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_495), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_511), .B(n_505), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_513), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_500), .B(n_515), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_482), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_513), .B(n_482), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_508), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_484), .B(n_485), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_498), .B(n_484), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g552 ( .A(n_500), .B(n_515), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_490), .B(n_483), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_496), .B(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_508), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_499), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_479), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_490), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_474), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_504), .B(n_474), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_497), .B(n_514), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_476), .B(n_507), .C(n_504), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_501), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_497), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_514), .B(n_486), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_514), .B(n_486), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_507), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_545), .B(n_514), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_545), .B(n_503), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_529), .B(n_476), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_517), .B(n_503), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_525), .A2(n_496), .B1(n_493), .B2(n_492), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_530), .B(n_493), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_527), .B(n_496), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_530), .B(n_492), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_552), .B(n_491), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_539), .B(n_491), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_517), .B(n_489), .Y(n_582) );
NAND2x1_ASAP7_75t_L g583 ( .A(n_552), .B(n_561), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_520), .B(n_489), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_520), .B(n_487), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_548), .B(n_487), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_521), .B(n_512), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_536), .Y(n_589) );
NAND2x1_ASAP7_75t_L g590 ( .A(n_561), .B(n_515), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_544), .B(n_512), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_509), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_518), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_544), .B(n_516), .Y(n_595) );
INVxp33_ASAP7_75t_L g596 ( .A(n_563), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_548), .B(n_516), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_531), .B(n_516), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_567), .B(n_568), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_528), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_567), .B(n_488), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_536), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_532), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
CKINVDCx16_ASAP7_75t_R g605 ( .A(n_561), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_564), .B(n_469), .C(n_471), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_509), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_568), .B(n_488), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_534), .B(n_562), .Y(n_610) );
NOR2x1p5_ASAP7_75t_L g611 ( .A(n_561), .B(n_469), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_534), .B(n_488), .Y(n_612) );
INVx3_ASAP7_75t_SL g613 ( .A(n_542), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_535), .B(n_547), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_488), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_562), .B(n_469), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_535), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_469), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_540), .B(n_471), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_543), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_537), .B(n_471), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_610), .B(n_546), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_610), .B(n_546), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_570), .B(n_546), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_613), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_614), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_573), .B(n_551), .Y(n_629) );
NOR2xp67_ASAP7_75t_L g630 ( .A(n_599), .B(n_546), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_596), .B(n_554), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_570), .B(n_526), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_572), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_581), .B(n_526), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_584), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_597), .B(n_566), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_600), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_589), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_583), .B(n_542), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_603), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_592), .B(n_537), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_608), .B(n_569), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_602), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_599), .B(n_524), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_569), .B(n_524), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_596), .B(n_550), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_587), .B(n_560), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_612), .B(n_531), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_613), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_612), .B(n_531), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_582), .B(n_531), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_591), .B(n_550), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_591), .B(n_547), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_582), .B(n_565), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_593), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_585), .B(n_565), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_622), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_607), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_577), .B(n_519), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_575), .B(n_564), .C(n_523), .D(n_557), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_645), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_646), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_635), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_631), .A2(n_575), .B1(n_601), .B2(n_609), .Y(n_665) );
OAI32xp33_ASAP7_75t_L g666 ( .A1(n_627), .A2(n_605), .A3(n_588), .B1(n_578), .B2(n_576), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_637), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_631), .A2(n_601), .B1(n_609), .B2(n_574), .C1(n_571), .C2(n_616), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_627), .B(n_586), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_661), .A2(n_585), .B1(n_586), .B2(n_571), .C(n_574), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_629), .A2(n_579), .B1(n_616), .B2(n_558), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_640), .Y(n_672) );
OA21x2_ASAP7_75t_SL g673 ( .A1(n_652), .A2(n_598), .B(n_579), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_659), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_628), .B(n_615), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_638), .B(n_606), .C(n_619), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_626), .B(n_595), .Y(n_677) );
AOI22xp5_ASAP7_75t_SL g678 ( .A1(n_649), .A2(n_598), .B1(n_595), .B2(n_579), .Y(n_678) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_639), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_660), .A2(n_617), .B1(n_598), .B2(n_540), .C(n_558), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_644), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_654), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_642), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_647), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_649), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_675), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_668), .B(n_632), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_665), .A2(n_633), .B1(n_630), .B2(n_643), .C(n_639), .Y(n_688) );
OAI21xp5_ASAP7_75t_SL g689 ( .A1(n_679), .A2(n_625), .B(n_623), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_679), .A2(n_625), .B(n_623), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_685), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_670), .B(n_658), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_678), .A2(n_579), .B1(n_590), .B2(n_651), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_664), .Y(n_694) );
NAND3xp33_ASAP7_75t_SL g695 ( .A(n_680), .B(n_673), .C(n_665), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_669), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_666), .A2(n_648), .B(n_650), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_667), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_676), .B(n_660), .C(n_634), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_695), .A2(n_671), .B(n_663), .C(n_662), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_688), .A2(n_671), .B1(n_681), .B2(n_682), .C(n_683), .Y(n_701) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_695), .A2(n_684), .A3(n_626), .B1(n_648), .B2(n_650), .C1(n_657), .C2(n_655), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_687), .A2(n_674), .B1(n_672), .B2(n_657), .C(n_655), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_696), .A2(n_651), .B1(n_677), .B2(n_636), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_689), .A2(n_641), .B1(n_611), .B2(n_622), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_692), .A2(n_656), .B1(n_653), .B2(n_624), .C(n_618), .Y(n_706) );
NOR2x1p5_ASAP7_75t_L g707 ( .A(n_699), .B(n_618), .Y(n_707) );
NOR2xp33_ASAP7_75t_SL g708 ( .A(n_705), .B(n_691), .Y(n_708) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_700), .B(n_690), .C(n_693), .Y(n_709) );
NAND3x2_ASAP7_75t_L g710 ( .A(n_702), .B(n_686), .C(n_701), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_703), .A2(n_698), .B1(n_694), .B2(n_697), .C(n_656), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_706), .B(n_653), .C(n_624), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_710), .B(n_707), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_709), .B(n_704), .C(n_555), .D(n_549), .Y(n_714) );
NAND3xp33_ASAP7_75t_SL g715 ( .A(n_708), .B(n_560), .C(n_559), .Y(n_715) );
OR5x1_ASAP7_75t_L g716 ( .A(n_714), .B(n_711), .C(n_712), .D(n_541), .E(n_510), .Y(n_716) );
AND3x2_ASAP7_75t_L g717 ( .A(n_713), .B(n_621), .C(n_620), .Y(n_717) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_716), .A2(n_715), .B(n_555), .Y(n_718) );
OA22x2_ASAP7_75t_L g719 ( .A1(n_717), .A2(n_621), .B1(n_593), .B2(n_620), .Y(n_719) );
OAI21x1_ASAP7_75t_SL g720 ( .A1(n_718), .A2(n_594), .B(n_604), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_721), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_719), .B1(n_541), .B2(n_549), .Y(n_723) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_541), .B1(n_594), .B2(n_604), .C1(n_556), .C2(n_471), .Y(n_724) );
endmodule