module fake_jpeg_24052_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_2),
.Y(n_63)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_41),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_15),
.Y(n_52)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_29),
.Y(n_58)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_1),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_22),
.B(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_50),
.B1(n_27),
.B2(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_30),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_25),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_15),
.C(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_45),
.B1(n_51),
.B2(n_10),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_17),
.B(n_14),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_90),
.B(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_37),
.B1(n_38),
.B2(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_85),
.B1(n_88),
.B2(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_82),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_48),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_65),
.C(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_96),
.C(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_99),
.B1(n_76),
.B2(n_92),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_64),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_62),
.B(n_26),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_3),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_45),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_109),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_80),
.B1(n_82),
.B2(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_7),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_73),
.Y(n_116)
);

BUFx12f_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_119),
.B(n_105),
.C(n_107),
.Y(n_129)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_77),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_104),
.C(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_97),
.B(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_117),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_97),
.C(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_112),
.C(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_140),
.C(n_141),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_118),
.B(n_113),
.C(n_122),
.D(n_114),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_112),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_146),
.B(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_150),
.C(n_140),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_149),
.B(n_151),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_131),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_83),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_108),
.B1(n_103),
.B2(n_51),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.C(n_72),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_141),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_143),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_108),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_160),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_155),
.B1(n_156),
.B2(n_72),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_8),
.C(n_11),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);


endmodule