module real_aes_3625_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_905;
wire n_357;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_892;
wire n_372;
wire n_202;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g239 ( .A(n_0), .B(n_171), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_1), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_2), .A2(n_16), .B1(n_903), .B2(n_904), .Y(n_902) );
INVx1_ASAP7_75t_L g904 ( .A(n_2), .Y(n_904) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_3), .A2(n_135), .B(n_176), .C(n_178), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g244 ( .A1(n_4), .A2(n_85), .B1(n_134), .B2(n_140), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_5), .A2(n_33), .B1(n_549), .B2(n_550), .Y(n_548) );
INVxp67_ASAP7_75t_L g510 ( .A(n_6), .Y(n_510) );
INVx1_ASAP7_75t_L g893 ( .A(n_6), .Y(n_893) );
INVx1_ASAP7_75t_L g896 ( .A(n_6), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_7), .A2(n_92), .B1(n_585), .B2(n_586), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_8), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_9), .A2(n_71), .B1(n_138), .B2(n_140), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_10), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_11), .A2(n_34), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_12), .A2(n_105), .B1(n_917), .B2(n_924), .Y(n_104) );
INVx2_ASAP7_75t_L g609 ( .A(n_13), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_14), .A2(n_63), .B1(n_132), .B2(n_134), .Y(n_131) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_15), .A2(n_70), .B(n_149), .Y(n_148) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_15), .A2(n_70), .B(n_149), .Y(n_151) );
INVx1_ASAP7_75t_L g903 ( .A(n_16), .Y(n_903) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_17), .B(n_618), .Y(n_617) );
XOR2x2_ASAP7_75t_L g503 ( .A(n_18), .B(n_52), .Y(n_503) );
INVx1_ASAP7_75t_SL g607 ( .A(n_19), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_20), .B(n_146), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_21), .Y(n_268) );
BUFx3_ASAP7_75t_L g110 ( .A(n_22), .Y(n_110) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_23), .A2(n_183), .B(n_184), .C(n_186), .Y(n_182) );
OAI22xp33_ASAP7_75t_SL g242 ( .A1(n_24), .A2(n_49), .B1(n_134), .B2(n_161), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_25), .A2(n_31), .B1(n_161), .B2(n_166), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g624 ( .A1(n_26), .A2(n_538), .B(n_625), .C(n_628), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_27), .B(n_555), .Y(n_615) );
O2A1O1Ixp5_ASAP7_75t_L g198 ( .A1(n_28), .A2(n_135), .B(n_199), .C(n_201), .Y(n_198) );
INVx1_ASAP7_75t_L g515 ( .A(n_29), .Y(n_515) );
INVx1_ASAP7_75t_SL g633 ( .A(n_30), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_32), .Y(n_115) );
AND2x2_ASAP7_75t_L g922 ( .A(n_35), .B(n_923), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_36), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_37), .B(n_216), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_38), .A2(n_42), .B1(n_554), .B2(n_556), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_39), .A2(n_69), .B1(n_556), .B2(n_573), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_40), .B(n_551), .Y(n_614) );
INVx2_ASAP7_75t_L g566 ( .A(n_41), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_43), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_44), .B(n_297), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_45), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_46), .A2(n_186), .B(n_605), .C(n_606), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_47), .A2(n_898), .B1(n_899), .B2(n_905), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_47), .Y(n_905) );
INVx1_ASAP7_75t_L g682 ( .A(n_48), .Y(n_682) );
INVx2_ASAP7_75t_L g634 ( .A(n_50), .Y(n_634) );
INVx1_ASAP7_75t_L g149 ( .A(n_51), .Y(n_149) );
AND2x4_ASAP7_75t_L g144 ( .A(n_53), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g189 ( .A(n_53), .B(n_145), .Y(n_189) );
INVx2_ASAP7_75t_L g574 ( .A(n_54), .Y(n_574) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_55), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_56), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_57), .Y(n_208) );
INVx2_ASAP7_75t_L g167 ( .A(n_58), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_59), .A2(n_135), .B(n_270), .C(n_271), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_60), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_61), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_61), .Y(n_900) );
INVx1_ASAP7_75t_SL g629 ( .A(n_62), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_64), .A2(n_80), .B1(n_177), .B2(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_65), .B(n_146), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_66), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_67), .Y(n_254) );
NAND2xp33_ASAP7_75t_R g150 ( .A(n_68), .B(n_151), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_68), .A2(n_103), .B1(n_216), .B2(n_353), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_72), .A2(n_186), .B(n_549), .C(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_73), .B(n_517), .Y(n_516) );
OR2x6_ASAP7_75t_L g512 ( .A(n_74), .B(n_513), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_75), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g668 ( .A(n_76), .Y(n_668) );
INVx1_ASAP7_75t_L g678 ( .A(n_77), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_78), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_79), .B(n_534), .Y(n_619) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_81), .B(n_199), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_82), .A2(n_135), .B(n_570), .C(n_572), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_82), .A2(n_135), .B(n_570), .C(n_572), .Y(n_658) );
INVx1_ASAP7_75t_L g514 ( .A(n_83), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_84), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_86), .A2(n_96), .B1(n_540), .B2(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g923 ( .A(n_87), .Y(n_923) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
BUFx5_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx1_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVx2_ASAP7_75t_L g191 ( .A(n_89), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_90), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g274 ( .A(n_91), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_93), .Y(n_185) );
INVx2_ASAP7_75t_SL g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g206 ( .A(n_95), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_97), .B(n_151), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_98), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_113) );
INVx1_ASAP7_75t_SL g118 ( .A(n_98), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_98), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_99), .B(n_578), .Y(n_636) );
INVx2_ASAP7_75t_L g211 ( .A(n_100), .Y(n_211) );
AND2x2_ASAP7_75t_L g544 ( .A(n_101), .B(n_158), .Y(n_544) );
OAI21xp33_ASAP7_75t_SL g266 ( .A1(n_102), .A2(n_134), .B(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_103), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_103), .B(n_216), .Y(n_215) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_518), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_110), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_504), .C(n_516), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_118), .B(n_354), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g504 ( .A1(n_119), .A2(n_505), .B(n_506), .Y(n_504) );
XNOR2x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_503), .Y(n_119) );
OAI22x1_ASAP7_75t_L g520 ( .A1(n_120), .A2(n_521), .B1(n_892), .B2(n_894), .Y(n_520) );
AO22x2_ASAP7_75t_L g906 ( .A1(n_120), .A2(n_521), .B1(n_907), .B2(n_908), .Y(n_906) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_400), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_311), .C(n_359), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_256), .Y(n_122) );
OAI21xp33_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_192), .B(n_223), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_124), .A2(n_471), .B(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_152), .Y(n_125) );
OR2x2_ASAP7_75t_L g398 ( .A(n_126), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_126), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g279 ( .A(n_128), .Y(n_279) );
INVx2_ASAP7_75t_L g310 ( .A(n_128), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_128), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g450 ( .A(n_128), .B(n_154), .Y(n_450) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_150), .Y(n_128) );
AND2x2_ASAP7_75t_L g351 ( .A(n_129), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_142), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B1(n_137), .B2(n_141), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_132), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_164) );
INVx1_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_132), .A2(n_134), .B1(n_253), .B2(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g535 ( .A(n_132), .Y(n_535) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_132), .Y(n_605) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g140 ( .A(n_133), .Y(n_140) );
INVx6_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
INVx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_134), .A2(n_161), .B1(n_162), .B2(n_163), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_134), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_134), .B(n_208), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_134), .A2(n_161), .B1(n_250), .B2(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_134), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g534 ( .A(n_134), .Y(n_534) );
INVx2_ASAP7_75t_L g542 ( .A(n_134), .Y(n_542) );
INVx2_ASAP7_75t_L g555 ( .A(n_134), .Y(n_555) );
INVx1_ASAP7_75t_L g571 ( .A(n_134), .Y(n_571) );
INVx2_ASAP7_75t_L g585 ( .A(n_134), .Y(n_585) );
NAND2xp33_ASAP7_75t_L g599 ( .A(n_134), .B(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g159 ( .A1(n_135), .A2(n_141), .B1(n_160), .B2(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g222 ( .A(n_135), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g248 ( .A1(n_135), .A2(n_144), .B1(n_186), .B2(n_249), .C(n_252), .Y(n_248) );
INVx2_ASAP7_75t_SL g590 ( .A(n_135), .Y(n_590) );
INVx1_ASAP7_75t_L g602 ( .A(n_135), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_135), .B(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_135), .B(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
INVx3_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_136), .B(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
INVx1_ASAP7_75t_L g234 ( .A(n_136), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_136), .B(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g588 ( .A(n_136), .Y(n_588) );
INVx2_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx2_ASAP7_75t_L g573 ( .A(n_140), .Y(n_573) );
INVx1_ASAP7_75t_L g673 ( .A(n_140), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_141), .A2(n_204), .B1(n_205), .B2(n_207), .Y(n_203) );
INVx2_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
O2A1O1Ixp5_ASAP7_75t_SL g667 ( .A1(n_141), .A2(n_668), .B(n_669), .C(n_672), .Y(n_667) );
NOR2xp67_ASAP7_75t_L g142 ( .A(n_143), .B(n_146), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_143), .B(n_297), .Y(n_635) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_144), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_144), .B(n_172), .Y(n_245) );
AND2x2_ASAP7_75t_L g543 ( .A(n_144), .B(n_296), .Y(n_543) );
INVx3_ASAP7_75t_L g560 ( .A(n_144), .Y(n_560) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_147), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_147), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
BUFx3_ASAP7_75t_L g297 ( .A(n_148), .Y(n_297) );
BUFx3_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g264 ( .A(n_151), .Y(n_264) );
INVx2_ASAP7_75t_L g354 ( .A(n_151), .Y(n_354) );
INVx1_ASAP7_75t_L g567 ( .A(n_151), .Y(n_567) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_153), .B(n_283), .Y(n_403) );
AND2x2_ASAP7_75t_L g490 ( .A(n_153), .B(n_434), .Y(n_490) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_173), .Y(n_153) );
INVx1_ASAP7_75t_L g307 ( .A(n_154), .Y(n_307) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_159), .B(n_168), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_156), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_156), .B(n_296), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_157), .B(n_189), .Y(n_228) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
INVx2_ASAP7_75t_L g179 ( .A(n_161), .Y(n_179) );
INVx2_ASAP7_75t_SL g233 ( .A(n_161), .Y(n_233) );
INVx1_ASAP7_75t_L g618 ( .A(n_161), .Y(n_618) );
INVx2_ASAP7_75t_L g627 ( .A(n_161), .Y(n_627) );
INVx1_ASAP7_75t_L g671 ( .A(n_161), .Y(n_671) );
INVx1_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_166), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_166), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g541 ( .A(n_166), .Y(n_541) );
INVx2_ASAP7_75t_L g556 ( .A(n_166), .Y(n_556) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx2_ASAP7_75t_L g247 ( .A(n_170), .Y(n_247) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g187 ( .A(n_171), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g190 ( .A(n_172), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g216 ( .A(n_172), .Y(n_216) );
OR2x2_ASAP7_75t_L g213 ( .A(n_173), .B(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_173), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_173), .B(n_196), .Y(n_288) );
INVx2_ASAP7_75t_L g309 ( .A(n_173), .Y(n_309) );
INVx1_ASAP7_75t_L g348 ( .A(n_173), .Y(n_348) );
INVx1_ASAP7_75t_L g389 ( .A(n_173), .Y(n_389) );
AND2x2_ASAP7_75t_L g424 ( .A(n_173), .B(n_214), .Y(n_424) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_173), .Y(n_479) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_181), .A3(n_187), .B(n_190), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g549 ( .A(n_177), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_179), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_183), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_186), .A2(n_244), .B(n_245), .Y(n_243) );
INVx3_ASAP7_75t_L g536 ( .A(n_186), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g197 ( .A(n_188), .B(n_198), .C(n_203), .Y(n_197) );
AOI221xp5_ASAP7_75t_L g218 ( .A1(n_188), .A2(n_219), .B1(n_220), .B2(n_221), .C(n_222), .Y(n_218) );
NOR4xp25_ASAP7_75t_L g568 ( .A(n_188), .B(n_569), .C(n_575), .D(n_578), .Y(n_568) );
NOR2x1_ASAP7_75t_SL g596 ( .A(n_188), .B(n_247), .Y(n_596) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g263 ( .A(n_189), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_213), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g278 ( .A(n_196), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g317 ( .A(n_196), .B(n_309), .Y(n_317) );
INVx2_ASAP7_75t_L g332 ( .A(n_196), .Y(n_332) );
INVx2_ASAP7_75t_L g358 ( .A(n_196), .Y(n_358) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_209), .B(n_210), .Y(n_196) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g204 ( .A(n_200), .Y(n_204) );
INVx1_ASAP7_75t_L g270 ( .A(n_200), .Y(n_270) );
INVx2_ASAP7_75t_L g551 ( .A(n_200), .Y(n_551) );
INVx2_ASAP7_75t_L g586 ( .A(n_200), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_209), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g684 ( .A(n_209), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_213), .Y(n_314) );
OR2x2_ASAP7_75t_L g329 ( .A(n_213), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g406 ( .A(n_213), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_214), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_214), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_214), .B(n_414), .Y(n_440) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g558 ( .A(n_216), .Y(n_558) );
AND2x2_ASAP7_75t_L g350 ( .A(n_217), .B(n_351), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_219), .A2(n_266), .B(n_269), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_219), .A2(n_614), .B(n_615), .Y(n_613) );
AOI322xp5_ASAP7_75t_L g432 ( .A1(n_223), .A2(n_372), .A3(n_410), .B1(n_433), .B2(n_435), .C1(n_436), .C2(n_437), .Y(n_432) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_236), .Y(n_223) );
AND2x2_ASAP7_75t_L g437 ( .A(n_224), .B(n_417), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_224), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g488 ( .A(n_224), .B(n_380), .Y(n_488) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_225), .B(n_285), .Y(n_303) );
AND2x2_ASAP7_75t_L g364 ( .A(n_225), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_225), .B(n_326), .Y(n_408) );
AND2x4_ASAP7_75t_L g445 ( .A(n_225), .B(n_236), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_225), .B(n_367), .Y(n_486) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g275 ( .A(n_226), .B(n_246), .Y(n_275) );
INVx1_ASAP7_75t_L g324 ( .A(n_226), .Y(n_324) );
AND2x2_ASAP7_75t_L g468 ( .A(n_226), .B(n_301), .Y(n_468) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g286 ( .A(n_227), .Y(n_286) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
INVx1_ASAP7_75t_L g295 ( .A(n_229), .Y(n_295) );
OA22x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B1(n_232), .B2(n_234), .Y(n_229) );
INVx4_ASAP7_75t_L g538 ( .A(n_230), .Y(n_538) );
INVx1_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
INVx1_ASAP7_75t_SL g393 ( .A(n_236), .Y(n_393) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
AND2x2_ASAP7_75t_L g285 ( .A(n_237), .B(n_261), .Y(n_285) );
INVx1_ASAP7_75t_L g326 ( .A(n_237), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_237), .B(n_260), .Y(n_502) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
INVx1_ASAP7_75t_L g343 ( .A(n_238), .Y(n_343) );
AND2x2_ASAP7_75t_L g367 ( .A(n_238), .B(n_246), .Y(n_367) );
AND2x2_ASAP7_75t_L g417 ( .A(n_238), .B(n_261), .Y(n_417) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_238), .Y(n_421) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
OR2x2_ASAP7_75t_L g293 ( .A(n_246), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g323 ( .A(n_246), .B(n_324), .Y(n_323) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_255), .Y(n_246) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_247), .A2(n_248), .B(n_255), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_276), .B1(n_283), .B2(n_287), .C(n_289), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_275), .Y(n_258) );
AND2x2_ASAP7_75t_L g463 ( .A(n_259), .B(n_323), .Y(n_463) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g477 ( .A(n_260), .B(n_358), .Y(n_477) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g300 ( .A(n_261), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
AND2x2_ASAP7_75t_L g344 ( .A(n_261), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g366 ( .A(n_261), .Y(n_366) );
BUFx2_ASAP7_75t_L g454 ( .A(n_261), .Y(n_454) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_273), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_275), .A2(n_299), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g466 ( .A(n_275), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_276), .A2(n_313), .B1(n_318), .B2(n_325), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
OR2x2_ASAP7_75t_L g374 ( .A(n_277), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g405 ( .A(n_278), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g423 ( .A(n_278), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g497 ( .A(n_282), .B(n_413), .Y(n_497) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_SL g409 ( .A(n_284), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g385 ( .A(n_286), .B(n_366), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_286), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g472 ( .A(n_286), .Y(n_472) );
OR2x2_ASAP7_75t_L g501 ( .A(n_286), .B(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g469 ( .A(n_287), .B(n_450), .Y(n_469) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI21xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_302), .B(n_304), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_299), .Y(n_291) );
AND2x2_ASAP7_75t_L g325 ( .A(n_292), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g427 ( .A(n_292), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g336 ( .A(n_294), .B(n_337), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_298), .Y(n_294) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g380 ( .A(n_301), .B(n_337), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_302), .A2(n_387), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g480 ( .A(n_306), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g355 ( .A(n_308), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g439 ( .A(n_308), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
INVx1_ASAP7_75t_L g415 ( .A(n_310), .Y(n_415) );
AND2x4_ASAP7_75t_L g434 ( .A(n_310), .B(n_358), .Y(n_434) );
INVx1_ASAP7_75t_SL g481 ( .A(n_310), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_327), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g449 ( .A(n_317), .B(n_450), .Y(n_449) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g433 ( .A(n_320), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_321), .B(n_345), .Y(n_495) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_325), .B(n_346), .Y(n_381) );
AND2x2_ASAP7_75t_L g372 ( .A(n_326), .B(n_336), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_333), .B1(n_339), .B2(n_341), .C1(n_346), .C2(n_355), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI21xp33_ASAP7_75t_L g378 ( .A1(n_329), .A2(n_379), .B(n_381), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_329), .A2(n_447), .B1(n_448), .B2(n_451), .C(n_455), .Y(n_446) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g361 ( .A(n_331), .Y(n_361) );
AND2x2_ASAP7_75t_L g390 ( .A(n_332), .B(n_350), .Y(n_390) );
INVx1_ASAP7_75t_L g414 ( .A(n_332), .Y(n_414) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_332), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_333), .A2(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g457 ( .A(n_336), .B(n_428), .Y(n_457) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g345 ( .A(n_338), .Y(n_345) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
INVx2_ASAP7_75t_L g422 ( .A(n_345), .Y(n_422) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g478 ( .A(n_349), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g444 ( .A(n_350), .Y(n_444) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g578 ( .A(n_354), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_355), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_376), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_368), .C(n_377), .D(n_382), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_361), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_372), .B(n_373), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp33_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_380), .B(n_454), .Y(n_459) );
AND2x4_ASAP7_75t_L g471 ( .A(n_380), .B(n_472), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_380), .B(n_395), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_391), .B2(n_397), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2x1p5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g456 ( .A(n_389), .Y(n_456) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
OR2x2_ASAP7_75t_L g447 ( .A(n_394), .B(n_420), .Y(n_447) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_460), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_425), .C(n_446), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .C(n_416), .Y(n_402) );
AOI22x1_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_409), .B2(n_411), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
OAI21xp33_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_423), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g494 ( .A(n_421), .Y(n_494) );
INVx1_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_424), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_432), .C(n_438), .Y(n_425) );
INVx1_ASAP7_75t_L g467 ( .A(n_428), .Y(n_467) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B(n_445), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_439), .A2(n_457), .B1(n_492), .B2(n_496), .Y(n_491) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_483), .C(n_498), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_470), .Y(n_461) );
OAI31xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .A3(n_468), .B(n_469), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_480), .B2(n_482), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B(n_489), .C(n_491), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g517 ( .A(n_508), .Y(n_517) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
OR2x6_ASAP7_75t_L g892 ( .A(n_511), .B(n_893), .Y(n_892) );
INVx8_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g895 ( .A(n_512), .B(n_896), .Y(n_895) );
OR2x6_ASAP7_75t_L g913 ( .A(n_512), .B(n_896), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_516), .A2(n_519), .B(n_914), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_897), .B1(n_906), .B2(n_910), .C(n_911), .Y(n_519) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_804), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_724), .C(n_768), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_694), .C(n_712), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_648), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_592), .B1(n_637), .B2(n_645), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g780 ( .A(n_528), .Y(n_780) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_562), .Y(n_528) );
NOR2x1p5_ASAP7_75t_L g795 ( .A(n_529), .B(n_700), .Y(n_795) );
NAND2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_545), .Y(n_529) );
INVx2_ASAP7_75t_L g640 ( .A(n_530), .Y(n_640) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g704 ( .A(n_531), .Y(n_704) );
AO31x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_537), .A3(n_543), .B(n_544), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_536), .A2(n_553), .B(n_557), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_538), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g676 ( .A(n_542), .Y(n_676) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_545), .B(n_654), .Y(n_705) );
INVx1_ASAP7_75t_L g755 ( .A(n_545), .Y(n_755) );
AND2x2_ASAP7_75t_L g815 ( .A(n_545), .B(n_642), .Y(n_815) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g653 ( .A(n_546), .Y(n_653) );
AOI21x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_552), .B(n_561), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_549), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AOI21x1_ASAP7_75t_L g642 ( .A1(n_558), .A2(n_643), .B(n_644), .Y(n_642) );
OAI21x1_ASAP7_75t_L g612 ( .A1(n_559), .A2(n_613), .B(n_616), .Y(n_612) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_560), .A2(n_679), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g772 ( .A(n_563), .B(n_703), .Y(n_772) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_579), .Y(n_563) );
AND2x2_ASAP7_75t_L g728 ( .A(n_564), .B(n_704), .Y(n_728) );
INVx1_ASAP7_75t_L g794 ( .A(n_564), .Y(n_794) );
AND2x4_ASAP7_75t_L g802 ( .A(n_564), .B(n_640), .Y(n_802) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_564), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_564), .B(n_857), .Y(n_856) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_565), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g581 ( .A(n_567), .Y(n_581) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_573), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g632 ( .A(n_573), .Y(n_632) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_575), .Y(n_659) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_580), .Y(n_700) );
AND2x2_ASAP7_75t_L g723 ( .A(n_580), .B(n_652), .Y(n_723) );
INVx1_ASAP7_75t_L g851 ( .A(n_580), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_580), .B(n_704), .Y(n_854) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_591), .Y(n_580) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_581), .A2(n_612), .B(n_620), .Y(n_611) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B1(n_589), .B2(n_590), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_587), .A2(n_631), .B(n_635), .Y(n_630) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g644 ( .A(n_591), .Y(n_644) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_610), .Y(n_592) );
OR2x6_ASAP7_75t_L g710 ( .A(n_593), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g822 ( .A(n_593), .B(n_732), .Y(n_822) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g763 ( .A(n_594), .B(n_764), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_594), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g811 ( .A(n_594), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g646 ( .A(n_595), .Y(n_646) );
OR2x2_ASAP7_75t_L g664 ( .A(n_595), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g718 ( .A(n_595), .B(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g737 ( .A(n_595), .B(n_665), .Y(n_737) );
AND2x2_ASAP7_75t_L g787 ( .A(n_595), .B(n_719), .Y(n_787) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_595), .Y(n_865) );
AO31x2_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .A3(n_603), .B(n_608), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_602), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_602), .A2(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_621), .Y(n_610) );
AND2x2_ASAP7_75t_L g647 ( .A(n_611), .B(n_622), .Y(n_647) );
OR2x2_ASAP7_75t_L g770 ( .A(n_611), .B(n_718), .Y(n_770) );
AND2x2_ASAP7_75t_L g812 ( .A(n_611), .B(n_666), .Y(n_812) );
OAI21x1_ASAP7_75t_L g688 ( .A1(n_612), .A2(n_620), .B(n_684), .Y(n_688) );
AND2x2_ASAP7_75t_L g686 ( .A(n_621), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g862 ( .A(n_621), .B(n_646), .Y(n_862) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_622), .B(n_741), .Y(n_740) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g693 ( .A(n_623), .Y(n_693) );
INVx1_ASAP7_75t_L g751 ( .A(n_623), .Y(n_751) );
OA21x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_630), .B(n_636), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g873 ( .A(n_638), .B(n_705), .Y(n_873) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
BUFx2_ASAP7_75t_SL g650 ( .A(n_640), .Y(n_650) );
INVx1_ASAP7_75t_L g716 ( .A(n_640), .Y(n_716) );
AND2x2_ASAP7_75t_L g756 ( .A(n_640), .B(n_654), .Y(n_756) );
AND2x2_ASAP7_75t_L g778 ( .A(n_641), .B(n_767), .Y(n_778) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g758 ( .A(n_642), .B(n_652), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_645), .B(n_797), .Y(n_796) );
INVxp33_ASAP7_75t_L g803 ( .A(n_645), .Y(n_803) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g741 ( .A(n_646), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_646), .Y(n_744) );
OR2x2_ASAP7_75t_L g823 ( .A(n_646), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g872 ( .A(n_646), .B(n_691), .Y(n_872) );
INVx1_ASAP7_75t_L g764 ( .A(n_647), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_661), .Y(n_648) );
INVx1_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
AND2x4_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_651), .B(n_700), .Y(n_747) );
INVx3_ASAP7_75t_L g849 ( .A(n_651), .Y(n_849) );
AND2x4_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g767 ( .A(n_653), .Y(n_767) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_654), .Y(n_890) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_660), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_685), .B(n_689), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g838 ( .A(n_664), .Y(n_838) );
OR2x2_ASAP7_75t_L g869 ( .A(n_664), .B(n_841), .Y(n_869) );
AND2x2_ASAP7_75t_L g692 ( .A(n_665), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_665), .B(n_691), .Y(n_732) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g825 ( .A(n_666), .B(n_687), .Y(n_825) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_674), .B(n_683), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_667), .A2(n_674), .B(n_683), .Y(n_719) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_670), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND3x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .C(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g762 ( .A(n_686), .B(n_737), .Y(n_762) );
INVxp67_ASAP7_75t_L g775 ( .A(n_686), .Y(n_775) );
INVx2_ASAP7_75t_L g691 ( .A(n_687), .Y(n_691) );
AND2x2_ASAP7_75t_L g745 ( .A(n_687), .B(n_693), .Y(n_745) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g781 ( .A(n_689), .Y(n_781) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVx2_ASAP7_75t_L g791 ( .A(n_690), .Y(n_791) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_SL g711 ( .A(n_691), .Y(n_711) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_691), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_692), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g759 ( .A(n_692), .Y(n_759) );
INVx2_ASAP7_75t_SL g709 ( .A(n_693), .Y(n_709) );
BUFx2_ASAP7_75t_L g814 ( .A(n_693), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_699), .B(n_703), .Y(n_783) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g846 ( .A(n_700), .Y(n_846) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
NOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g717 ( .A(n_709), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g786 ( .A(n_709), .Y(n_786) );
AND2x2_ASAP7_75t_L g866 ( .A(n_709), .B(n_825), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_709), .B(n_787), .Y(n_870) );
NOR3xp33_ASAP7_75t_L g889 ( .A(n_709), .B(n_715), .C(n_890), .Y(n_889) );
AND2x2_ASAP7_75t_L g828 ( .A(n_710), .B(n_774), .Y(n_828) );
INVx1_ASAP7_75t_L g736 ( .A(n_711), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_717), .B(n_720), .C(n_722), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g832 ( .A(n_715), .B(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g757 ( .A(n_716), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g777 ( .A(n_716), .B(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_L g800 ( .A(n_718), .B(n_786), .Y(n_800) );
INVx1_ASAP7_75t_L g878 ( .A(n_718), .Y(n_878) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_719), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_722), .A2(n_832), .B1(n_861), .B2(n_863), .C(n_867), .Y(n_860) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g727 ( .A(n_723), .B(n_728), .Y(n_727) );
NOR4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_738), .C(n_748), .D(n_760), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_729), .B1(n_733), .B2(n_734), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_726), .A2(n_739), .B1(n_742), .B2(n_746), .Y(n_738) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI21xp33_ASAP7_75t_SL g807 ( .A1(n_727), .A2(n_808), .B(n_809), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_728), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g784 ( .A(n_728), .Y(n_784) );
AND2x2_ASAP7_75t_L g845 ( .A(n_728), .B(n_846), .Y(n_845) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g840 ( .A(n_731), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g842 ( .A1(n_734), .A2(n_843), .B(n_844), .C(n_847), .Y(n_842) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_737), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g818 ( .A(n_737), .B(n_791), .Y(n_818) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x4_ASAP7_75t_L g858 ( .A(n_744), .B(n_812), .Y(n_858) );
INVx1_ASAP7_75t_L g883 ( .A(n_745), .Y(n_883) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g833 ( .A(n_747), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_757), .B2(n_759), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_750), .B(n_881), .Y(n_880) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_R g841 ( .A(n_751), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_752), .A2(n_800), .B1(n_801), .B2(n_803), .Y(n_799) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
NOR2xp33_ASAP7_75t_SL g891 ( .A(n_754), .B(n_850), .Y(n_891) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g885 ( .A(n_755), .B(n_772), .Y(n_885) );
AND2x4_ASAP7_75t_L g830 ( .A(n_756), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g875 ( .A(n_757), .Y(n_875) );
INVx2_ASAP7_75t_L g831 ( .A(n_758), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_763), .A2(n_828), .B1(n_829), .B2(n_832), .C(n_834), .Y(n_827) );
AND2x2_ASAP7_75t_L g839 ( .A(n_766), .B(n_794), .Y(n_839) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_767), .Y(n_820) );
INVx1_ASAP7_75t_L g857 ( .A(n_767), .Y(n_857) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_788), .C(n_799), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_773), .B2(n_776), .C(n_779), .Y(n_769) );
INVx1_ASAP7_75t_L g874 ( .A(n_770), .Y(n_874) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_774), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_778), .B(n_793), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_782), .B2(n_785), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_789), .B(n_796), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_795), .Y(n_835) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g808 ( .A(n_800), .Y(n_808) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g819 ( .A(n_802), .B(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g826 ( .A(n_802), .B(n_815), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_859), .Y(n_804) );
NOR3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_827), .C(n_842), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_817), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .C(n_816), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_811), .A2(n_819), .B(n_845), .Y(n_844) );
AND2x2_ASAP7_75t_L g886 ( .A(n_812), .B(n_841), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g837 ( .A(n_814), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_821), .B2(n_826), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_830), .A2(n_878), .B1(n_879), .B2(n_882), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_835), .A2(n_836), .B1(n_839), .B2(n_840), .Y(n_834) );
INVx1_ASAP7_75t_L g843 ( .A(n_835), .Y(n_843) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
OAI21xp5_ASAP7_75t_SL g847 ( .A1(n_848), .A2(n_852), .B(n_858), .Y(n_847) );
NOR2x1_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_854), .B(n_856), .Y(n_881) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_876), .Y(n_859) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_868), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .C(n_871), .Y(n_868) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_884), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_891), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_892), .Y(n_907) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx8_ASAP7_75t_L g909 ( .A(n_895), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_897), .Y(n_910) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
BUFx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_913), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
BUFx2_ASAP7_75t_L g924 ( .A(n_918), .Y(n_924) );
BUFx3_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
CKINVDCx16_ASAP7_75t_R g921 ( .A(n_922), .Y(n_921) );
endmodule