module fake_jpeg_19404_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_47),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_54),
.B(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_27),
.B1(n_35),
.B2(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_65),
.B1(n_20),
.B2(n_16),
.Y(n_98)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_27),
.B1(n_35),
.B2(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_72),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_27),
.B1(n_35),
.B2(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_75),
.B1(n_23),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_17),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_18),
.B1(n_23),
.B2(n_36),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_79),
.A2(n_84),
.B1(n_87),
.B2(n_96),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_59),
.B1(n_53),
.B2(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_34),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_21),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_113),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_18),
.B1(n_23),
.B2(n_36),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_28),
.B1(n_30),
.B2(n_21),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_17),
.B1(n_41),
.B2(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_24),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_20),
.B1(n_44),
.B2(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_110),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_41),
.B1(n_38),
.B2(n_21),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_19),
.B1(n_28),
.B2(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_25),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_34),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_34),
.C(n_21),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_126),
.B1(n_129),
.B2(n_133),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_30),
.C(n_31),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_21),
.B1(n_34),
.B2(n_30),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_86),
.B1(n_104),
.B2(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_101),
.C(n_95),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_21),
.B1(n_31),
.B2(n_24),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_24),
.B1(n_31),
.B2(n_2),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_137),
.B1(n_151),
.B2(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_14),
.B(n_13),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_97),
.B1(n_88),
.B2(n_81),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_106),
.B1(n_107),
.B2(n_90),
.Y(n_177)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_91),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_15),
.B(n_12),
.C(n_2),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_12),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_149),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_95),
.B(n_104),
.C(n_80),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_166),
.B(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_104),
.B1(n_101),
.B2(n_96),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_184),
.B1(n_185),
.B2(n_5),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_161),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_100),
.C(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_163),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_120),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_112),
.C(n_77),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_7),
.C(n_8),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_169),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_102),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_139),
.B(n_127),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_1),
.B(n_3),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_102),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_119),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_139),
.B1(n_133),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_125),
.B1(n_134),
.B2(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_138),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_12),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_148),
.B1(n_141),
.B2(n_130),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_195),
.B1(n_199),
.B2(n_204),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_191),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_142),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_142),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_193),
.B(n_197),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_124),
.B(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_149),
.B1(n_135),
.B2(n_131),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_3),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_170),
.B(n_153),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_161),
.B(n_166),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_135),
.B1(n_131),
.B2(n_7),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_152),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_179),
.B(n_182),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_159),
.A2(n_135),
.B1(n_6),
.B2(n_7),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_172),
.B1(n_191),
.B2(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_184),
.C(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_156),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_229),
.B1(n_187),
.B2(n_199),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_178),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_215),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_219),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_158),
.B1(n_177),
.B2(n_156),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_182),
.B1(n_185),
.B2(n_181),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_208),
.B1(n_197),
.B2(n_204),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_181),
.B1(n_183),
.B2(n_168),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_9),
.C(n_10),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_241),
.C(n_243),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_9),
.B1(n_10),
.B2(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_188),
.C(n_209),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_10),
.C(n_188),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_205),
.B(n_207),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_259),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_253),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_196),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_264),
.B1(n_235),
.B2(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_205),
.B1(n_190),
.B2(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_186),
.B1(n_216),
.B2(n_212),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_264),
.B1(n_253),
.B2(n_257),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_244),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_221),
.B(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_248),
.B1(n_246),
.B2(n_221),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_222),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_241),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_227),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_283),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_218),
.C(n_243),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_273),
.B1(n_265),
.B2(n_262),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_267),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_251),
.B1(n_256),
.B2(n_259),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_245),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_294),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_251),
.B1(n_218),
.B2(n_186),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_245),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_244),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_245),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.C(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_247),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_277),
.C(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_278),
.C(n_274),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_294),
.C(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_234),
.C(n_282),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_282),
.C(n_194),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_286),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_314),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_295),
.B(n_293),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_194),
.B1(n_265),
.B2(n_284),
.C(n_255),
.Y(n_314)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_275),
.C(n_269),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_275),
.C(n_269),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_321),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_260),
.C(n_249),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_308),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_320),
.B(n_201),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.B(n_324),
.C(n_270),
.D(n_254),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_319),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_201),
.C(n_239),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_239),
.B1(n_213),
.B2(n_210),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_193),
.B(n_237),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_233),
.C(n_210),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_233),
.B(n_10),
.Y(n_332)
);


endmodule