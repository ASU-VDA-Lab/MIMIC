module fake_jpeg_15676_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_19),
.B1(n_15),
.B2(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_25),
.B1(n_18),
.B2(n_5),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_14),
.B1(n_5),
.B2(n_0),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_39),
.B2(n_29),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_39),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_29),
.B1(n_22),
.B2(n_37),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_47),
.Y(n_53)
);


endmodule