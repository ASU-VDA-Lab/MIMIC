module real_aes_2095_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_0), .B(n_115), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_1), .A2(n_128), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_2), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_3), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g122 ( .A(n_4), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_5), .B(n_137), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_6), .B(n_124), .Y(n_497) );
INVx1_ASAP7_75t_L g473 ( .A(n_7), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g830 ( .A(n_8), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_9), .Y(n_488) );
NAND2xp33_ASAP7_75t_L g200 ( .A(n_10), .B(n_135), .Y(n_200) );
INVx2_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
AOI221x1_ASAP7_75t_L g144 ( .A1(n_12), .A2(n_24), .B1(n_115), .B2(n_128), .C(n_145), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_13), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_14), .B(n_115), .Y(n_196) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_15), .A2(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g505 ( .A(n_16), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_17), .B(n_142), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_18), .B(n_137), .Y(n_188) );
AO21x1_ASAP7_75t_L g114 ( .A1(n_19), .A2(n_115), .B(n_123), .Y(n_114) );
INVx1_ASAP7_75t_L g438 ( .A(n_20), .Y(n_438) );
INVx1_ASAP7_75t_L g503 ( .A(n_21), .Y(n_503) );
INVx1_ASAP7_75t_SL g554 ( .A(n_22), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_23), .B(n_116), .Y(n_517) );
NAND2x1_ASAP7_75t_L g155 ( .A(n_25), .B(n_137), .Y(n_155) );
AOI33xp33_ASAP7_75t_L g541 ( .A1(n_26), .A2(n_52), .A3(n_454), .B1(n_461), .B2(n_542), .B3(n_543), .Y(n_541) );
NAND2x1_ASAP7_75t_L g214 ( .A(n_27), .B(n_135), .Y(n_214) );
INVx1_ASAP7_75t_L g481 ( .A(n_28), .Y(n_481) );
OR2x2_ASAP7_75t_L g125 ( .A(n_29), .B(n_86), .Y(n_125) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_29), .A2(n_86), .B(n_126), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_30), .B(n_452), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_31), .B(n_135), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_32), .B(n_137), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_33), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_34), .A2(n_128), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g799 ( .A(n_35), .Y(n_799) );
AND2x2_ASAP7_75t_L g121 ( .A(n_36), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g129 ( .A(n_36), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g460 ( .A(n_36), .Y(n_460) );
OR2x6_ASAP7_75t_L g436 ( .A(n_37), .B(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_38), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_39), .B(n_115), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_40), .B(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_124), .B1(n_160), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_42), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_43), .B(n_116), .Y(n_555) );
OAI222xp33_ASAP7_75t_L g101 ( .A1(n_44), .A2(n_102), .B1(n_103), .B2(n_790), .C1(n_796), .C2(n_799), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_44), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_45), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_46), .B(n_135), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_47), .B(n_194), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_48), .B(n_116), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_49), .A2(n_128), .B(n_213), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_50), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_51), .B(n_135), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_53), .B(n_116), .Y(n_466) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
INVx1_ASAP7_75t_L g132 ( .A(n_54), .Y(n_132) );
AND2x2_ASAP7_75t_L g467 ( .A(n_55), .B(n_142), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_56), .A2(n_75), .B1(n_452), .B2(n_458), .C(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_57), .B(n_452), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_58), .B(n_137), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_59), .B(n_160), .Y(n_490) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_60), .A2(n_458), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_61), .A2(n_128), .B(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_62), .A2(n_106), .B1(n_819), .B2(n_820), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_62), .Y(n_820) );
INVx1_ASAP7_75t_L g500 ( .A(n_63), .Y(n_500) );
AO21x1_ASAP7_75t_L g127 ( .A1(n_64), .A2(n_128), .B(n_133), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_65), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_66), .B(n_115), .Y(n_205) );
INVx1_ASAP7_75t_L g464 ( .A(n_67), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_68), .B(n_115), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_69), .A2(n_458), .B(n_463), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_70), .Y(n_832) );
AND2x2_ASAP7_75t_L g172 ( .A(n_71), .B(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g130 ( .A(n_72), .Y(n_130) );
AND2x2_ASAP7_75t_L g218 ( .A(n_73), .B(n_159), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_74), .B(n_452), .Y(n_544) );
AND2x2_ASAP7_75t_L g556 ( .A(n_76), .B(n_159), .Y(n_556) );
INVx1_ASAP7_75t_L g501 ( .A(n_77), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_78), .A2(n_458), .B(n_553), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_79), .A2(n_458), .B(n_516), .C(n_520), .Y(n_515) );
INVx1_ASAP7_75t_L g439 ( .A(n_80), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_81), .B(n_115), .Y(n_190) );
AND2x2_ASAP7_75t_L g203 ( .A(n_82), .B(n_159), .Y(n_203) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_83), .B(n_159), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_84), .A2(n_458), .B1(n_539), .B2(n_540), .Y(n_538) );
AND2x2_ASAP7_75t_L g123 ( .A(n_85), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g162 ( .A(n_87), .B(n_159), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_88), .B(n_135), .Y(n_189) );
INVx1_ASAP7_75t_L g527 ( .A(n_89), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_90), .B(n_137), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_91), .B(n_135), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_92), .A2(n_128), .B(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g545 ( .A(n_93), .B(n_159), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_94), .B(n_137), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_95), .A2(n_479), .B(n_480), .C(n_483), .Y(n_478) );
BUFx2_ASAP7_75t_L g803 ( .A(n_96), .Y(n_803) );
BUFx2_ASAP7_75t_SL g816 ( .A(n_96), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_97), .A2(n_128), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_98), .B(n_116), .Y(n_528) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_824), .B(n_831), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_800), .B(n_812), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_431), .B1(n_440), .B2(n_786), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_106), .A2(n_792), .B1(n_794), .B2(n_795), .Y(n_791) );
INVx1_ASAP7_75t_L g819 ( .A(n_106), .Y(n_819) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_330), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_267), .C(n_290), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_219), .C(n_236), .Y(n_108) );
OAI31xp33_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_149), .A3(n_173), .B(n_180), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_110), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_141), .Y(n_111) );
AND2x4_ASAP7_75t_L g222 ( .A(n_112), .B(n_141), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_112), .B(n_164), .Y(n_251) );
AND2x4_ASAP7_75t_L g253 ( .A(n_112), .B(n_247), .Y(n_253) );
AND2x2_ASAP7_75t_L g384 ( .A(n_112), .B(n_177), .Y(n_384) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g229 ( .A(n_113), .Y(n_229) );
OAI21x1_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_127), .B(n_139), .Y(n_113) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_121), .Y(n_115) );
INVx1_ASAP7_75t_L g482 ( .A(n_116), .Y(n_482) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
AND2x6_ASAP7_75t_L g135 ( .A(n_117), .B(n_130), .Y(n_135) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g137 ( .A(n_119), .B(n_132), .Y(n_137) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx5_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_121), .Y(n_483) );
AND2x2_ASAP7_75t_L g131 ( .A(n_122), .B(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_122), .Y(n_455) );
INVx1_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_124), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_SL g184 ( .A(n_124), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_124), .A2(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_124), .B(n_138), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_124), .A2(n_525), .B(n_529), .Y(n_524) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_125), .B(n_126), .Y(n_143) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
BUFx3_ASAP7_75t_L g456 ( .A(n_129), .Y(n_456) );
INVx2_ASAP7_75t_L g462 ( .A(n_130), .Y(n_462) );
AND2x4_ASAP7_75t_L g458 ( .A(n_131), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g454 ( .A(n_132), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_136), .B(n_138), .Y(n_133) );
INVxp67_ASAP7_75t_L g504 ( .A(n_135), .Y(n_504) );
INVxp67_ASAP7_75t_L g506 ( .A(n_137), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_138), .A2(n_146), .B(n_147), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_138), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_138), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_138), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_138), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_138), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_138), .A2(n_214), .B(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_138), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_138), .A2(n_465), .B(n_473), .C(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_138), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_138), .A2(n_465), .B(n_527), .C(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g539 ( .A(n_138), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_138), .A2(n_465), .B(n_554), .C(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g163 ( .A(n_141), .B(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_141), .B(n_228), .Y(n_320) );
AND2x2_ASAP7_75t_L g326 ( .A(n_141), .B(n_165), .Y(n_326) );
AND2x2_ASAP7_75t_L g415 ( .A(n_141), .B(n_416), .Y(n_415) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_148), .Y(n_141) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_142), .A2(n_144), .B(n_148), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_142), .A2(n_205), .B(n_206), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_142), .Y(n_217) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_SL g397 ( .A(n_149), .Y(n_397) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_163), .Y(n_149) );
BUFx2_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
AND2x2_ASAP7_75t_L g260 ( .A(n_150), .B(n_164), .Y(n_260) );
AND2x2_ASAP7_75t_L g309 ( .A(n_150), .B(n_165), .Y(n_309) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g266 ( .A(n_151), .B(n_165), .Y(n_266) );
INVxp67_ASAP7_75t_L g278 ( .A(n_151), .Y(n_278) );
BUFx3_ASAP7_75t_L g323 ( .A(n_151), .Y(n_323) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_158), .B(n_162), .Y(n_151) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_158), .B(n_162), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_158), .A2(n_166), .B(n_172), .Y(n_165) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_158), .A2(n_166), .B(n_172), .Y(n_179) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_158), .A2(n_450), .B(n_467), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_158), .A2(n_159), .B1(n_478), .B2(n_484), .Y(n_477) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_158), .A2(n_450), .B(n_467), .Y(n_606) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_160), .B(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
OAI31xp33_ASAP7_75t_L g219 ( .A1(n_163), .A2(n_220), .A3(n_225), .B(n_230), .Y(n_219) );
AND2x2_ASAP7_75t_L g227 ( .A(n_164), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g246 ( .A(n_165), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_167), .B(n_171), .Y(n_166) );
AOI322xp5_ASAP7_75t_L g420 ( .A1(n_173), .A2(n_295), .A3(n_324), .B1(n_329), .B2(n_421), .C1(n_424), .C2(n_425), .Y(n_420) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_176), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_174), .B(n_266), .Y(n_271) );
NAND2x1_ASAP7_75t_L g308 ( .A(n_174), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g352 ( .A(n_174), .B(n_256), .Y(n_352) );
INVx1_ASAP7_75t_SL g366 ( .A(n_174), .Y(n_366) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_175), .Y(n_390) );
AND2x2_ASAP7_75t_L g319 ( .A(n_176), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_176), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_177), .B(n_178), .Y(n_176) );
BUFx2_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
INVx1_ASAP7_75t_L g416 ( .A(n_177), .Y(n_416) );
OR2x2_ASAP7_75t_L g283 ( .A(n_178), .B(n_228), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_178), .B(n_253), .Y(n_317) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g256 ( .A(n_179), .B(n_228), .Y(n_256) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_201), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g312 ( .A(n_182), .Y(n_312) );
OR2x2_ASAP7_75t_L g339 ( .A(n_182), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
NOR2x1_ASAP7_75t_SL g233 ( .A(n_183), .B(n_202), .Y(n_233) );
AND2x2_ASAP7_75t_L g240 ( .A(n_183), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g412 ( .A(n_183), .B(n_274), .Y(n_412) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_184), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
OR2x2_ASAP7_75t_L g234 ( .A(n_193), .B(n_235), .Y(n_234) );
BUFx3_ASAP7_75t_L g243 ( .A(n_193), .Y(n_243) );
INVx2_ASAP7_75t_L g274 ( .A(n_193), .Y(n_274) );
INVx1_ASAP7_75t_L g315 ( .A(n_193), .Y(n_315) );
AND2x2_ASAP7_75t_L g346 ( .A(n_193), .B(n_202), .Y(n_346) );
AND2x2_ASAP7_75t_L g377 ( .A(n_193), .B(n_304), .Y(n_377) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_194), .A2(n_471), .B(n_475), .Y(n_470) );
INVx2_ASAP7_75t_SL g520 ( .A(n_194), .Y(n_520) );
AND2x2_ASAP7_75t_L g273 ( .A(n_201), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_201), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_201), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g381 ( .A(n_201), .B(n_243), .Y(n_381) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
INVx5_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_202), .B(n_235), .Y(n_313) );
BUFx2_ASAP7_75t_L g373 ( .A(n_202), .Y(n_373) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx4_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
AND2x2_ASAP7_75t_L g358 ( .A(n_210), .B(n_241), .Y(n_358) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_217), .A2(n_550), .B(n_556), .Y(n_549) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_221), .A2(n_348), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g369 ( .A(n_222), .B(n_260), .Y(n_369) );
INVx1_ASAP7_75t_SL g395 ( .A(n_222), .Y(n_395) );
AND2x2_ASAP7_75t_L g380 ( .A(n_223), .B(n_352), .Y(n_380) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_224), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
AND2x2_ASAP7_75t_L g249 ( .A(n_226), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g255 ( .A(n_226), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
AND2x2_ASAP7_75t_L g337 ( .A(n_227), .B(n_265), .Y(n_337) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
OR2x2_ASAP7_75t_L g426 ( .A(n_234), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g242 ( .A(n_235), .Y(n_242) );
AND2x4_ASAP7_75t_L g298 ( .A(n_235), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_235), .B(n_303), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_235), .B(n_241), .Y(n_340) );
AND2x2_ASAP7_75t_L g400 ( .A(n_235), .B(n_303), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_244), .B1(n_257), .B2(n_259), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_237), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND3x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .C(n_243), .Y(n_239) );
AND2x4_ASAP7_75t_L g257 ( .A(n_240), .B(n_258), .Y(n_257) );
INVx4_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_241), .B(n_298), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_242), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g342 ( .A(n_243), .Y(n_342) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_243), .A2(n_372), .A3(n_408), .B1(n_410), .B2(n_413), .C1(n_417), .C2(n_418), .Y(n_407) );
NAND4xp25_ASAP7_75t_SL g244 ( .A(n_245), .B(n_248), .C(n_252), .D(n_254), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_246), .B(n_262), .Y(n_374) );
BUFx2_ASAP7_75t_L g265 ( .A(n_247), .Y(n_265) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g389 ( .A(n_250), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g403 ( .A(n_251), .B(n_278), .Y(n_403) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g269 ( .A(n_253), .B(n_270), .Y(n_269) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_253), .A2(n_322), .B(n_324), .C(n_327), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_253), .B(n_260), .Y(n_379) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_255), .A2(n_337), .B1(n_338), .B2(n_341), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_256), .A2(n_292), .B1(n_296), .B2(n_300), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_256), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_256), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_256), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g423 ( .A(n_256), .Y(n_423) );
INVx1_ASAP7_75t_L g362 ( .A(n_257), .Y(n_362) );
OAI21xp33_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_261), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g270 ( .A(n_260), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_260), .B(n_265), .Y(n_419) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g355 ( .A(n_262), .B(n_266), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_264), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g422 ( .A(n_265), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g396 ( .A(n_266), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_272), .C(n_275), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_270), .A2(n_301), .B1(n_348), .B2(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_274), .B(n_297), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_274), .B(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_280), .B(n_284), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI211xp5_ASAP7_75t_SL g333 ( .A1(n_281), .A2(n_334), .B(n_336), .C(n_344), .Y(n_333) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp67_ASAP7_75t_SL g367 ( .A(n_286), .B(n_313), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_286), .Y(n_370) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_288), .B(n_297), .Y(n_427) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g299 ( .A(n_289), .Y(n_299) );
INVx2_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
NAND4xp25_ASAP7_75t_L g290 ( .A(n_291), .B(n_306), .C(n_318), .D(n_321), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_294), .A2(n_426), .B1(n_428), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x4_ASAP7_75t_L g393 ( .A(n_297), .B(n_323), .Y(n_393) );
AND2x2_ASAP7_75t_L g314 ( .A(n_298), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
AND2x2_ASAP7_75t_L g345 ( .A(n_298), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
INVx1_ASAP7_75t_L g349 ( .A(n_305), .Y(n_349) );
AOI32xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .A3(n_313), .B1(n_314), .B2(n_316), .Y(n_306) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_307), .A2(n_355), .B(n_356), .Y(n_354) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_310), .A2(n_387), .B1(n_389), .B2(n_391), .C(n_394), .Y(n_386) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g371 ( .A(n_312), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g329 ( .A(n_313), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_314), .A2(n_352), .B1(n_402), .B2(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
AND2x2_ASAP7_75t_L g406 ( .A(n_315), .B(n_359), .Y(n_406) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_322), .B(n_374), .Y(n_409) );
INVx1_ASAP7_75t_L g428 ( .A(n_322), .Y(n_428) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g330 ( .A(n_331), .B(n_385), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_375), .Y(n_331) );
NOR3xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_347), .C(n_360), .Y(n_332) );
INVx1_ASAP7_75t_L g350 ( .A(n_335), .Y(n_350) );
INVx1_ASAP7_75t_SL g361 ( .A(n_337), .Y(n_361) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g343 ( .A(n_340), .Y(n_343) );
INVx2_ASAP7_75t_L g353 ( .A(n_341), .Y(n_353) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x4_ASAP7_75t_L g399 ( .A(n_342), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g417 ( .A(n_346), .B(n_400), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g368 ( .A1(n_357), .A2(n_369), .A3(n_370), .B1(n_371), .B2(n_374), .Y(n_368) );
NOR2xp33_ASAP7_75t_SL g387 ( .A(n_357), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g388 ( .A(n_359), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B(n_363), .C(n_368), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_412), .Y(n_424) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_373), .B(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_380), .B2(n_381), .C(n_382), .Y(n_375) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
CKINVDCx16_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_401), .C(n_407), .D(n_420), .Y(n_385) );
INVxp33_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_397), .C(n_398), .Y(n_394) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
CKINVDCx11_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
INVx4_ASAP7_75t_SL g795 ( .A(n_432), .Y(n_795) );
INVx3_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
AND2x6_ASAP7_75t_SL g434 ( .A(n_435), .B(n_436), .Y(n_434) );
OR2x6_ASAP7_75t_SL g788 ( .A(n_435), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g798 ( .A(n_435), .B(n_436), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_435), .B(n_789), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_436), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g794 ( .A(n_440), .Y(n_794) );
NAND4xp75_ASAP7_75t_L g440 ( .A(n_441), .B(n_658), .C(n_703), .D(n_772), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_618), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_574), .C(n_599), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_492), .B1(n_530), .B2(n_546), .C1(n_561), .C2(n_568), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_468), .Y(n_446) );
AND2x2_ASAP7_75t_L g783 ( .A(n_447), .B(n_597), .Y(n_783) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_449), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_449), .B(n_476), .Y(n_573) );
INVx3_ASAP7_75t_L g588 ( .A(n_449), .Y(n_588) );
AND2x2_ASAP7_75t_L g721 ( .A(n_449), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g491 ( .A(n_452), .Y(n_491) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g512 ( .A(n_453), .Y(n_512) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
OR2x6_ASAP7_75t_L g465 ( .A(n_454), .B(n_462), .Y(n_465) );
INVxp33_ASAP7_75t_L g542 ( .A(n_454), .Y(n_542) );
INVx1_ASAP7_75t_L g513 ( .A(n_456), .Y(n_513) );
INVxp67_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
NOR2x1p5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g543 ( .A(n_461), .Y(n_543) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_465), .A2(n_482), .B1(n_500), .B2(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
AND2x2_ASAP7_75t_L g651 ( .A(n_468), .B(n_604), .Y(n_651) );
AND2x2_ASAP7_75t_L g653 ( .A(n_468), .B(n_654), .Y(n_653) );
INVx3_ASAP7_75t_L g688 ( .A(n_468), .Y(n_688) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_476), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g571 ( .A(n_470), .Y(n_571) );
INVx1_ASAP7_75t_L g590 ( .A(n_470), .Y(n_590) );
AND2x4_ASAP7_75t_L g597 ( .A(n_470), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_470), .B(n_536), .Y(n_613) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_470), .Y(n_722) );
INVx1_ASAP7_75t_L g732 ( .A(n_470), .Y(n_732) );
INVx1_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
INVx2_ASAP7_75t_L g585 ( .A(n_476), .Y(n_585) );
INVx1_ASAP7_75t_L g666 ( .A(n_476), .Y(n_666) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_494), .B(n_521), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_494), .B(n_548), .Y(n_641) );
INVx2_ASAP7_75t_L g662 ( .A(n_494), .Y(n_662) );
AND2x2_ASAP7_75t_L g670 ( .A(n_494), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_508), .Y(n_494) );
AND2x4_ASAP7_75t_L g560 ( .A(n_495), .B(n_509), .Y(n_560) );
INVx1_ASAP7_75t_L g567 ( .A(n_495), .Y(n_567) );
AND2x2_ASAP7_75t_L g743 ( .A(n_495), .B(n_549), .Y(n_743) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g581 ( .A(n_496), .B(n_509), .Y(n_581) );
INVx2_ASAP7_75t_L g617 ( .A(n_496), .Y(n_617) );
AND2x2_ASAP7_75t_L g696 ( .A(n_496), .B(n_549), .Y(n_696) );
NOR2x1_ASAP7_75t_SL g739 ( .A(n_496), .B(n_522), .Y(n_739) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B(n_507), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g579 ( .A(n_508), .Y(n_579) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g593 ( .A(n_509), .B(n_522), .Y(n_593) );
INVx1_ASAP7_75t_L g609 ( .A(n_509), .Y(n_609) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_509), .Y(n_717) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .C(n_514), .Y(n_511) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_520), .A2(n_537), .B(n_545), .Y(n_536) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_520), .A2(n_537), .B(n_545), .Y(n_586) );
AND2x2_ASAP7_75t_L g580 ( .A(n_521), .B(n_581), .Y(n_580) );
OR2x6_ASAP7_75t_L g661 ( .A(n_521), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g699 ( .A(n_521), .B(n_696), .Y(n_699) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_522), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g628 ( .A(n_522), .Y(n_628) );
OR2x2_ASAP7_75t_L g634 ( .A(n_522), .B(n_549), .Y(n_634) );
AND2x4_ASAP7_75t_L g648 ( .A(n_522), .B(n_609), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_522), .B(n_617), .Y(n_649) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g693 ( .A(n_533), .B(n_612), .Y(n_693) );
BUFx2_ASAP7_75t_L g745 ( .A(n_533), .Y(n_745) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g776 ( .A(n_535), .B(n_688), .Y(n_776) );
INVx2_ASAP7_75t_L g570 ( .A(n_536), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_544), .Y(n_537) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_557), .Y(n_546) );
AND2x2_ASAP7_75t_L g592 ( .A(n_547), .B(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_SL g577 ( .A(n_548), .B(n_567), .Y(n_577) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g565 ( .A(n_549), .Y(n_565) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_549), .Y(n_671) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_549), .Y(n_738) );
INVx1_ASAP7_75t_L g778 ( .A(n_549), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
BUFx2_ASAP7_75t_L g692 ( .A(n_557), .Y(n_692) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x4_ASAP7_75t_L g608 ( .A(n_558), .B(n_609), .Y(n_608) );
NOR2xp67_ASAP7_75t_SL g640 ( .A(n_558), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g713 ( .A(n_558), .B(n_696), .Y(n_713) );
AND2x4_ASAP7_75t_SL g716 ( .A(n_558), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g765 ( .A(n_558), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g632 ( .A(n_559), .Y(n_632) );
INVx4_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g627 ( .A(n_560), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_560), .B(n_625), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_560), .B(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_560), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g710 ( .A(n_564), .B(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
AND2x2_ASAP7_75t_L g744 ( .A(n_569), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g752 ( .A(n_569), .B(n_681), .Y(n_752) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g621 ( .A(n_570), .B(n_606), .Y(n_621) );
AND2x4_ASAP7_75t_L g654 ( .A(n_570), .B(n_588), .Y(n_654) );
INVx1_ASAP7_75t_L g771 ( .A(n_570), .Y(n_771) );
AND2x2_ASAP7_75t_L g657 ( .A(n_572), .B(n_597), .Y(n_657) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g678 ( .A(n_573), .B(n_613), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_582), .B1(n_591), .B2(n_594), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B(n_580), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_576), .A2(n_645), .B1(n_753), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_577), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g646 ( .A(n_577), .B(n_578), .Y(n_646) );
AND2x2_ASAP7_75t_SL g676 ( .A(n_577), .B(n_648), .Y(n_676) );
AOI211xp5_ASAP7_75t_SL g764 ( .A1(n_577), .A2(n_765), .B(n_767), .C(n_768), .Y(n_764) );
AND2x2_ASAP7_75t_SL g695 ( .A(n_578), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_578), .B(n_624), .Y(n_750) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g655 ( .A(n_580), .Y(n_655) );
INVx2_ASAP7_75t_L g711 ( .A(n_581), .Y(n_711) );
AND2x2_ASAP7_75t_L g785 ( .A(n_581), .B(n_778), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_582), .A2(n_734), .B(n_740), .Y(n_733) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g720 ( .A(n_584), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g730 ( .A(n_584), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AND2x2_ASAP7_75t_L g637 ( .A(n_585), .B(n_590), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_585), .B(n_606), .Y(n_639) );
AND2x2_ASAP7_75t_L g681 ( .A(n_585), .B(n_606), .Y(n_681) );
INVx2_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
AND2x4_ASAP7_75t_L g604 ( .A(n_586), .B(n_605), .Y(n_604) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx3_ASAP7_75t_L g596 ( .A(n_588), .Y(n_596) );
INVx3_ASAP7_75t_L g602 ( .A(n_589), .Y(n_602) );
BUFx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_593), .A2(n_699), .B(n_775), .Y(n_779) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g611 ( .A(n_596), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_596), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_596), .B(n_671), .Y(n_686) );
OR2x2_ASAP7_75t_L g701 ( .A(n_596), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g708 ( .A(n_596), .B(n_612), .Y(n_708) );
AND2x2_ASAP7_75t_L g664 ( .A(n_597), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g680 ( .A(n_597), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g697 ( .A(n_597), .B(n_666), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_607), .B1(n_610), .B2(n_614), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_602), .B(n_603), .Y(n_674) );
NOR2xp67_ASAP7_75t_SL g712 ( .A(n_602), .B(n_620), .Y(n_712) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_606), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g615 ( .A(n_608), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g679 ( .A(n_608), .B(n_625), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_608), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g782 ( .A(n_616), .B(n_648), .Y(n_782) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_617), .B(n_728), .Y(n_727) );
NOR2xp67_ASAP7_75t_SL g618 ( .A(n_619), .B(n_642), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B(n_629), .C(n_638), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_620), .A2(n_673), .B(n_683), .C(n_687), .Y(n_682) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g762 ( .A(n_621), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g673 ( .A(n_625), .B(n_649), .Y(n_673) );
AND2x2_ASAP7_75t_L g760 ( .A(n_625), .B(n_739), .Y(n_760) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g728 ( .A(n_628), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_632), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g702 ( .A(n_637), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_650), .B1(n_652), .B2(n_655), .C(n_656), .Y(n_642) );
NOR4xp25_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .C(n_647), .D(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g761 ( .A(n_648), .B(n_724), .Y(n_761) );
INVx2_ASAP7_75t_L g767 ( .A(n_648), .Y(n_767) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_651), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g754 ( .A(n_654), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND4xp75_ASAP7_75t_L g659 ( .A(n_660), .B(n_682), .C(n_689), .D(n_698), .Y(n_659) );
OA211x2_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B(n_667), .C(n_675), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_661), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g755 ( .A(n_665), .Y(n_755) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g763 ( .A(n_666), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_674), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g724 ( .A(n_671), .Y(n_724) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g784 ( .A1(n_679), .A2(n_730), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g758 ( .A(n_680), .Y(n_758) );
NAND2x1p5_ASAP7_75t_L g770 ( .A(n_681), .B(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_694), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVxp67_ASAP7_75t_L g756 ( .A(n_692), .Y(n_756) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_696), .B(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_697), .A2(n_760), .B1(n_782), .B2(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND3x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_746), .C(n_759), .Y(n_704) );
NOR3x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_718), .C(n_733), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_714), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_712), .B2(n_713), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_723), .B1(n_725), .B2(n_729), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g777 ( .A(n_727), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .Y(n_740) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g766 ( .A(n_743), .Y(n_766) );
OAI21xp5_ASAP7_75t_SL g774 ( .A1(n_744), .A2(n_775), .B(n_777), .Y(n_774) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_757), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B1(n_753), .B2(n_756), .Y(n_747) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
O2A1O1Ixp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B(n_762), .C(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NOR2x1_ASAP7_75t_SL g772 ( .A(n_773), .B(n_780), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_779), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_781), .B(n_784), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_787), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
BUFx4f_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_797), .B(n_828), .Y(n_827) );
INVx3_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_804), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
INVxp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_805), .A2(n_818), .B(n_821), .Y(n_817) );
NOR2xp33_ASAP7_75t_SL g805 ( .A(n_806), .B(n_811), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx2_ASAP7_75t_R g823 ( .A(n_810), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g833 ( .A(n_827), .Y(n_833) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
endmodule