module fake_jpeg_11579_n_560 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_560);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_560;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_65),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_64),
.Y(n_139)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_68),
.Y(n_175)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_75),
.Y(n_182)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_98),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_86),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_90),
.Y(n_166)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_32),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_97),
.Y(n_169)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_15),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_23),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_99),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_107),
.Y(n_181)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_32),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_119),
.Y(n_190)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_44),
.B(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_3),
.Y(n_180)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_28),
.B(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_48),
.Y(n_159)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_20),
.B1(n_42),
.B2(n_59),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_124),
.A2(n_133),
.B1(n_142),
.B2(n_153),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_54),
.B1(n_59),
.B2(n_42),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_127),
.A2(n_150),
.B1(n_173),
.B2(n_177),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_20),
.B1(n_45),
.B2(n_47),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_57),
.B(n_4),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_134),
.A2(n_100),
.A3(n_78),
.B1(n_15),
.B2(n_103),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_47),
.C(n_37),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_137),
.A2(n_68),
.B(n_78),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_45),
.B1(n_55),
.B2(n_50),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_67),
.A2(n_58),
.B1(n_56),
.B2(n_52),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_152),
.A2(n_192),
.B1(n_115),
.B2(n_114),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_70),
.A2(n_56),
.B1(n_30),
.B2(n_52),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_72),
.A2(n_55),
.B1(n_50),
.B2(n_21),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_157),
.A2(n_163),
.B1(n_170),
.B2(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_159),
.B(n_195),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_74),
.A2(n_40),
.B1(n_37),
.B2(n_21),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_40),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_75),
.A2(n_48),
.B1(n_34),
.B2(n_33),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_69),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_180),
.B(n_165),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_188),
.B1(n_112),
.B2(n_108),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_86),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_79),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_111),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_204),
.B(n_234),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_206),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_207),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_218),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_95),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_258),
.C(n_260),
.Y(n_291)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_210),
.Y(n_300)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_228),
.Y(n_288)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_213),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_102),
.B1(n_118),
.B2(n_105),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_145),
.Y(n_216)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_217),
.A2(n_266),
.B1(n_269),
.B2(n_271),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_169),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_135),
.B(n_63),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_12),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_221),
.B(n_222),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_14),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_164),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_79),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_240),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_225),
.A2(n_226),
.B1(n_251),
.B2(n_253),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_157),
.A2(n_89),
.B1(n_94),
.B2(n_106),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_162),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_257),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_162),
.Y(n_234)
);

BUFx12_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_235),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_173),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_238),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_127),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_168),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_131),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_163),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_243),
.B(n_244),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_130),
.B(n_100),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_85),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_265),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_146),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_248),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_155),
.B(n_126),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_149),
.Y(n_249)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_249),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_154),
.B(n_189),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_253),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_133),
.A2(n_129),
.B1(n_160),
.B2(n_136),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_156),
.B(n_200),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_256),
.Y(n_308)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_255),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_175),
.B(n_179),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_132),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_261),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_179),
.B(n_158),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_264),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_165),
.B(n_174),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_183),
.C(n_187),
.Y(n_293)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_144),
.B(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_129),
.B(n_136),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_267),
.B(n_214),
.Y(n_302)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_268),
.Y(n_314)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_174),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_188),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_285),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_204),
.A2(n_185),
.B(n_177),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_280),
.A2(n_306),
.B(n_231),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_143),
.B1(n_178),
.B2(n_182),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_284),
.A2(n_286),
.B1(n_299),
.B2(n_305),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_245),
.A2(n_143),
.B1(n_178),
.B2(n_182),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_245),
.A2(n_187),
.B1(n_183),
.B2(n_164),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_318),
.B1(n_320),
.B2(n_327),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_214),
.A2(n_267),
.B1(n_209),
.B2(n_221),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_205),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_228),
.A2(n_209),
.B1(n_202),
.B2(n_222),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_244),
.A2(n_220),
.B1(n_242),
.B2(n_264),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_236),
.A2(n_263),
.B1(n_260),
.B2(n_223),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_263),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_313),
.B(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_268),
.A2(n_232),
.B1(n_206),
.B2(n_213),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_216),
.A2(n_266),
.B1(n_241),
.B2(n_256),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_258),
.B(n_210),
.CI(n_260),
.CON(n_321),
.SN(n_321)
);

MAJIxp5_ASAP7_75t_SL g369 ( 
.A(n_321),
.B(n_273),
.C(n_291),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_270),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_233),
.A2(n_259),
.B1(n_239),
.B2(n_230),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_255),
.B1(n_249),
.B2(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_212),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_331),
.B(n_346),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_332),
.B(n_368),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_274),
.A2(n_227),
.B(n_229),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_269),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_349),
.Y(n_384)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_352),
.B1(n_353),
.B2(n_283),
.Y(n_375)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_343),
.Y(n_389)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_345),
.A2(n_292),
.B(n_275),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_261),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_296),
.B(n_252),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_350),
.B(n_351),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_315),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_272),
.A2(n_235),
.B1(n_252),
.B2(n_290),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_272),
.A2(n_235),
.B1(n_276),
.B2(n_325),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_298),
.B(n_288),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_354),
.B(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_299),
.A2(n_304),
.B1(n_286),
.B2(n_306),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_313),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_281),
.B(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_361),
.B(n_365),
.Y(n_400)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_303),
.B(n_281),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_273),
.A2(n_294),
.B(n_280),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_366),
.A2(n_275),
.B(n_321),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_275),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_367),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_281),
.B(n_276),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_276),
.B(n_285),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_371),
.Y(n_374)
);

OA22x2_ASAP7_75t_L g373 ( 
.A1(n_353),
.A2(n_284),
.B1(n_283),
.B2(n_273),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_358),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_375),
.A2(n_385),
.B1(n_391),
.B2(n_402),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_377),
.A2(n_403),
.B1(n_345),
.B2(n_366),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_349),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_396),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_334),
.A2(n_352),
.B1(n_289),
.B2(n_347),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_388),
.B(n_319),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_334),
.A2(n_293),
.B1(n_314),
.B2(n_309),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_343),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_397),
.A2(n_398),
.B(n_348),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_347),
.A2(n_328),
.B1(n_320),
.B2(n_321),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_341),
.A2(n_309),
.B1(n_282),
.B2(n_316),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_297),
.B1(n_316),
.B2(n_300),
.Y(n_403)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_405),
.Y(n_409)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_410),
.A2(n_411),
.B1(n_429),
.B2(n_430),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_371),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_424),
.C(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_381),
.B(n_360),
.Y(n_414)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_376),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_421),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_404),
.B(n_400),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_417),
.B(n_425),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_330),
.Y(n_420)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_420),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_405),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_341),
.B1(n_336),
.B2(n_332),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_422),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_364),
.B1(n_368),
.B2(n_344),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_364),
.C(n_329),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_339),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_426),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_405),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_427),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_383),
.B(n_361),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_428),
.Y(n_439)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_377),
.A2(n_364),
.B1(n_340),
.B2(n_369),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_436),
.B1(n_373),
.B2(n_387),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_342),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_432),
.A2(n_433),
.B(n_435),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_384),
.B(n_356),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_402),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_357),
.B1(n_355),
.B2(n_370),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_384),
.B(n_337),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_437),
.B(n_393),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_446),
.C(n_449),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_399),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_448),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_445),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_392),
.C(n_374),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_427),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_374),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_388),
.C(n_389),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_398),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_451),
.C(n_453),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_389),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_373),
.C(n_393),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_410),
.B(n_387),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_426),
.C(n_373),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_464),
.A2(n_419),
.B1(n_437),
.B2(n_418),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_433),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_470),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_417),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_466),
.B(n_475),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_411),
.B1(n_416),
.B2(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_458),
.A2(n_413),
.B1(n_415),
.B2(n_408),
.Y(n_468)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_434),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_409),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_477),
.Y(n_492)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_463),
.Y(n_473)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_473),
.Y(n_504)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_476),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_452),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_448),
.B(n_435),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_409),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_479),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_439),
.B1(n_453),
.B2(n_456),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_441),
.A2(n_421),
.B(n_418),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_481),
.A2(n_441),
.B(n_461),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_419),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_484),
.C(n_485),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_420),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_425),
.C(n_395),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_460),
.C(n_447),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_487),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_489),
.A2(n_395),
.B(n_394),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_491),
.A2(n_470),
.B1(n_472),
.B2(n_430),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_493),
.B(n_496),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_469),
.A2(n_460),
.B(n_455),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_464),
.C(n_455),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_502),
.C(n_482),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_484),
.A2(n_459),
.B1(n_444),
.B2(n_457),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_482),
.B1(n_472),
.B2(n_477),
.Y(n_509)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_485),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_469),
.B(n_406),
.C(n_462),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_429),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_505),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_511),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_509),
.B(n_490),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_432),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_510),
.B(n_512),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_471),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_498),
.B(n_497),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_491),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_483),
.B(n_465),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_517),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_505),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_506),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_406),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_519),
.B(n_521),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_489),
.B(n_503),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_494),
.A2(n_394),
.B1(n_401),
.B2(n_407),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_527),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_526),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_492),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_512),
.B(n_508),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_516),
.B(n_504),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_529),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_500),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_515),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_511),
.C(n_488),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_535),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_518),
.B1(n_520),
.B2(n_507),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_507),
.Y(n_536)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_536),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_499),
.C(n_493),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_541),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_539),
.B(n_543),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_531),
.A2(n_506),
.B1(n_509),
.B2(n_521),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_524),
.A2(n_505),
.B1(n_514),
.B2(n_495),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_540),
.B(n_526),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_538),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_495),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_550),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_525),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_546),
.A2(n_536),
.B(n_542),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_552),
.A2(n_553),
.B(n_554),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_544),
.A2(n_539),
.B1(n_538),
.B2(n_492),
.Y(n_554)
);

AOI321xp33_ASAP7_75t_L g556 ( 
.A1(n_551),
.A2(n_547),
.A3(n_549),
.B1(n_407),
.B2(n_401),
.C(n_372),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_549),
.C(n_362),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_557),
.A2(n_555),
.B(n_372),
.Y(n_558)
);

OAI33xp33_ASAP7_75t_L g559 ( 
.A1(n_558),
.A2(n_295),
.A3(n_319),
.B1(n_326),
.B2(n_363),
.B3(n_528),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_295),
.Y(n_560)
);


endmodule