module real_jpeg_7109_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_5;
wire n_36;
wire n_39;
wire n_40;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g4 ( 
.A(n_5),
.Y(n_4)
);

AOI211xp5_ASAP7_75t_L g5 ( 
.A1(n_6),
.A2(n_19),
.B(n_34),
.C(n_35),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_6),
.B(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

OA22x2_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_12),
.B1(n_14),
.B2(n_18),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_9),
.B(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);


endmodule