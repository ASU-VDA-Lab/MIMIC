module real_aes_8990_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g260 ( .A1(n_0), .A2(n_261), .B(n_262), .C(n_266), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_1), .B(n_255), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_2), .B(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_3), .A2(n_249), .B(n_334), .Y(n_333) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_4), .A2(n_222), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g213 ( .A(n_5), .Y(n_213) );
AND2x6_ASAP7_75t_L g247 ( .A(n_5), .B(n_211), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_5), .B(n_532), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_6), .A2(n_230), .B(n_247), .C(n_312), .Y(n_311) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_7), .A2(n_21), .B1(n_90), .B2(n_95), .Y(n_98) );
INVx1_ASAP7_75t_L g227 ( .A(n_8), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_9), .B(n_241), .Y(n_348) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_10), .A2(n_23), .B1(n_90), .B2(n_91), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_11), .A2(n_230), .B(n_275), .C(n_282), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_12), .A2(n_53), .B1(n_109), .B2(n_114), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_13), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_14), .A2(n_230), .B(n_282), .C(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_15), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_16), .A2(n_81), .B1(n_185), .B2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_16), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_17), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_18), .A2(n_249), .B(n_257), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_19), .Y(n_143) );
INVx2_ASAP7_75t_L g232 ( .A(n_20), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_22), .A2(n_245), .B(n_298), .C(n_299), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g204 ( .A1(n_23), .A2(n_38), .B1(n_49), .B2(n_205), .C(n_206), .Y(n_204) );
INVxp67_ASAP7_75t_L g207 ( .A(n_23), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_24), .B(n_347), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_25), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_26), .B(n_273), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_27), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_28), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_29), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_30), .B(n_241), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_31), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_32), .B(n_249), .Y(n_343) );
AOI22xp5_ASAP7_75t_SL g527 ( .A1(n_32), .A2(n_81), .B1(n_185), .B2(n_528), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_32), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_33), .A2(n_245), .B(n_298), .C(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g263 ( .A(n_34), .Y(n_263) );
INVx1_ASAP7_75t_L g326 ( .A(n_35), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_36), .B(n_249), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_37), .Y(n_287) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_38), .A2(n_59), .B1(n_90), .B2(n_91), .Y(n_89) );
INVxp67_ASAP7_75t_L g208 ( .A(n_38), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_39), .Y(n_131) );
INVx1_ASAP7_75t_L g211 ( .A(n_40), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_41), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_42), .B(n_255), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_43), .A2(n_237), .B(n_281), .C(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g226 ( .A(n_44), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_45), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_46), .B(n_241), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_47), .A2(n_56), .B1(n_133), .B2(n_137), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_48), .B(n_242), .Y(n_313) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_49), .A2(n_66), .B1(n_90), .B2(n_95), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_50), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_51), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_52), .B(n_277), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_54), .A2(n_230), .B(n_235), .C(n_245), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_55), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_57), .B(n_279), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_58), .Y(n_304) );
INVx2_ASAP7_75t_L g224 ( .A(n_60), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_61), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_62), .B(n_265), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_63), .A2(n_192), .B1(n_198), .B2(n_199), .Y(n_191) );
INVx1_ASAP7_75t_L g198 ( .A(n_63), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_64), .A2(n_72), .B1(n_189), .B2(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_64), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_65), .A2(n_75), .B1(n_196), .B2(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_65), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_65), .B(n_249), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_67), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_68), .Y(n_101) );
INVxp67_ASAP7_75t_L g338 ( .A(n_69), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_70), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_70), .Y(n_193) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
INVx1_ASAP7_75t_L g189 ( .A(n_72), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_73), .A2(n_81), .B1(n_184), .B2(n_185), .Y(n_80) );
INVx2_ASAP7_75t_L g184 ( .A(n_73), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_74), .Y(n_148) );
INVx1_ASAP7_75t_L g197 ( .A(n_75), .Y(n_197) );
INVx1_ASAP7_75t_L g236 ( .A(n_76), .Y(n_236) );
AND2x2_ASAP7_75t_L g328 ( .A(n_77), .B(n_285), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_201), .B1(n_214), .B2(n_523), .C(n_526), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_186), .Y(n_79) );
INVx1_ASAP7_75t_L g185 ( .A(n_81), .Y(n_185) );
AND2x2_ASAP7_75t_SL g81 ( .A(n_82), .B(n_141), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_119), .Y(n_82) );
OAI221xp5_ASAP7_75t_SL g83 ( .A1(n_84), .A2(n_101), .B1(n_102), .B2(n_107), .C(n_108), .Y(n_83) );
INVx3_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_96), .Y(n_86) );
AND2x6_ASAP7_75t_L g111 ( .A(n_87), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g162 ( .A(n_87), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_94), .Y(n_106) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_89), .B(n_94), .Y(n_118) );
AND2x2_ASAP7_75t_L g129 ( .A(n_89), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g158 ( .A(n_89), .B(n_98), .Y(n_158) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g95 ( .A(n_92), .Y(n_95) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
INVx1_ASAP7_75t_L g157 ( .A(n_94), .Y(n_157) );
AND2x4_ASAP7_75t_L g105 ( .A(n_96), .B(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g116 ( .A(n_96), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_96), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_99), .Y(n_96) );
OR2x2_ASAP7_75t_L g113 ( .A(n_97), .B(n_100), .Y(n_113) );
AND2x2_ASAP7_75t_L g124 ( .A(n_97), .B(n_100), .Y(n_124) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g163 ( .A(n_98), .B(n_100), .Y(n_163) );
AND2x2_ASAP7_75t_L g156 ( .A(n_99), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g176 ( .A(n_99), .Y(n_176) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g147 ( .A(n_106), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g151 ( .A(n_106), .B(n_124), .Y(n_151) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx11_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g146 ( .A(n_113), .B(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_L g139 ( .A(n_118), .B(n_140), .Y(n_139) );
OAI221xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_125), .B1(n_126), .B2(n_131), .C(n_132), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx6_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g136 ( .A(n_124), .B(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx8_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx6_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_152), .C(n_171), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B1(n_148), .B2(n_149), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI222xp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .B1(n_160), .B2(n_164), .C1(n_165), .C2(n_170), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx4f_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g169 ( .A(n_157), .Y(n_169) );
AND2x4_ASAP7_75t_L g168 ( .A(n_158), .B(n_169), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_158), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx4f_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_177), .B2(n_178), .Y(n_171) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_191), .B2(n_200), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_191), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_192), .Y(n_199) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_197), .A2(n_310), .B(n_311), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
AND3x1_ASAP7_75t_SL g203 ( .A(n_204), .B(n_209), .C(n_212), .Y(n_203) );
INVxp67_ASAP7_75t_L g532 ( .A(n_204), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_SL g534 ( .A(n_209), .Y(n_534) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_209), .A2(n_250), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g542 ( .A(n_209), .Y(n_542) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_210), .B(n_213), .Y(n_536) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_SL g541 ( .A(n_212), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR3x1_ASAP7_75t_L g215 ( .A(n_216), .B(n_431), .C(n_480), .Y(n_215) );
NAND5xp2_ASAP7_75t_L g216 ( .A(n_217), .B(n_365), .C(n_394), .D(n_402), .E(n_417), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_289), .B(n_305), .C(n_349), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_269), .Y(n_218) );
AND2x2_ASAP7_75t_L g360 ( .A(n_219), .B(n_357), .Y(n_360) );
AND2x2_ASAP7_75t_L g393 ( .A(n_219), .B(n_270), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_219), .B(n_293), .Y(n_486) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_254), .Y(n_219) );
INVx2_ASAP7_75t_L g292 ( .A(n_220), .Y(n_292) );
BUFx2_ASAP7_75t_L g460 ( .A(n_220), .Y(n_460) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_228), .B(n_252), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_221), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g255 ( .A(n_221), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_221), .B(n_304), .Y(n_303) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_221), .A2(n_309), .B(n_318), .Y(n_308) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_222), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_222), .A2(n_343), .B(n_344), .Y(n_342) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g320 ( .A(n_223), .Y(n_320) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_224), .B(n_225), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_248), .Y(n_228) );
INVx5_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
AND2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
BUFx3_ASAP7_75t_L g267 ( .A(n_231), .Y(n_267) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g251 ( .A(n_232), .Y(n_251) );
INVx1_ASAP7_75t_L g317 ( .A(n_232), .Y(n_317) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_234), .Y(n_239) );
INVx3_ASAP7_75t_L g242 ( .A(n_234), .Y(n_242) );
AND2x2_ASAP7_75t_L g250 ( .A(n_234), .B(n_251), .Y(n_250) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
INVx1_ASAP7_75t_L g347 ( .A(n_234), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_240), .C(n_243), .Y(n_235) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g277 ( .A(n_239), .Y(n_277) );
INVx2_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_241), .B(n_338), .Y(n_337) );
INVx5_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_246), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_246), .A2(n_259), .B(n_335), .C(n_336), .Y(n_334) );
INVx4_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g249 ( .A(n_247), .B(n_250), .Y(n_249) );
BUFx3_ASAP7_75t_L g282 ( .A(n_247), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_247), .B(n_250), .Y(n_310) );
BUFx2_ASAP7_75t_L g273 ( .A(n_249), .Y(n_273) );
INVx1_ASAP7_75t_L g281 ( .A(n_251), .Y(n_281) );
AND2x2_ASAP7_75t_L g269 ( .A(n_254), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g358 ( .A(n_254), .Y(n_358) );
AND2x2_ASAP7_75t_L g444 ( .A(n_254), .B(n_357), .Y(n_444) );
AND2x2_ASAP7_75t_L g499 ( .A(n_254), .B(n_292), .Y(n_499) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_268), .Y(n_254) );
INVx2_ASAP7_75t_L g298 ( .A(n_259), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx4_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
INVx1_ASAP7_75t_L g416 ( .A(n_269), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_269), .B(n_293), .Y(n_463) );
INVx5_ASAP7_75t_L g357 ( .A(n_270), .Y(n_357) );
AND2x4_ASAP7_75t_L g378 ( .A(n_270), .B(n_358), .Y(n_378) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_270), .Y(n_400) );
AND2x2_ASAP7_75t_L g475 ( .A(n_270), .B(n_460), .Y(n_475) );
AND2x2_ASAP7_75t_L g478 ( .A(n_270), .B(n_294), .Y(n_478) );
OR2x6_ASAP7_75t_L g270 ( .A(n_271), .B(n_286), .Y(n_270) );
AOI21xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_274), .B(n_283), .Y(n_271) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_273), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .B(n_280), .Y(n_275) );
INVx2_ASAP7_75t_L g279 ( .A(n_277), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_279), .A2(n_300), .B(n_301), .C(n_302), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_279), .A2(n_302), .B(n_326), .C(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g288 ( .A(n_285), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_285), .A2(n_296), .B(n_297), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_323), .B(n_324), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_289), .B(n_358), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_289), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g383 ( .A(n_291), .B(n_358), .Y(n_383) );
AND2x2_ASAP7_75t_L g401 ( .A(n_291), .B(n_294), .Y(n_401) );
INVx1_ASAP7_75t_L g421 ( .A(n_291), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_291), .B(n_357), .Y(n_466) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_291), .Y(n_508) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_292), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_293), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_293), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_293), .A2(n_353), .B(n_414), .C(n_416), .Y(n_413) );
AND2x2_ASAP7_75t_L g420 ( .A(n_293), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g429 ( .A(n_293), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g433 ( .A(n_293), .B(n_357), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_293), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g448 ( .A(n_293), .B(n_358), .Y(n_448) );
AND2x2_ASAP7_75t_L g498 ( .A(n_293), .B(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g362 ( .A(n_294), .Y(n_362) );
AND2x2_ASAP7_75t_L g403 ( .A(n_294), .B(n_356), .Y(n_403) );
AND2x2_ASAP7_75t_L g415 ( .A(n_294), .B(n_390), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_294), .B(n_444), .Y(n_462) );
OR2x6_ASAP7_75t_L g294 ( .A(n_295), .B(n_303), .Y(n_294) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_329), .Y(n_305) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_321), .Y(n_306) );
OR2x2_ASAP7_75t_L g353 ( .A(n_307), .B(n_321), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_307), .B(n_360), .C(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_307), .B(n_331), .Y(n_370) );
OR2x2_ASAP7_75t_L g385 ( .A(n_307), .B(n_373), .Y(n_385) );
AND2x2_ASAP7_75t_L g391 ( .A(n_307), .B(n_340), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_307), .B(n_522), .Y(n_521) );
INVx5_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_308), .B(n_331), .Y(n_388) );
AND2x2_ASAP7_75t_L g427 ( .A(n_308), .B(n_341), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_308), .B(n_340), .Y(n_455) );
OR2x2_ASAP7_75t_L g458 ( .A(n_308), .B(n_340), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_315), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_315), .A2(n_346), .B(n_348), .Y(n_345) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx5_ASAP7_75t_SL g373 ( .A(n_321), .Y(n_373) );
OR2x2_ASAP7_75t_L g379 ( .A(n_321), .B(n_330), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_321), .B(n_396), .Y(n_395) );
AOI321xp33_ASAP7_75t_L g402 ( .A1(n_321), .A2(n_403), .A3(n_404), .B1(n_405), .B2(n_411), .C(n_413), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_321), .B(n_329), .Y(n_412) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_321), .Y(n_425) );
OR2x2_ASAP7_75t_L g472 ( .A(n_321), .B(n_370), .Y(n_472) );
AND2x2_ASAP7_75t_L g494 ( .A(n_321), .B(n_391), .Y(n_494) );
AND2x2_ASAP7_75t_L g513 ( .A(n_321), .B(n_331), .Y(n_513) );
OR2x6_ASAP7_75t_L g321 ( .A(n_322), .B(n_328), .Y(n_321) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_340), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_331), .B(n_340), .Y(n_354) );
AND2x2_ASAP7_75t_L g363 ( .A(n_331), .B(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
AND2x2_ASAP7_75t_L g396 ( .A(n_331), .B(n_391), .Y(n_396) );
INVxp67_ASAP7_75t_L g426 ( .A(n_331), .Y(n_426) );
OR2x2_ASAP7_75t_L g468 ( .A(n_331), .B(n_373), .Y(n_468) );
OA21x2_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_339), .Y(n_331) );
OR2x2_ASAP7_75t_L g350 ( .A(n_340), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g364 ( .A(n_340), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_340), .B(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g446 ( .A(n_340), .B(n_390), .Y(n_446) );
AND2x2_ASAP7_75t_L g484 ( .A(n_340), .B(n_373), .Y(n_484) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_341), .B(n_373), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B(n_355), .C(n_359), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_350), .A2(n_352), .B1(n_477), .B2(n_479), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_352), .A2(n_375), .B1(n_430), .B2(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_SL g504 ( .A(n_353), .Y(n_504) );
INVx1_ASAP7_75t_SL g404 ( .A(n_354), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_356), .B(n_376), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g417 ( .A1(n_356), .A2(n_397), .B1(n_404), .B2(n_418), .C1(n_422), .C2(n_428), .Y(n_417) );
AND2x2_ASAP7_75t_L g507 ( .A(n_356), .B(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_357), .B(n_377), .Y(n_452) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_357), .Y(n_489) );
AND2x2_ASAP7_75t_L g492 ( .A(n_357), .B(n_401), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_357), .B(n_508), .Y(n_518) );
INVx1_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_358), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_360), .A2(n_501), .B(n_502), .C(n_505), .Y(n_500) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_362), .B(n_424), .C(n_427), .Y(n_423) );
OR2x2_ASAP7_75t_L g451 ( .A(n_362), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_362), .B(n_378), .Y(n_479) );
OR2x2_ASAP7_75t_L g384 ( .A(n_364), .B(n_385), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B(n_374), .C(n_386), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_367), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g473 ( .A(n_368), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_369), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g387 ( .A(n_372), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_373), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g441 ( .A(n_373), .B(n_391), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_373), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_373), .B(n_390), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_379), .B1(n_380), .B2(n_384), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_376), .B(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_378), .B(n_420), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g442 ( .A1(n_379), .A2(n_443), .B1(n_445), .B2(n_447), .C(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g497 ( .A(n_382), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g510 ( .A(n_382), .B(n_499), .Y(n_510) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx1_ASAP7_75t_L g501 ( .A(n_384), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_385), .A2(n_468), .B(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_392), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g434 ( .A(n_395), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_396), .A2(n_482), .B1(n_485), .B2(n_487), .C(n_490), .Y(n_481) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_404), .A2(n_494), .B1(n_495), .B2(n_497), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g470 ( .A(n_406), .Y(n_470) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp67_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g474 ( .A(n_410), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g439 ( .A(n_415), .Y(n_439) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_420), .B(n_444), .Y(n_496) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_426), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g512 ( .A(n_427), .B(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g519 ( .A(n_427), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_434), .B(n_435), .C(n_469), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B(n_442), .C(n_461), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g522 ( .A(n_446), .Y(n_522) );
AND2x2_ASAP7_75t_L g459 ( .A(n_448), .B(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B1(n_457), .B2(n_459), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OR2x2_ASAP7_75t_L g467 ( .A(n_455), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g520 ( .A(n_456), .Y(n_520) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI31xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .A3(n_464), .B(n_467), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_473), .C(n_476), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
NAND5xp2_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .C(n_500), .D(n_514), .E(n_517), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_492), .A2(n_518), .B1(n_519), .B2(n_521), .Y(n_517) );
INVx1_ASAP7_75t_SL g516 ( .A(n_494), .Y(n_516) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B(n_511), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
OAI322xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .A3(n_529), .B1(n_533), .B2(n_535), .C1(n_537), .C2(n_539), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
endmodule