module fake_jpeg_17589_n_23 (n_3, n_2, n_1, n_0, n_4, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_8),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_8),
.C(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_7),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_14),
.B(n_11),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_17),
.B(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_8),
.B(n_3),
.Y(n_19)
);

AOI322xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_20),
.A3(n_5),
.B1(n_18),
.B2(n_9),
.C1(n_2),
.C2(n_4),
.Y(n_21)
);

OAI31xp33_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_5),
.A3(n_9),
.B(n_4),
.Y(n_22)
);

AOI221xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_2),
.B1(n_3),
.B2(n_9),
.C(n_19),
.Y(n_23)
);


endmodule