module fake_jpeg_7843_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2x1_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_29),
.B1(n_16),
.B2(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_51),
.B1(n_22),
.B2(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_32),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_34),
.B1(n_20),
.B2(n_23),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_16),
.B1(n_31),
.B2(n_27),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_59),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_40),
.B1(n_28),
.B2(n_19),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_69),
.B1(n_80),
.B2(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_36),
.B1(n_39),
.B2(n_33),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_68),
.B1(n_81),
.B2(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_70),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_39),
.B1(n_33),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_19),
.B1(n_28),
.B2(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_26),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_79),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_41),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_88),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_56),
.B1(n_55),
.B2(n_52),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_130)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_30),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_43),
.B(n_35),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_109),
.B(n_20),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_43),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_83),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_22),
.B1(n_17),
.B2(n_26),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_41),
.B(n_35),
.C(n_20),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_78),
.B1(n_65),
.B2(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_35),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_70),
.C(n_64),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_116),
.C(n_127),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_82),
.C(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_123),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_67),
.B1(n_62),
.B2(n_71),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_126),
.B1(n_94),
.B2(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_133),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_64),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_30),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_30),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_17),
.B1(n_78),
.B2(n_23),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_106),
.B1(n_108),
.B2(n_23),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_91),
.B1(n_104),
.B2(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_141),
.B(n_148),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_85),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_147),
.C(n_111),
.Y(n_164)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_99),
.CON(n_143),
.SN(n_143)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_149),
.B(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_109),
.C(n_94),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_108),
.B(n_99),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_110),
.B1(n_130),
.B2(n_115),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_98),
.A3(n_30),
.B1(n_15),
.B2(n_14),
.C1(n_13),
.C2(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_13),
.C(n_3),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_143),
.A3(n_137),
.B1(n_154),
.B2(n_138),
.C(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_174),
.C(n_4),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_111),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_175),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_1),
.C(n_3),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_3),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_165),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_150),
.B(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_158),
.B(n_167),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_135),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_186),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_185),
.B1(n_171),
.B2(n_159),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_142),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.C(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_4),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_190),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_4),
.C(n_5),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_192),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_199),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_173),
.C(n_167),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_183),
.B1(n_179),
.B2(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_206),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_171),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_157),
.B(n_200),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_177),
.B1(n_176),
.B2(n_182),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_208),
.B1(n_203),
.B2(n_205),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_5),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_7),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_200),
.B1(n_195),
.B2(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_217),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_213),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_6),
.B(n_7),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_215),
.B(n_9),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_6),
.B(n_7),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_8),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_219),
.C(n_9),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_10),
.B(n_227),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_10),
.Y(n_230)
);


endmodule