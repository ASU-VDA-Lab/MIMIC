module fake_jpeg_21548_n_314 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_25),
.B1(n_21),
.B2(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_25),
.B1(n_21),
.B2(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_25),
.B1(n_32),
.B2(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_42),
.B1(n_34),
.B2(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_67),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_42),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_38),
.C(n_37),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_70),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_19),
.B(n_18),
.C(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_77),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_81),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_16),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_89),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVxp33_ASAP7_75t_SL g90 ( 
.A(n_46),
.Y(n_90)
);

AND2x4_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_38),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_92),
.Y(n_129)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_122),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_121),
.B(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_38),
.C(n_37),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_122),
.C(n_33),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_62),
.A2(n_36),
.B1(n_20),
.B2(n_28),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_82),
.B1(n_23),
.B2(n_84),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_38),
.C(n_37),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_38),
.B(n_23),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_143),
.Y(n_166)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_24),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_150),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_19),
.B1(n_18),
.B2(n_28),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_92),
.B1(n_99),
.B2(n_66),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_146),
.B1(n_115),
.B2(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_15),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_101),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_149),
.A2(n_152),
.B(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_61),
.B(n_14),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_157),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_88),
.B(n_73),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_68),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_33),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_110),
.B(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_74),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_172),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_104),
.B1(n_132),
.B2(n_113),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_33),
.B(n_157),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_187),
.B(n_24),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_114),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_182),
.B1(n_183),
.B2(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_104),
.B1(n_118),
.B2(n_110),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_127),
.B1(n_20),
.B2(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_89),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_181),
.C(n_188),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_112),
.C(n_110),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_141),
.B1(n_146),
.B2(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_128),
.B1(n_130),
.B2(n_103),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_109),
.B(n_125),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_109),
.C(n_125),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_138),
.A2(n_128),
.B1(n_103),
.B2(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_197),
.B(n_202),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_13),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_200),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_91),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_190),
.B1(n_193),
.B2(n_162),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_0),
.B(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_127),
.B1(n_20),
.B2(n_27),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_215),
.B1(n_174),
.B2(n_184),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_217),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_218),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_79),
.B(n_65),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_31),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_31),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_185),
.C(n_176),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_219),
.C(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_166),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_189),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_14),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_216),
.A2(n_174),
.B1(n_178),
.B2(n_184),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_29),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_29),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_14),
.B(n_29),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_178),
.B(n_167),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_225),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_231),
.B(n_236),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_169),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_6),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_205),
.B(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_228),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_253),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_204),
.B1(n_201),
.B2(n_192),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_248),
.B1(n_260),
.B2(n_208),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_199),
.B1(n_215),
.B2(n_220),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_213),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_195),
.C(n_218),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_242),
.C(n_221),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_219),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_207),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_199),
.B1(n_196),
.B2(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_251),
.C(n_257),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_211),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_274),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_234),
.B1(n_239),
.B2(n_222),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_212),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_275),
.B(n_259),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_240),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_240),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_248),
.B1(n_260),
.B2(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_262),
.C(n_274),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_287),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_222),
.C(n_252),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_255),
.B1(n_202),
.B2(n_197),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_278),
.B1(n_286),
.B2(n_290),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_208),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_6),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_276),
.B(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_282),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_27),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_302),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_287),
.B1(n_279),
.B2(n_283),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_291),
.B(n_7),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_10),
.B(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_27),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.C(n_27),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.C(n_305),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_297),
.B(n_11),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_31),
.C(n_6),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_0),
.Y(n_314)
);


endmodule