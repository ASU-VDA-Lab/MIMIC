module real_jpeg_33049_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_1),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_1),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_1),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_1),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_1),
.B(n_412),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_1),
.Y(n_435)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_202),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_2),
.B(n_428),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_2),
.B(n_459),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_3),
.B(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_4),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_4),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_4),
.B(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_6),
.Y(n_103)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_7),
.B(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_7),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_7),
.B(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_9),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_9),
.B(n_35),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_9),
.B(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_10),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_10),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_10),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_10),
.B(n_152),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_10),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_10),
.B(n_470),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_13),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_14),
.A2(n_29),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_14),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_14),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_14),
.B(n_312),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_14),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_14),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_14),
.B(n_475),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_15),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_16),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_17),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_149),
.Y(n_148)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_17),
.B(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_21),
.B(n_519),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_189),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_187),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_156),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_24),
.B(n_156),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_68),
.C(n_126),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_25),
.B(n_68),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_56),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_27),
.B(n_42),
.C(n_56),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_34),
.C(n_37),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_28),
.A2(n_34),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_32),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_33),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_34),
.A2(n_89),
.B1(n_292),
.B2(n_296),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XOR2x2_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_41),
.Y(n_167)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_41),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_41),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.C(n_53),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_44),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_43),
.B(n_58),
.C(n_64),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_43),
.A2(n_44),
.B1(n_212),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_44),
.B(n_212),
.C(n_215),
.Y(n_211)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_47),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_76),
.C(n_81),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_53),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_53),
.B(n_227),
.Y(n_262)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_55),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_55),
.Y(n_410)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_55),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_57),
.A2(n_58),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_57),
.A2(n_58),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_57),
.B(n_198),
.C(n_201),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_60),
.Y(n_340)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2x1_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_91),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_69),
.B(n_108),
.C(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.C(n_87),
.Y(n_69)
);

XOR2x2_ASAP7_75t_L g375 ( 
.A(n_70),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_73),
.A2(n_227),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_73),
.B(n_227),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_L g446 ( 
.A1(n_73),
.A2(n_227),
.B(n_415),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_74),
.A2(n_75),
.B1(n_87),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_83),
.Y(n_143)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_80),
.Y(n_319)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_82),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_85),
.Y(n_272)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_89),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_108),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_95),
.B(n_96),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_95),
.B(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_110),
.C(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_101),
.B(n_104),
.C(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_101),
.B(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_103),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_134),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_107),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.C(n_124),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_115),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_112),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_110),
.B(n_130),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_110),
.B(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_110),
.B(n_408),
.Y(n_442)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_111),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_115),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_115),
.B(n_275),
.C(n_280),
.Y(n_297)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_129),
.C(n_132),
.Y(n_128)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_124),
.A2(n_132),
.B1(n_133),
.B2(n_140),
.Y(n_362)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_127),
.B(n_515),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.C(n_141),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_128),
.A2(n_137),
.B1(n_138),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_128),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_129),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_130),
.B(n_205),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_131),
.Y(n_477)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_141),
.B(n_379),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_142),
.B(n_146),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_144),
.B(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_148),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_151),
.B(n_154),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_184),
.B2(n_185),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_176),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_182),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_512),
.B(n_517),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_392),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_355),
.B(n_388),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_322),
.B(n_354),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_298),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_194),
.B(n_298),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_250),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_195),
.B(n_251),
.C(n_282),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_221),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_196),
.B(n_222),
.C(n_231),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.C(n_210),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g320 ( 
.A(n_197),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_204),
.B(n_211),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_209),
.B(n_410),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_209),
.B(n_487),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_212),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_214),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_215),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_218),
.Y(n_424)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_220),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_224)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_226),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_227),
.B(n_230),
.C(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_229),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_249),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_236),
.Y(n_463)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_237),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_238),
.Y(n_490)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_241),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_242),
.B(n_331),
.C(n_332),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OA21x2_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_253),
.B(n_257),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_282),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_260),
.C(n_273),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_273),
.Y(n_300)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx4f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_260),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.C(n_268),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_261),
.A2(n_262),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_263),
.A2(n_264),
.B1(n_268),
.B2(n_269),
.Y(n_404)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_297),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_285),
.C(n_297),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_292),
.C(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_320),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_299),
.B(n_396),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_302),
.B(n_320),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.C(n_308),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_304),
.B(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.C(n_317),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_310),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_450)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_317),
.B(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_323),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_325),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_326),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_344),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_343),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_367),
.C(n_368),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_337),
.C(n_342),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_339),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_343),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_386),
.C(n_387),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_349),
.C(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_SL g392 ( 
.A(n_355),
.B(n_393),
.C(n_510),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_371),
.B1(n_381),
.B2(n_384),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_372),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_372),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_365),
.C(n_369),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_369),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_364),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_363),
.C(n_364),
.Y(n_373)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_SL g516 ( 
.A(n_373),
.B(n_375),
.C(n_378),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_385),
.Y(n_390)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B(n_391),
.Y(n_388)
);

AO21x2_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_416),
.B(n_509),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_395),
.B(n_397),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.C(n_405),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_398),
.A2(n_399),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_399),
.B(n_503),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_402),
.B(n_405),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_402),
.B(n_405),
.Y(n_508)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.C(n_414),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_445),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_414),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_501),
.B(n_505),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_452),
.B(n_500),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_443),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_443),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_432),
.C(n_442),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_497),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_426),
.C(n_431),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_423),
.B(n_482),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_430),
.B2(n_431),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_426),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AO22x1_ASAP7_75t_L g497 ( 
.A1(n_432),
.A2(n_433),
.B1(n_442),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_434),
.A2(n_437),
.B1(n_438),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_448),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_444),
.B(n_449),
.C(n_451),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_494),
.B(n_499),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_478),
.B(n_493),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_467),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_467),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_464),
.B2(n_465),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_461),
.C(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_473),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_468),
.A2(n_469),
.B1(n_473),
.B2(n_474),
.Y(n_491)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_SL g470 ( 
.A(n_471),
.Y(n_470)
);

INVx8_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_485),
.B(n_492),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_491),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_491),
.Y(n_492)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_496),
.Y(n_499)
);

NOR2x1p5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_514),
.B(n_516),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_518),
.Y(n_517)
);


endmodule