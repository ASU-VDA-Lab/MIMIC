module fake_jpeg_263_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_23),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_13),
.C(n_18),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_1),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_18),
.B(n_16),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_17),
.B(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_21),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_14),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_26),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_11),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_31),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_38),
.C(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_27),
.A3(n_33),
.B1(n_37),
.B2(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_44),
.B1(n_6),
.B2(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_5),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_53),
.A3(n_49),
.B1(n_54),
.B2(n_51),
.C1(n_50),
.C2(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.C(n_53),
.Y(n_61)
);


endmodule