module real_aes_316_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g101 ( .A1(n_0), .A2(n_56), .B1(n_91), .B2(n_102), .Y(n_101) );
AOI22xp33_ASAP7_75t_SL g79 ( .A1(n_1), .A2(n_80), .B1(n_81), .B2(n_158), .Y(n_79) );
INVx1_ASAP7_75t_L g158 ( .A(n_1), .Y(n_158) );
INVx1_ASAP7_75t_L g179 ( .A(n_2), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_3), .B(n_209), .Y(n_259) );
INVx1_ASAP7_75t_L g305 ( .A(n_4), .Y(n_305) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_5), .A2(n_18), .B1(n_91), .B2(n_99), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_6), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_7), .A2(n_34), .B1(n_153), .B2(n_156), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_8), .A2(n_47), .B1(n_149), .B2(n_150), .Y(n_148) );
INVx2_ASAP7_75t_L g208 ( .A(n_9), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g163 ( .A1(n_10), .A2(n_76), .B1(n_164), .B2(n_165), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_10), .Y(n_164) );
INVx1_ASAP7_75t_L g269 ( .A(n_11), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_12), .A2(n_50), .B1(n_114), .B2(n_119), .Y(n_113) );
INVx1_ASAP7_75t_L g266 ( .A(n_13), .Y(n_266) );
INVx1_ASAP7_75t_SL g252 ( .A(n_14), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_15), .B(n_219), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_15), .A2(n_80), .B1(n_81), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_15), .Y(n_543) );
AOI33xp33_ASAP7_75t_L g285 ( .A1(n_16), .A2(n_39), .A3(n_199), .B1(n_214), .B2(n_286), .B3(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g313 ( .A(n_17), .Y(n_313) );
OAI221xp5_ASAP7_75t_L g171 ( .A1(n_18), .A2(n_56), .B1(n_58), .B2(n_172), .C(n_174), .Y(n_171) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_19), .A2(n_69), .B(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g210 ( .A(n_19), .B(n_69), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_20), .B(n_240), .Y(n_249) );
INVx3_ASAP7_75t_L g91 ( .A(n_21), .Y(n_91) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_22), .A2(n_72), .B1(n_135), .B2(n_137), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_23), .A2(n_24), .B1(n_125), .B2(n_129), .Y(n_124) );
INVx1_ASAP7_75t_SL g92 ( .A(n_25), .Y(n_92) );
INVx1_ASAP7_75t_L g181 ( .A(n_26), .Y(n_181) );
AND2x2_ASAP7_75t_L g203 ( .A(n_26), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g228 ( .A(n_26), .B(n_179), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_27), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_28), .B(n_240), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_29), .A2(n_196), .B1(n_206), .B2(n_209), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_30), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_31), .B(n_219), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_32), .A2(n_161), .B1(n_162), .B2(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_32), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_33), .B(n_230), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_35), .B(n_219), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_36), .A2(n_68), .B1(n_104), .B2(n_109), .Y(n_103) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_37), .A2(n_58), .B1(n_91), .B2(n_95), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_38), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_40), .B(n_219), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_41), .A2(n_74), .B1(n_141), .B2(n_144), .Y(n_140) );
INVx1_ASAP7_75t_L g200 ( .A(n_42), .Y(n_200) );
INVx1_ASAP7_75t_L g221 ( .A(n_42), .Y(n_221) );
AND2x2_ASAP7_75t_L g298 ( .A(n_43), .B(n_246), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_44), .A2(n_60), .B1(n_212), .B2(n_240), .C(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_45), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_48), .B(n_206), .Y(n_321) );
AOI21xp5_ASAP7_75t_SL g235 ( .A1(n_49), .A2(n_212), .B(n_236), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_51), .A2(n_80), .B1(n_81), .B2(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_51), .Y(n_551) );
INVx1_ASAP7_75t_L g262 ( .A(n_52), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_53), .A2(n_160), .B1(n_166), .B2(n_167), .Y(n_159) );
INVx1_ASAP7_75t_L g166 ( .A(n_53), .Y(n_166) );
INVx1_ASAP7_75t_L g296 ( .A(n_54), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_55), .A2(n_212), .B(n_295), .Y(n_294) );
INVxp33_ASAP7_75t_L g176 ( .A(n_56), .Y(n_176) );
INVx1_ASAP7_75t_L g204 ( .A(n_57), .Y(n_204) );
INVx1_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVxp67_ASAP7_75t_L g175 ( .A(n_58), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_59), .B(n_240), .Y(n_288) );
AND2x2_ASAP7_75t_L g254 ( .A(n_61), .B(n_233), .Y(n_254) );
INVx1_ASAP7_75t_L g263 ( .A(n_62), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_63), .A2(n_212), .B(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_64), .A2(n_212), .B(n_217), .C(n_229), .Y(n_211) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_65), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_66), .B(n_85), .Y(n_84) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_67), .A2(n_212), .B1(n_283), .B2(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g237 ( .A(n_70), .Y(n_237) );
AND2x2_ASAP7_75t_L g289 ( .A(n_71), .B(n_233), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_73), .A2(n_311), .B(n_312), .C(n_314), .Y(n_310) );
BUFx2_ASAP7_75t_SL g173 ( .A(n_75), .Y(n_173) );
INVx1_ASAP7_75t_L g165 ( .A(n_76), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_76), .B(n_219), .Y(n_238) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_168), .B1(n_182), .B2(n_539), .C(n_541), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_159), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_133), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_103), .C(n_113), .D(n_124), .Y(n_83) );
INVx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx6_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_96), .Y(n_87) );
AND2x4_ASAP7_75t_L g111 ( .A(n_88), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g130 ( .A(n_88), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
AND2x2_ASAP7_75t_L g117 ( .A(n_89), .B(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
OAI22x1_ASAP7_75t_L g89 ( .A1(n_90), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx2_ASAP7_75t_L g99 ( .A(n_91), .Y(n_99) );
INVx1_ASAP7_75t_L g102 ( .A(n_91), .Y(n_102) );
AND2x2_ASAP7_75t_L g107 ( .A(n_94), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g118 ( .A(n_94), .Y(n_118) );
BUFx2_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
AND2x2_ASAP7_75t_L g143 ( .A(n_96), .B(n_107), .Y(n_143) );
AND2x4_ASAP7_75t_L g149 ( .A(n_96), .B(n_117), .Y(n_149) );
AND2x4_ASAP7_75t_L g155 ( .A(n_96), .B(n_147), .Y(n_155) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_100), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x4_ASAP7_75t_L g106 ( .A(n_98), .B(n_100), .Y(n_106) );
AND2x2_ASAP7_75t_L g122 ( .A(n_98), .B(n_101), .Y(n_122) );
INVx1_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
INVxp67_ASAP7_75t_L g112 ( .A(n_100), .Y(n_112) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g127 ( .A(n_101), .B(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g116 ( .A(n_106), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g157 ( .A(n_106), .B(n_147), .Y(n_157) );
AND2x2_ASAP7_75t_L g136 ( .A(n_107), .B(n_127), .Y(n_136) );
AND2x4_ASAP7_75t_L g147 ( .A(n_108), .B(n_118), .Y(n_147) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g126 ( .A(n_117), .B(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g138 ( .A(n_122), .B(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g151 ( .A(n_122), .B(n_147), .Y(n_151) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g146 ( .A(n_127), .B(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_128), .Y(n_132) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_140), .C(n_148), .D(n_152), .Y(n_133) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx8_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_160), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
AND3x1_ASAP7_75t_SL g170 ( .A(n_171), .B(n_177), .C(n_180), .Y(n_170) );
INVxp67_ASAP7_75t_L g549 ( .A(n_171), .Y(n_549) );
CKINVDCx8_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_177), .Y(n_547) );
AOI21xp33_ASAP7_75t_L g556 ( .A1(n_177), .A2(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g198 ( .A(n_178), .B(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_SL g554 ( .A(n_178), .B(n_180), .Y(n_554) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g216 ( .A(n_179), .B(n_200), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_180), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g213 ( .A(n_181), .B(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND4xp75_ASAP7_75t_L g187 ( .A(n_188), .B(n_390), .C(n_456), .D(n_519), .Y(n_187) );
NOR2x1_ASAP7_75t_L g188 ( .A(n_189), .B(n_353), .Y(n_188) );
OR3x1_ASAP7_75t_L g189 ( .A(n_190), .B(n_323), .C(n_350), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_255), .B(n_278), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_241), .Y(n_192) );
AND2x2_ASAP7_75t_L g453 ( .A(n_193), .B(n_423), .Y(n_453) );
INVx1_ASAP7_75t_L g526 ( .A(n_193), .Y(n_526) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_231), .Y(n_193) );
INVx2_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_194), .Y(n_341) );
AND2x2_ASAP7_75t_L g345 ( .A(n_194), .B(n_258), .Y(n_345) );
AND2x4_ASAP7_75t_L g361 ( .A(n_194), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_194), .Y(n_365) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_211), .Y(n_194) );
NOR3xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_201), .C(n_205), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x4_ASAP7_75t_L g240 ( .A(n_198), .B(n_202), .Y(n_240) );
OR2x6_ASAP7_75t_L g226 ( .A(n_199), .B(n_215), .Y(n_226) );
INVxp33_ASAP7_75t_L g286 ( .A(n_199), .Y(n_286) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_199), .Y(n_557) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g271 ( .A(n_200), .B(n_222), .Y(n_271) );
INVxp67_ASAP7_75t_L g558 ( .A(n_201), .Y(n_558) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g215 ( .A(n_204), .Y(n_215) );
AND2x6_ASAP7_75t_L g268 ( .A(n_204), .B(n_220), .Y(n_268) );
OAI222xp33_ASAP7_75t_L g541 ( .A1(n_205), .A2(n_542), .B1(n_544), .B2(n_550), .C1(n_552), .C2(n_555), .Y(n_541) );
INVx4_ASAP7_75t_L g233 ( .A(n_206), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_206), .B(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_207), .Y(n_230) );
AND2x4_ASAP7_75t_L g209 ( .A(n_208), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_208), .B(n_210), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_235), .B(n_239), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_209), .B(n_227), .Y(n_272) );
INVxp67_ASAP7_75t_L g320 ( .A(n_212), .Y(n_320) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_216), .Y(n_212) );
INVx1_ASAP7_75t_L g287 ( .A(n_214), .Y(n_287) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_227), .Y(n_217) );
INVx1_ASAP7_75t_L g264 ( .A(n_219), .Y(n_264) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_227), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_226), .A2(n_227), .B(n_252), .C(n_253), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_226), .A2(n_262), .B1(n_263), .B2(n_264), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_226), .A2(n_227), .B(n_296), .C(n_297), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_SL g304 ( .A1(n_226), .A2(n_227), .B(n_305), .C(n_306), .Y(n_304) );
INVxp67_ASAP7_75t_L g311 ( .A(n_226), .Y(n_311) );
INVx1_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_229), .A2(n_281), .B(n_289), .Y(n_280) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_229), .A2(n_281), .B(n_289), .Y(n_329) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_230), .A2(n_303), .B(n_307), .Y(n_302) );
AND2x2_ASAP7_75t_L g256 ( .A(n_231), .B(n_257), .Y(n_256) );
INVx4_ASAP7_75t_L g342 ( .A(n_231), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_231), .B(n_332), .Y(n_346) );
INVx2_ASAP7_75t_L g360 ( .A(n_231), .Y(n_360) );
AND2x4_ASAP7_75t_L g364 ( .A(n_231), .B(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_231), .Y(n_399) );
OR2x2_ASAP7_75t_L g405 ( .A(n_231), .B(n_244), .Y(n_405) );
NOR2x1_ASAP7_75t_SL g434 ( .A(n_231), .B(n_258), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_231), .B(n_508), .Y(n_536) );
OR2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx3_ASAP7_75t_L g291 ( .A(n_233), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_233), .A2(n_291), .B1(n_310), .B2(n_315), .Y(n_309) );
INVx1_ASAP7_75t_L g322 ( .A(n_240), .Y(n_322) );
AND2x2_ASAP7_75t_L g433 ( .A(n_241), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_242), .B(n_257), .Y(n_467) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g274 ( .A(n_244), .Y(n_274) );
INVx2_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
AND2x2_ASAP7_75t_L g356 ( .A(n_244), .B(n_258), .Y(n_356) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_244), .Y(n_383) );
INVx1_ASAP7_75t_L g424 ( .A(n_244), .Y(n_424) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .B(n_254), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_246), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_273), .Y(n_255) );
AND2x2_ASAP7_75t_L g436 ( .A(n_256), .B(n_331), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_257), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g503 ( .A(n_257), .Y(n_503) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g362 ( .A(n_258), .Y(n_362) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_265), .B(n_272), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_264), .B(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_269), .B2(n_270), .Y(n_265) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_273), .A2(n_440), .B(n_444), .C(n_450), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_275), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g486 ( .A(n_275), .Y(n_486) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g408 ( .A(n_277), .B(n_362), .Y(n_408) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_299), .Y(n_278) );
AOI32xp33_ASAP7_75t_L g444 ( .A1(n_279), .A2(n_428), .A3(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_290), .Y(n_279) );
INVx2_ASAP7_75t_L g370 ( .A(n_280), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_280), .B(n_302), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_288), .Y(n_281) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g382 ( .A(n_290), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_290), .B(n_308), .Y(n_413) );
AND2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_290), .Y(n_500) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_298), .Y(n_290) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_291), .A2(n_292), .B(n_298), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g401 ( .A(n_299), .B(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_326), .Y(n_352) );
AND2x2_ASAP7_75t_L g501 ( .A(n_300), .B(n_499), .Y(n_501) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_308), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
AND2x4_ASAP7_75t_L g377 ( .A(n_302), .B(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g411 ( .A(n_302), .Y(n_411) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_302), .Y(n_419) );
AND2x2_ASAP7_75t_L g428 ( .A(n_302), .B(n_308), .Y(n_428) );
INVx1_ASAP7_75t_L g512 ( .A(n_302), .Y(n_512) );
INVx2_ASAP7_75t_L g349 ( .A(n_308), .Y(n_349) );
INVx1_ASAP7_75t_L g376 ( .A(n_308), .Y(n_376) );
INVx1_ASAP7_75t_L g443 ( .A(n_308), .Y(n_443) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_316), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B1(n_321), .B2(n_322), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_322), .Y(n_540) );
OAI32xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_334), .A3(n_339), .B1(n_343), .B2(n_347), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_325), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_326), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g427 ( .A(n_326), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g452 ( .A(n_326), .Y(n_452) );
AND2x2_ASAP7_75t_L g533 ( .A(n_326), .B(n_375), .Y(n_533) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g348 ( .A(n_328), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g447 ( .A(n_328), .B(n_370), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_328), .B(n_349), .Y(n_469) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_328), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
INVx1_ASAP7_75t_L g402 ( .A(n_329), .Y(n_402) );
AND2x2_ASAP7_75t_L g417 ( .A(n_329), .B(n_349), .Y(n_417) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g445 ( .A(n_331), .B(n_434), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_331), .B(n_364), .Y(n_515) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_332), .Y(n_484) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_333), .Y(n_466) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g367 ( .A(n_336), .B(n_368), .Y(n_367) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_336), .B(n_452), .Y(n_451) );
NOR2xp67_ASAP7_75t_SL g538 ( .A(n_336), .B(n_476), .Y(n_538) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g395 ( .A(n_338), .B(n_349), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_339), .B(n_405), .Y(n_463) );
INVx2_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_340), .B(n_356), .Y(n_429) );
AND2x4_ASAP7_75t_SL g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_342), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g494 ( .A(n_342), .B(n_365), .Y(n_494) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_342), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_343), .B(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
OR2x2_ASAP7_75t_L g465 ( .A(n_344), .B(n_466), .Y(n_465) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_344), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g454 ( .A(n_345), .B(n_399), .Y(n_454) );
INVxp33_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_348), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g528 ( .A(n_348), .B(n_410), .Y(n_528) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_371), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_366), .Y(n_354) );
AND2x2_ASAP7_75t_L g489 ( .A(n_356), .B(n_364), .Y(n_489) );
NAND2xp33_ASAP7_75t_R g357 ( .A(n_358), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g531 ( .A(n_360), .Y(n_531) );
INVx4_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
INVx1_ASAP7_75t_L g508 ( .A(n_362), .Y(n_508) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g502 ( .A(n_364), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_SL g506 ( .A(n_364), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_367), .A2(n_432), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g396 ( .A(n_370), .B(n_382), .Y(n_396) );
AND2x2_ASAP7_75t_L g410 ( .A(n_370), .B(n_411), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_379), .B(n_384), .C(n_387), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g458 ( .A(n_374), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g386 ( .A(n_375), .Y(n_386) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g446 ( .A(n_376), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g455 ( .A(n_376), .B(n_377), .Y(n_455) );
INVx1_ASAP7_75t_L g487 ( .A(n_376), .Y(n_487) );
AND2x4_ASAP7_75t_L g468 ( .A(n_377), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g490 ( .A(n_377), .B(n_381), .Y(n_490) );
AND2x2_ASAP7_75t_L g498 ( .A(n_377), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g473 ( .A(n_381), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_381), .B(n_395), .Y(n_475) );
AND2x2_ASAP7_75t_L g478 ( .A(n_381), .B(n_428), .Y(n_478) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_382), .B(n_443), .Y(n_492) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_408), .Y(n_420) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g516 ( .A(n_386), .B(n_396), .Y(n_516) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_388), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g400 ( .A(n_389), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_389), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_430), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_414), .Y(n_391) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_397), .B1(n_401), .B2(n_403), .C1(n_406), .C2(n_409), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_399), .B(n_408), .Y(n_407) );
OR2x6_ASAP7_75t_L g479 ( .A(n_399), .B(n_449), .Y(n_479) );
NAND5xp2_ASAP7_75t_L g482 ( .A(n_399), .B(n_402), .C(n_418), .D(n_483), .E(n_485), .Y(n_482) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_400), .B(n_404), .Y(n_518) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_405), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_407), .A2(n_498), .B1(n_501), .B2(n_502), .Y(n_497) );
INVx2_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_408), .B(n_424), .Y(n_461) );
INVx3_ASAP7_75t_L g496 ( .A(n_409), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
AND2x2_ASAP7_75t_L g441 ( .A(n_410), .B(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
INVx2_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g437 ( .A(n_413), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_426), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_420), .B(n_421), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g425 ( .A(n_417), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_420), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_SL g507 ( .A(n_424), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_439), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g476 ( .A(n_447), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_450) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_480), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .C(n_470), .Y(n_457) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OA21x2_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B(n_468), .Y(n_462) );
NAND2xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_467), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_477), .B(n_479), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B(n_475), .C(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_474), .A2(n_514), .B1(n_516), .B2(n_517), .Y(n_513) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_504), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_488), .C(n_495), .D(n_497), .Y(n_481) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g493 ( .A(n_484), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g524 ( .A(n_487), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_491), .B2(n_493), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_493), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI21xp5_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_509), .B(n_513), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVxp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_534), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_524), .B(n_525), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_529), .B2(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
endmodule