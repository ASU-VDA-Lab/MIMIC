module fake_jpeg_28627_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_54),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_22),
.B(n_10),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_101),
.Y(n_106)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_10),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_66),
.B(n_88),
.Y(n_156)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_10),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_37),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_24),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_46),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_108),
.B(n_131),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_51),
.B1(n_50),
.B2(n_38),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_111),
.A2(n_130),
.B1(n_141),
.B2(n_147),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_138),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_51),
.B1(n_50),
.B2(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_24),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_61),
.A2(n_39),
.B1(n_37),
.B2(n_45),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_136),
.A2(n_155),
.B1(n_103),
.B2(n_79),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_88),
.B(n_42),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_55),
.A2(n_50),
.B1(n_41),
.B2(n_45),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_26),
.C(n_43),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_25),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_60),
.A2(n_50),
.B1(n_41),
.B2(n_45),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_162),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_45),
.B1(n_41),
.B2(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_59),
.B(n_35),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_96),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_70),
.B(n_35),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_47),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_42),
.B1(n_46),
.B2(n_43),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_106),
.A2(n_92),
.B1(n_91),
.B2(n_82),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_188),
.B1(n_202),
.B2(n_214),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_42),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_171),
.B(n_172),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_46),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_180),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_118),
.A2(n_63),
.B(n_43),
.C(n_36),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_199),
.Y(n_266)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_179),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_178),
.B(n_181),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_124),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_36),
.B1(n_26),
.B2(n_30),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_112),
.B(n_117),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_189),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_185),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_186),
.Y(n_262)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_34),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_105),
.A2(n_37),
.B1(n_39),
.B2(n_25),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_190),
.A2(n_142),
.B1(n_146),
.B2(n_127),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_33),
.B1(n_26),
.B2(n_30),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_119),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_195),
.B(n_197),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_36),
.B(n_34),
.C(n_33),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_165),
.Y(n_200)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_200),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_107),
.B(n_31),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_111),
.A2(n_39),
.B1(n_25),
.B2(n_33),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_132),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_205),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_115),
.A2(n_34),
.B1(n_30),
.B2(n_39),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_215),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_148),
.A2(n_47),
.B1(n_40),
.B2(n_31),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_130),
.A2(n_47),
.B1(n_40),
.B2(n_31),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_155),
.A2(n_40),
.B1(n_31),
.B2(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_11),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_18),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_137),
.B1(n_142),
.B2(n_134),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_120),
.A2(n_31),
.B1(n_12),
.B2(n_3),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_225),
.Y(n_234)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_9),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_132),
.A2(n_9),
.B(n_17),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_229),
.B(n_8),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_148),
.A2(n_9),
.B1(n_17),
.B2(n_3),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_0),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_139),
.A2(n_12),
.B1(n_17),
.B2(n_4),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_157),
.C(n_151),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_255),
.C(n_178),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_236),
.A2(n_261),
.B1(n_225),
.B2(n_200),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_169),
.A2(n_134),
.B1(n_146),
.B2(n_125),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_263),
.B1(n_269),
.B2(n_203),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_173),
.A2(n_159),
.B(n_150),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_243),
.A2(n_276),
.B(n_229),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_13),
.C(n_18),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_129),
.C(n_137),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_196),
.A2(n_158),
.B1(n_9),
.B2(n_4),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_174),
.A2(n_158),
.B1(n_13),
.B2(n_5),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_198),
.A2(n_186),
.B1(n_182),
.B2(n_211),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_186),
.A2(n_8),
.B1(n_16),
.B2(n_5),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_176),
.B(n_7),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_226),
.A2(n_7),
.B(n_8),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_219),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_180),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_280),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_204),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_15),
.B1(n_250),
.B2(n_231),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_287),
.A2(n_291),
.B(n_294),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_271),
.A2(n_215),
.B1(n_172),
.B2(n_171),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_181),
.B(n_189),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_245),
.A2(n_170),
.B1(n_183),
.B2(n_188),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_292),
.A2(n_296),
.B1(n_297),
.B2(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_260),
.B(n_271),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_245),
.A2(n_218),
.B1(n_192),
.B2(n_187),
.Y(n_297)
);

OA22x2_ASAP7_75t_L g361 ( 
.A1(n_298),
.A2(n_316),
.B1(n_327),
.B2(n_230),
.Y(n_361)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_299),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_175),
.B1(n_194),
.B2(n_193),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_301),
.A2(n_311),
.B1(n_318),
.B2(n_319),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_209),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_239),
.B(n_209),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_309),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_209),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_256),
.A2(n_199),
.B1(n_220),
.B2(n_195),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_281),
.A2(n_205),
.B1(n_197),
.B2(n_224),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_257),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_312),
.B(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_216),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_314),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_228),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_SL g316 ( 
.A1(n_260),
.A2(n_200),
.A3(n_184),
.B1(n_177),
.B2(n_223),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_317),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_213),
.B1(n_210),
.B2(n_208),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_266),
.A2(n_207),
.B1(n_206),
.B2(n_14),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_320),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_256),
.A2(n_0),
.B1(n_1),
.B2(n_14),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_330),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_269),
.A2(n_1),
.B1(n_15),
.B2(n_235),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_280),
.A2(n_1),
.B1(n_15),
.B2(n_235),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_254),
.B1(n_240),
.B2(n_231),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_238),
.B(n_1),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_325),
.B(n_248),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_326),
.A2(n_231),
.B1(n_232),
.B2(n_262),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_238),
.A2(n_243),
.B1(n_255),
.B2(n_242),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_276),
.A2(n_268),
.B(n_257),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_251),
.B(n_253),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_255),
.A2(n_242),
.B1(n_234),
.B2(n_268),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_351),
.B1(n_366),
.B2(n_283),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_251),
.B(n_253),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_333),
.A2(n_327),
.B(n_325),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_309),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_336),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_338),
.B(n_343),
.Y(n_382)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_339),
.A2(n_361),
.B(n_319),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_282),
.C(n_249),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_352),
.C(n_356),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_248),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_291),
.B(n_294),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_345),
.A2(n_354),
.B(n_293),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_312),
.B(n_249),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_346),
.B(n_355),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_302),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_349),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_292),
.A2(n_297),
.B1(n_316),
.B2(n_310),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_314),
.A2(n_254),
.B(n_267),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_267),
.C(n_240),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_285),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_364),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_230),
.B1(n_233),
.B2(n_241),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_344),
.B1(n_301),
.B2(n_366),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_288),
.C(n_313),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_322),
.A2(n_233),
.B1(n_241),
.B2(n_273),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_306),
.B(n_259),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_300),
.B(n_273),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_370),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_327),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_324),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_389),
.C(n_399),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_374),
.A2(n_362),
.B1(n_355),
.B2(n_360),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_375),
.A2(n_395),
.B1(n_401),
.B2(n_406),
.Y(n_416)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_363),
.A2(n_295),
.B(n_315),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_363),
.Y(n_413)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_387),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_388),
.B(n_394),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_311),
.Y(n_389)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_364),
.B(n_318),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_321),
.B1(n_296),
.B2(n_286),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_290),
.B1(n_284),
.B2(n_320),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_403),
.B1(n_336),
.B2(n_354),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_368),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_402),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_356),
.C(n_367),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_408),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_371),
.A2(n_326),
.B1(n_323),
.B2(n_305),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_359),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_365),
.A2(n_303),
.B1(n_307),
.B2(n_304),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_349),
.A2(n_304),
.B1(n_317),
.B2(n_299),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_347),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_293),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_405),
.Y(n_412)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_413),
.A2(n_380),
.B(n_406),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_345),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_426),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_424),
.B1(n_395),
.B2(n_398),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_348),
.C(n_339),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_425),
.C(n_427),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_422),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_386),
.A2(n_361),
.B1(n_348),
.B2(n_333),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_361),
.C(n_353),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_353),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_350),
.C(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_390),
.B(n_332),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_428),
.B(n_382),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_433),
.B1(n_439),
.B2(n_383),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_350),
.C(n_342),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_388),
.C(n_390),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_404),
.A2(n_357),
.B1(n_369),
.B2(n_372),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_436),
.B(n_384),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_397),
.A2(n_357),
.B1(n_369),
.B2(n_347),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_389),
.B(n_357),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_394),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_441),
.A2(n_456),
.B1(n_461),
.B2(n_430),
.Y(n_478)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_392),
.Y(n_445)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_446),
.B(n_467),
.Y(n_479)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

FAx1_ASAP7_75t_SL g449 ( 
.A(n_429),
.B(n_400),
.CI(n_408),
.CON(n_449),
.SN(n_449)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_457),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_424),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_407),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_466),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_376),
.Y(n_453)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_465),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_411),
.B(n_386),
.C(n_387),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_427),
.C(n_431),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_423),
.A2(n_401),
.B1(n_375),
.B2(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_376),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_464),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_393),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_437),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_416),
.A2(n_402),
.B1(n_381),
.B2(n_385),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_377),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_440),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_477),
.C(n_482),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_453),
.B(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_463),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_425),
.C(n_420),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_461),
.B1(n_456),
.B2(n_441),
.Y(n_499)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_423),
.C(n_458),
.Y(n_481)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_436),
.C(n_414),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_414),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_484),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_429),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_446),
.B(n_416),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_486),
.B(n_487),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_488),
.B(n_471),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_495),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_457),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_496),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_447),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_489),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_486),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_504),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_471),
.B(n_483),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_501),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_466),
.C(n_460),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_502),
.B(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_443),
.C(n_452),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_474),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_443),
.C(n_467),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_506),
.Y(n_519)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_479),
.B(n_449),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_476),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_491),
.A2(n_470),
.B(n_485),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_515),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_494),
.A2(n_465),
.B(n_478),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_517),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_490),
.B(n_484),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_516),
.A2(n_500),
.B1(n_507),
.B2(n_449),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_497),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_521),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_487),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_508),
.A2(n_496),
.B1(n_499),
.B2(n_498),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_528),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_503),
.C(n_502),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_525),
.B(n_526),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_476),
.C(n_498),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_514),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_529),
.B(n_530),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_510),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_448),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_531),
.B(n_480),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_510),
.A2(n_464),
.B(n_409),
.Y(n_532)
);

AOI21x1_ASAP7_75t_L g537 ( 
.A1(n_532),
.A2(n_524),
.B(n_523),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_525),
.A2(n_511),
.B(n_513),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_533),
.A2(n_517),
.B(n_434),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_521),
.C(n_516),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_539),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_SL g543 ( 
.A1(n_537),
.A2(n_479),
.B(n_434),
.C(n_415),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_538),
.A2(n_522),
.B(n_526),
.Y(n_541)
);

MAJx2_ASAP7_75t_L g544 ( 
.A(n_541),
.B(n_543),
.C(n_535),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_534),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_545),
.B(n_540),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_545),
.A2(n_539),
.B(n_435),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_438),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_438),
.C(n_299),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_317),
.Y(n_551)
);


endmodule