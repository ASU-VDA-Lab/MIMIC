module real_jpeg_16810_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_155;
wire n_120;
wire n_572;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_1),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_1),
.B(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_145),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

NAND2x1_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_2),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_2),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_2),
.B(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_3),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_5),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_7),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_7),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_7),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_7),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_7),
.B(n_145),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_7),
.B(n_147),
.Y(n_451)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

BUFx4f_ASAP7_75t_L g259 ( 
.A(n_8),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_8),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_9),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_9),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_9),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_9),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_9),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_9),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_9),
.B(n_496),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_10),
.B(n_58),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_10),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_155),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_10),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_10),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_11),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_11),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_11),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_11),
.B(n_209),
.Y(n_351)
);

AOI22x1_ASAP7_75t_L g152 ( 
.A1(n_12),
.A2(n_15),
.B1(n_153),
.B2(n_157),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_12),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_12),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_12),
.B(n_305),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g380 ( 
.A1(n_12),
.A2(n_152),
.A3(n_381),
.B(n_384),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_12),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_12),
.B(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_12),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_12),
.B(n_483),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_13),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_14),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_14),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_14),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_14),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_14),
.B(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_14),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_14),
.B(n_156),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

NAND2x1_ASAP7_75t_L g346 ( 
.A(n_15),
.B(n_347),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_15),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_16),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_16),
.Y(n_277)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_16),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_578),
.B(n_586),
.C(n_588),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_127),
.B(n_577),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_80),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_27),
.B(n_80),
.Y(n_577)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_27),
.Y(n_590)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_46),
.CI(n_60),
.CON(n_27),
.SN(n_27)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_28),
.B(n_46),
.C(n_60),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.C(n_40),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_29),
.A2(n_35),
.B1(n_53),
.B2(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g580 ( 
.A(n_29),
.B(n_48),
.C(n_55),
.Y(n_580)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_34),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_70),
.C(n_75),
.Y(n_69)
);

AOI22x1_ASAP7_75t_L g122 ( 
.A1(n_35),
.A2(n_64),
.B1(n_75),
.B2(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_39),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_55),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_48),
.A2(n_54),
.B1(n_582),
.B2(n_586),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_116),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_52),
.B(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.C(n_69),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_61),
.A2(n_62),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_65),
.B(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2x1_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_73),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_75),
.A2(n_76),
.B1(n_115),
.B2(n_338),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_111),
.C(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_79),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_123),
.C(n_124),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_81),
.B(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_110),
.C(n_120),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_82),
.B(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_88),
.C(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_87),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.C(n_107),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_92),
.A2(n_93),
.B1(n_100),
.B2(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_99),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_99),
.Y(n_336)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_101),
.Y(n_541)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_105),
.Y(n_228)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_105),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_107),
.B(n_540),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_110),
.B(n_121),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_111),
.B(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_115),
.A2(n_257),
.B1(n_260),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_115),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_115),
.B(n_260),
.C(n_333),
.Y(n_546)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_119),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_123),
.B(n_124),
.Y(n_552)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_532),
.B(n_572),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_365),
.B(n_529),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_326),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_280),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_131),
.B(n_280),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_204),
.Y(n_131)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_132),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_169),
.C(n_192),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_134),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.C(n_161),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_135),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g542 ( 
.A(n_136),
.B(n_248),
.C(n_358),
.Y(n_542)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_137),
.B(n_248),
.Y(n_355)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_142),
.C(n_146),
.Y(n_195)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_140),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_145),
.Y(n_298)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_151),
.A2(n_152),
.B1(n_161),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_161),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_162),
.A2(n_163),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_163),
.B(n_235),
.C(n_257),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_166),
.B(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_168),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_170),
.A2(n_193),
.B1(n_194),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_170),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_182),
.C(n_187),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_171),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_172),
.A2(n_178),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_172),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_172),
.B(n_432),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_174),
.Y(n_479)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_176),
.B(n_377),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_178),
.Y(n_379)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_180),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_187),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_197),
.C(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_197),
.A2(n_198),
.B1(n_393),
.B2(n_394),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_198),
.Y(n_392)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_203),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_253),
.B1(n_278),
.B2(n_279),
.Y(n_204)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_243),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g328 ( 
.A(n_206),
.B(n_244),
.C(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.C(n_229),
.Y(n_206)
);

XNOR2x2_ASAP7_75t_SL g286 ( 
.A(n_207),
.B(n_287),
.Y(n_286)
);

XOR2x1_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_211),
.C(n_214),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_217),
.B(n_229),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_218),
.A2(n_226),
.B1(n_227),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_218),
.Y(n_325)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_221),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_222),
.B(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_226),
.B(n_412),
.C(n_414),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_226),
.A2(n_227),
.B1(n_412),
.B2(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_235),
.C(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_235),
.A2(n_242),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_236),
.Y(n_387)
);

INVx6_ASAP7_75t_L g484 ( 
.A(n_236),
.Y(n_484)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_246),
.B(n_252),
.C(n_360),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_248),
.Y(n_360)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_253),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_254),
.B(n_262),
.C(n_264),
.Y(n_361)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_257),
.Y(n_260)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_258),
.Y(n_450)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_259),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_265),
.B(n_270),
.C(n_274),
.Y(n_340)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_363),
.C(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.C(n_288),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_289),
.B(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_319),
.C(n_323),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_290),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.C(n_303),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_SL g419 ( 
.A(n_292),
.B(n_420),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_295),
.B(n_303),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_296),
.B(n_300),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.C(n_314),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_304),
.A2(n_310),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_304),
.Y(n_408)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_310),
.A2(n_409),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_310),
.B(n_477),
.C(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2x1_ASAP7_75t_SL g406 ( 
.A(n_314),
.B(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_323),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_326),
.A2(n_530),
.B(n_531),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_362),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_327),
.B(n_362),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_328),
.B(n_331),
.C(n_352),
.Y(n_568)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_352),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_339),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_332),
.B(n_340),
.C(n_341),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_342),
.B(n_346),
.C(n_351),
.Y(n_547)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_361),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_354),
.B(n_359),
.C(n_566),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_356),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_361),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_423),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.C(n_400),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_372),
.Y(n_425)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.C(n_396),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_373),
.B(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_397),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_380),
.C(n_388),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_380),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_433),
.C(n_437),
.Y(n_456)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_393),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_389),
.B(n_518),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_SL g463 ( 
.A(n_390),
.B(n_391),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_390),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_390),
.A2(n_481),
.B1(n_482),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_421),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_421),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_419),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_402),
.B(n_527),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_405),
.B(n_419),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.C(n_417),
.Y(n_405)
);

XOR2x1_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_418),
.Y(n_513)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

XOR2x2_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_458),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.C(n_426),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_427),
.A2(n_524),
.B(n_528),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_509),
.B(n_523),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_471),
.B(n_508),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_454),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_430),
.B(n_454),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_439),
.C(n_448),
.Y(n_430)
);

XOR2x1_ASAP7_75t_SL g502 ( 
.A(n_431),
.B(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_437),
.Y(n_432)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_439),
.A2(n_440),
.B1(n_448),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_447),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_447),
.Y(n_475)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

AO22x1_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_449),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_451),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_452),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_495),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_456),
.B(n_457),
.C(n_522),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_460),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g520 ( 
.A(n_461),
.B(n_463),
.C(n_464),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx6_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_501),
.B(n_507),
.Y(n_471)
);

OAI21x1_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_485),
.B(n_500),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_480),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_482),
.Y(n_493)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_494),
.B(n_499),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_492),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_492),
.Y(n_499)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_505),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_521),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_521),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_512),
.B1(n_514),
.B2(n_515),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_516),
.C(n_520),
.Y(n_525)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_526),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_SL g532 ( 
.A(n_533),
.B(n_553),
.C(n_567),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_533),
.A2(n_573),
.B(n_576),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_R g533 ( 
.A(n_534),
.B(n_551),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_551),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_543),
.C(n_548),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_556),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_538),
.C(n_542),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_537),
.B(n_562),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_542),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_543),
.A2(n_548),
.B1(n_549),
.B2(n_557),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_543),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_546),
.C(n_547),
.Y(n_543)
);

XNOR2x2_ASAP7_75t_SL g563 ( 
.A(n_544),
.B(n_564),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_547),
.Y(n_564)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_554),
.A2(n_574),
.B(n_575),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_558),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_558),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_563),
.C(n_565),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_560),
.A2(n_561),
.B1(n_563),
.B2(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_563),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_570),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_569),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_SL g574 ( 
.A(n_568),
.B(n_569),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_R g578 ( 
.A(n_579),
.B(n_587),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_579),
.B(n_587),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_581),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_582),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_584),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_589),
.Y(n_588)
);


endmodule