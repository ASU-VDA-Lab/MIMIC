module fake_jpeg_14510_n_425 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_425);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_58),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_66),
.Y(n_123)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_27),
.B(n_16),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_17),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_75),
.Y(n_171)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_82),
.Y(n_115)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_14),
.B1(n_12),
.B2(n_4),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_21),
.B1(n_52),
.B2(n_49),
.Y(n_165)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_28),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_83),
.B(n_85),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_1),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_87),
.B(n_89),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_39),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_2),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_93),
.B(n_99),
.Y(n_138)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_5),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_35),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_38),
.A2(n_5),
.B(n_6),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_25),
.Y(n_150)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_24),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_48),
.B1(n_23),
.B2(n_54),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_112),
.A2(n_119),
.B1(n_122),
.B2(n_125),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_113),
.A2(n_151),
.B1(n_74),
.B2(n_91),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_61),
.A2(n_48),
.B1(n_54),
.B2(n_51),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_24),
.B1(n_20),
.B2(n_46),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_124),
.B(n_126),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_139),
.A2(n_173),
.B1(n_174),
.B2(n_125),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_142),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_118),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_67),
.B1(n_107),
.B2(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_56),
.B(n_41),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_25),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_160),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_21),
.B(n_52),
.C(n_49),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_171),
.B(n_170),
.C(n_134),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_112),
.B1(n_119),
.B2(n_122),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_57),
.A2(n_60),
.B1(n_95),
.B2(n_92),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_73),
.A2(n_18),
.B1(n_40),
.B2(n_36),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_36),
.B1(n_40),
.B2(n_53),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_178),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_53),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_182),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_180),
.A2(n_208),
.B1(n_200),
.B2(n_185),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_59),
.B1(n_109),
.B2(n_98),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_86),
.B(n_110),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_194),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_9),
.C(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_217),
.C(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_156),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_192),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_195),
.A2(n_196),
.B1(n_218),
.B2(n_227),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_175),
.B1(n_145),
.B2(n_163),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_198),
.A2(n_200),
.B1(n_203),
.B2(n_190),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_154),
.B1(n_166),
.B2(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_210),
.B1(n_214),
.B2(n_220),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_139),
.B1(n_159),
.B2(n_175),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_212),
.B1(n_180),
.B2(n_213),
.Y(n_243)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_215),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_153),
.A2(n_136),
.B1(n_162),
.B2(n_130),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_123),
.B(n_154),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_143),
.B1(n_114),
.B2(n_146),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_225),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_134),
.A2(n_170),
.B(n_143),
.C(n_128),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_128),
.B(n_144),
.C(n_132),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_217),
.B(n_212),
.C(n_228),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_146),
.A2(n_164),
.B1(n_131),
.B2(n_120),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_132),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_136),
.A2(n_162),
.B1(n_147),
.B2(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_144),
.A2(n_48),
.B1(n_23),
.B2(n_84),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_116),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_228),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_112),
.A2(n_165),
.B1(n_119),
.B2(n_122),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_171),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_142),
.A2(n_48),
.B1(n_23),
.B2(n_84),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_192),
.B1(n_198),
.B2(n_232),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_252),
.B1(n_255),
.B2(n_258),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_256),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_225),
.B(n_179),
.C(n_194),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_257),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_200),
.A2(n_184),
.B1(n_211),
.B2(n_189),
.Y(n_255)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_203),
.B(n_204),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_222),
.C(n_229),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_184),
.A2(n_186),
.B1(n_221),
.B2(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_177),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_272),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_221),
.B(n_217),
.C(n_191),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_269),
.B(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_205),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_230),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_193),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_193),
.A2(n_232),
.B1(n_212),
.B2(n_202),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_201),
.B(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_253),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_222),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_278),
.B(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_285),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_258),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_249),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_288),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_246),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_244),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_293),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_294),
.Y(n_319)
);

AOI32xp33_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_236),
.A3(n_251),
.B1(n_255),
.B2(n_267),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_302),
.B(n_307),
.C(n_248),
.D(n_234),
.Y(n_323)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_250),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_235),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_271),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_256),
.C(n_259),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_242),
.B(n_257),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_242),
.B(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_239),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_277),
.A2(n_266),
.B1(n_243),
.B2(n_233),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_313),
.A2(n_314),
.B1(n_318),
.B2(n_332),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_266),
.B1(n_241),
.B2(n_243),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_284),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_329),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_243),
.B1(n_270),
.B2(n_265),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_318),
.A2(n_308),
.B1(n_280),
.B2(n_285),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_270),
.B1(n_256),
.B2(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_326),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_333),
.C(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_323),
.B(n_291),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_234),
.B1(n_240),
.B2(n_277),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_283),
.C(n_300),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_297),
.A2(n_286),
.B(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_297),
.B(n_289),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_292),
.CI(n_306),
.CON(n_329),
.SN(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_303),
.B1(n_283),
.B2(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_332),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_280),
.B1(n_297),
.B2(n_308),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_304),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_340),
.C(n_347),
.Y(n_357)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_342),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_339),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_307),
.C(n_278),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_328),
.A2(n_288),
.B(n_301),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_309),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_293),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_315),
.C(n_319),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_317),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_349),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_350),
.A2(n_351),
.B1(n_355),
.B2(n_338),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_324),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_279),
.B(n_285),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_343),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_312),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_353),
.A2(n_313),
.B1(n_316),
.B2(n_319),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_356),
.A2(n_370),
.B1(n_342),
.B2(n_352),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_327),
.Y(n_358)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_344),
.B(n_336),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_365),
.C(n_367),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_369),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_319),
.C(n_311),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_311),
.C(n_329),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_310),
.B1(n_325),
.B2(n_279),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_323),
.C(n_326),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_336),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_384),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_380),
.B1(n_381),
.B2(n_347),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_366),
.A2(n_353),
.B1(n_337),
.B2(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_345),
.B(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_342),
.B1(n_335),
.B2(n_345),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_364),
.A2(n_341),
.B1(n_355),
.B2(n_310),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_350),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx11_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_346),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_348),
.Y(n_384)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_385),
.B(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_390),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_380),
.A2(n_375),
.B1(n_381),
.B2(n_378),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_371),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_394),
.C(n_395),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_325),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_365),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_396),
.B(n_385),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_398),
.B(n_399),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_401),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g401 ( 
.A1(n_386),
.A2(n_369),
.B(n_363),
.C(n_358),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_392),
.A2(n_373),
.B(n_367),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_373),
.B(n_379),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_403),
.B(n_340),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_406),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_407),
.B(n_405),
.Y(n_416)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_388),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_411),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_395),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_387),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_412),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_416),
.B(n_394),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_415),
.B(n_405),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_419),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_417),
.B(n_414),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_408),
.C(n_413),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_420),
.B(n_415),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_382),
.B1(n_406),
.B2(n_383),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_411),
.Y(n_425)
);


endmodule