module fake_jpeg_7183_n_176 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_36),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_23),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_28),
.B(n_19),
.C(n_14),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_25),
.B(n_18),
.C(n_20),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_67),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_24),
.B1(n_18),
.B2(n_20),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_61),
.A3(n_51),
.B1(n_50),
.B2(n_63),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_13),
.C(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_21),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_32),
.C(n_35),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.C(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_27),
.B1(n_72),
.B2(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_51),
.B(n_21),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_60),
.C(n_44),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_54),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_32),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_56),
.C(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_36),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_26),
.Y(n_130)
);

XOR2x2_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_66),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_102),
.B1(n_109),
.B2(n_89),
.C(n_92),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_69),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_83),
.B(n_92),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_15),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_30),
.B1(n_39),
.B2(n_22),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_113),
.B1(n_83),
.B2(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_26),
.B1(n_41),
.B2(n_15),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_123),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_118),
.B1(n_96),
.B2(n_113),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_76),
.A3(n_90),
.B1(n_78),
.B2(n_93),
.C1(n_75),
.C2(n_85),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_126),
.A3(n_105),
.B1(n_112),
.B2(n_98),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_78),
.B(n_80),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_85),
.B(n_88),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_130),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_77),
.B1(n_86),
.B2(n_26),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_111),
.B(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_128),
.B1(n_119),
.B2(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_115),
.B1(n_122),
.B2(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_139),
.B(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_13),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_98),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_132),
.B1(n_142),
.B2(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_6),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_121),
.B1(n_125),
.B2(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_116),
.C(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_15),
.C(n_3),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_139),
.B(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_159),
.B1(n_8),
.B2(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_0),
.B(n_5),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_7),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_6),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_151),
.C(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_164),
.C(n_154),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_9),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_7),
.C(n_8),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_156),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_163),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_154),
.B(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.C(n_160),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_11),
.CI(n_171),
.CON(n_174),
.SN(n_174)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_9),
.B(n_10),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.C(n_11),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);


endmodule