module fake_jpeg_29106_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_1),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_19),
.Y(n_84)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_17),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_71),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.C(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_20),
.CI(n_23),
.CON(n_86),
.SN(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_24),
.B(n_25),
.Y(n_88)
);

AO21x2_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_26),
.B(n_27),
.Y(n_89)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_79),
.C(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_93),
.C(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_99),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_98),
.B(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_96),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_78),
.C(n_89),
.Y(n_110)
);


endmodule