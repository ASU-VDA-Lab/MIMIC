module fake_ariane_1843_n_131 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_131);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_131;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_124;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_117;
wire n_85;
wire n_130;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_122;
wire n_52;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_87;
wire n_81;
wire n_29;
wire n_41;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_11),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_0),
.Y(n_51)
);

OR2x6_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_47),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_7),
.B(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_9),
.C(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_11),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_48),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_50),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_52),
.B2(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_64),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_50),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_35),
.B1(n_42),
.B2(n_39),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_65),
.B(n_54),
.C(n_45),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_77),
.Y(n_85)
);

AO21x2_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_68),
.B(n_62),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_78),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_62),
.B(n_46),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_53),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_40),
.B1(n_43),
.B2(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_74),
.B(n_76),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_72),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_91),
.B1(n_86),
.B2(n_80),
.Y(n_102)
);

OR2x6_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_108),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_38),
.A3(n_32),
.B1(n_31),
.B2(n_81),
.C1(n_102),
.C2(n_39),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_112),
.Y(n_117)
);

OAI211xp5_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_83),
.B(n_95),
.C(n_96),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_110),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_60),
.C(n_89),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_121),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_86),
.B1(n_87),
.B2(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_88),
.Y(n_128)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_98),
.B1(n_97),
.B2(n_84),
.C(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_129),
.B1(n_18),
.B2(n_20),
.C(n_25),
.Y(n_131)
);


endmodule