module fake_jpeg_4902_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_15),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_64),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_37),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_71),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_76),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_36),
.B1(n_26),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_101),
.B1(n_69),
.B2(n_53),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_45),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_26),
.B1(n_40),
.B2(n_36),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_60),
.Y(n_113)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_54),
.B1(n_69),
.B2(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_82),
.B1(n_77),
.B2(n_83),
.Y(n_150)
);

OAI31xp33_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_25),
.A3(n_57),
.B(n_62),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_121),
.B1(n_50),
.B2(n_67),
.Y(n_137)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_70),
.CI(n_57),
.CON(n_112),
.SN(n_112)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_113),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_25),
.B(n_51),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_123),
.B1(n_128),
.B2(n_132),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_46),
.B1(n_38),
.B2(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_122),
.B1(n_116),
.B2(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_68),
.B1(n_51),
.B2(n_61),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_61),
.B1(n_67),
.B2(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_41),
.B(n_43),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_43),
.C(n_23),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_159),
.Y(n_167)
);

CKINVDCx10_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_145),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_117),
.B1(n_110),
.B2(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_96),
.B1(n_126),
.B2(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_158),
.B(n_34),
.Y(n_178)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_63),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_127),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_33),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_115),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_131),
.C(n_128),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_166),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_112),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_168),
.B(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_164),
.B1(n_177),
.B2(n_88),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_112),
.B1(n_117),
.B2(n_46),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_110),
.B(n_92),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

OAI22x1_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_76),
.B1(n_74),
.B2(n_46),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_179),
.B1(n_184),
.B2(n_108),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_118),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_158),
.B1(n_160),
.B2(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_186),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_136),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_85),
.B(n_118),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_42),
.B(n_27),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_102),
.B(n_27),
.Y(n_194)
);

OAI22x1_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_76),
.B1(n_42),
.B2(n_97),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_104),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_201),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_190),
.B(n_192),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_140),
.B1(n_152),
.B2(n_135),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_155),
.B(n_149),
.Y(n_192)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_205),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_32),
.B(n_18),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_202),
.B1(n_214),
.B2(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_93),
.B1(n_141),
.B2(n_108),
.Y(n_202)
);

NAND2x1_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_27),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_27),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_192),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_30),
.B(n_20),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_35),
.B(n_31),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_156),
.B1(n_142),
.B2(n_30),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_171),
.B1(n_167),
.B2(n_173),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_210),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_22),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_104),
.C(n_27),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_30),
.B1(n_32),
.B2(n_18),
.Y(n_214)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_193),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_221),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_180),
.B1(n_162),
.B2(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_203),
.B1(n_198),
.B2(n_200),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_173),
.B1(n_181),
.B2(n_165),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_232),
.B1(n_238),
.B2(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_234),
.C(n_195),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_181),
.B1(n_172),
.B2(n_35),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_198),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_191),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_172),
.C(n_104),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_19),
.B(n_28),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_214),
.B(n_205),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_19),
.B1(n_31),
.B2(n_28),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_97),
.B1(n_87),
.B2(n_107),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_245),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_200),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_242),
.B(n_247),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_195),
.B1(n_190),
.B2(n_211),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_209),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_261),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_107),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_97),
.B1(n_87),
.B2(n_29),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_222),
.B1(n_87),
.B2(n_224),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_29),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_0),
.B(n_1),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_232),
.B1(n_238),
.B2(n_235),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_262),
.B1(n_260),
.B2(n_259),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_254),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_217),
.C(n_226),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_236),
.C(n_230),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_216),
.C(n_223),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_241),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_221),
.C(n_29),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_279),
.B(n_281),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_29),
.C(n_24),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_292),
.C(n_282),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_298),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_266),
.A2(n_258),
.B(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_287),
.A2(n_299),
.B(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

XOR2x1_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_244),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_277),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_283),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_254),
.C(n_261),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_282),
.B1(n_279),
.B2(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_272),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_301),
.C(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_267),
.C(n_269),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_275),
.B1(n_246),
.B2(n_263),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_3),
.C(n_4),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_283),
.B1(n_11),
.B2(n_12),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_284),
.B(n_289),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_24),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_1),
.C(n_3),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_3),
.C(n_4),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_305),
.B1(n_306),
.B2(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_320),
.C(n_321),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_317),
.B(n_319),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_11),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_24),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_4),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_301),
.A2(n_13),
.B(n_12),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_310),
.C(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_5),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_328),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_300),
.B(n_5),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_321),
.C(n_6),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_24),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_330),
.C(n_5),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_4),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_5),
.B(n_6),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_338),
.B(n_331),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_318),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_337),
.Y(n_340)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_325),
.A2(n_318),
.B1(n_24),
.B2(n_8),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_339),
.Y(n_342)
);

OAI21x1_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_341),
.B(n_336),
.Y(n_343)
);

AOI222xp33_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_340),
.C2(n_338),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_7),
.B(n_8),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_7),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_7),
.Y(n_347)
);


endmodule