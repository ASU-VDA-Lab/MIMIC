module real_jpeg_10762_n_12 (n_5, n_4, n_8, n_0, n_283, n_1, n_11, n_2, n_284, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_283;
input n_1;
input n_11;
input n_2;
input n_284;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_11),
.B1(n_19),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_1),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_30),
.B1(n_64),
.B2(n_65),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_9),
.B(n_27),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_40),
.B(n_63),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_9),
.B(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_8),
.A2(n_11),
.B1(n_19),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_11),
.B1(n_19),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_9),
.A2(n_51),
.B1(n_64),
.B2(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_40),
.B1(n_42),
.B2(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_37),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_26),
.B(n_39),
.C(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_28),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_11),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_10),
.A2(n_20),
.B1(n_64),
.B2(n_65),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_20),
.B1(n_40),
.B2(n_42),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_23),
.B(n_51),
.C(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_73),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_72),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_31),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_18),
.A2(n_25),
.B(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_22),
.A2(n_25),
.B1(n_50),
.B2(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_22),
.B(n_25),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_38),
.B(n_39),
.C(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_28),
.A2(n_49),
.B(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_32),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_32),
.B(n_280),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_47),
.CI(n_52),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_37),
.B1(n_44),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_36),
.B(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_37),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_37),
.A2(n_44),
.B1(n_129),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_38),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_40),
.A2(n_43),
.B(n_51),
.Y(n_135)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_51),
.B(n_68),
.C(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_45),
.B(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_50),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_51),
.B(n_63),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.C(n_60),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_53),
.A2(n_60),
.B1(n_260),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_53),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_54),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_55),
.A2(n_56),
.B1(n_145),
.B2(n_151),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_55),
.B(n_145),
.C(n_188),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_55),
.A2(n_56),
.B1(n_128),
.B2(n_132),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_55),
.B(n_128),
.C(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_55),
.A2(n_56),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_60),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_69),
.B1(n_94),
.B2(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_223),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_279),
.B(n_281),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_252),
.A3(n_272),
.B1(n_277),
.B2(n_278),
.C(n_283),
.Y(n_74)
);

AOI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_207),
.A3(n_227),
.B1(n_246),
.B2(n_251),
.C(n_284),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_176),
.C(n_204),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_156),
.B(n_175),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_141),
.B(n_155),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_123),
.B(n_140),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_112),
.B(n_122),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_102),
.B(n_111),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_91),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_83),
.A2(n_104),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_83),
.B(n_145),
.C(n_150),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_86),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_86),
.A2(n_138),
.B1(n_183),
.B2(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_88),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_89),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_101),
.B1(n_128),
.B2(n_132),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_128),
.C(n_139),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_101),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_97),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_101),
.B(n_181),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B(n_110),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_117),
.C(n_120),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_121),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_114),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_120),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_119),
.A2(n_120),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_195),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_144),
.C(n_154),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_133),
.B2(n_139),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_128),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_132),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_162),
.C(n_166),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_130),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_143),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_152),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_151),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_233),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_158),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_168),
.C(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_165),
.B2(n_166),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_166),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_165),
.A2(n_166),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_165),
.A2(n_166),
.B1(n_266),
.B2(n_270),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_165),
.B(n_260),
.C(n_261),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_165),
.B(n_270),
.C(n_271),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_199),
.C(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_178),
.B(n_189),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_185),
.CI(n_186),
.CON(n_178),
.SN(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_203),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_198),
.C(n_203),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_247),
.B(n_250),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_209),
.B(n_210),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_226),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_219),
.C(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_221),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_222),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_236),
.B(n_238),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_244),
.B2(n_245),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_232),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_243),
.C(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_254),
.C(n_262),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_254),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_264),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_264),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_257),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_263),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);


endmodule