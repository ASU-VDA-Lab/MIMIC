module fake_netlist_5_1501_n_1741 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1741);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1741;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_51),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_57),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_4),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_98),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_20),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_37),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_86),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_43),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_92),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_68),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_13),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_42),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_79),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_32),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_112),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_21),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_0),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_130),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_49),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_105),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_88),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_35),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_50),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_123),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_14),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_60),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_25),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_122),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_89),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_154),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_39),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_55),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_23),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_91),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_144),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_120),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_107),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_96),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_145),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_87),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_40),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

HB1xp67_ASAP7_75t_SL g258 ( 
.A(n_28),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_117),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_58),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_158),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_6),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_85),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_95),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_55),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_135),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_101),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_0),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_42),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_77),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_82),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_67),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_28),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_148),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_34),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_75),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_34),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_115),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_151),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_147),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_16),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_3),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_17),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_119),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_125),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_7),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_44),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_14),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_84),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_70),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_22),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_56),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_30),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_27),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_141),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_83),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_16),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_146),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_171),
.B(n_1),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_4),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_306),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_222),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_222),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_262),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_309),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_171),
.B(n_5),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_222),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_222),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_212),
.B(n_237),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_183),
.B(n_7),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_225),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_165),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_212),
.B(n_8),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_246),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_193),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_165),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_298),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_160),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_167),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_172),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_163),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_172),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_173),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_173),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_225),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_180),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_174),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_184),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_175),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_166),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_169),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_184),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_170),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_205),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_225),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_176),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_261),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_205),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_232),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_237),
.B(n_9),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_261),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_210),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_179),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_186),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_210),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_181),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_182),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_188),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_189),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_185),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_190),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_211),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_191),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_183),
.B(n_9),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_187),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_225),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_322),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_169),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_349),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_352),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_339),
.B(n_276),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_363),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

CKINVDCx8_ASAP7_75t_R g402 ( 
.A(n_320),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_281),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_276),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_366),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_369),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_391),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_386),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_329),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_291),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_321),
.B(n_195),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_335),
.B(n_194),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_291),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_341),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_333),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_334),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_347),
.B(n_307),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_336),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_336),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_338),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_307),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_353),
.B(n_178),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_354),
.B(n_219),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_385),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_377),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_390),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_342),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_350),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_350),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_330),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_358),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_375),
.B1(n_319),
.B2(n_374),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_394),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_427),
.B(n_344),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_395),
.B(n_387),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_431),
.A2(n_346),
.B1(n_348),
.B2(n_323),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_426),
.B(n_358),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_395),
.B(n_362),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_431),
.A2(n_370),
.B1(n_376),
.B2(n_234),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_211),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_362),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_448),
.A2(n_370),
.B1(n_376),
.B2(n_234),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_397),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_379),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_460),
.B(n_345),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_396),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_419),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_444),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_379),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_439),
.B(n_219),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_383),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_439),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_429),
.B(n_383),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_419),
.B(n_384),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_463),
.B(n_384),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_226),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_413),
.B(n_388),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_413),
.B(n_226),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_411),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_453),
.B(n_388),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_440),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_461),
.B(n_278),
.C(n_215),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_440),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_394),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_461),
.B(n_393),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_393),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_448),
.B(n_229),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_440),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_453),
.B(n_218),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_429),
.B(n_178),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_421),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_437),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_437),
.B(n_268),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_421),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_461),
.B(n_465),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_448),
.A2(n_224),
.B1(n_242),
.B2(n_168),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_448),
.A2(n_278),
.B1(n_316),
.B2(n_332),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_448),
.A2(n_316),
.B1(n_337),
.B2(n_318),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_465),
.B(n_196),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_331),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_453),
.B(n_199),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_453),
.B(n_201),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_402),
.B(n_437),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

NOR2x1p5_ASAP7_75t_L g559 ( 
.A(n_400),
.B(n_268),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_405),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_405),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_446),
.A2(n_389),
.B1(n_304),
.B2(n_310),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_434),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_405),
.B(n_281),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_403),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_434),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_451),
.B(n_343),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_420),
.A2(n_275),
.B1(n_256),
.B2(n_208),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_402),
.B(n_204),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_404),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_446),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_404),
.B(n_206),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_406),
.B(n_207),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_454),
.B(n_238),
.C(n_229),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_454),
.B(n_200),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_455),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_402),
.B(n_446),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_447),
.B(n_317),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_447),
.B(n_213),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_455),
.A2(n_304),
.B1(n_310),
.B2(n_312),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_406),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_457),
.B(n_238),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_457),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_407),
.B(n_214),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_462),
.A2(n_233),
.B1(n_239),
.B2(n_236),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_398),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_396),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_396),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_407),
.B(n_223),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_405),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_396),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_399),
.B(n_164),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_408),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_408),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_410),
.B(n_230),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_405),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_399),
.B(n_281),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_410),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_401),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_456),
.A2(n_269),
.B1(n_216),
.B2(n_312),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_409),
.A2(n_265),
.B1(n_203),
.B2(n_221),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_412),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_412),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_456),
.B(n_281),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_456),
.A2(n_269),
.B1(n_192),
.B2(n_308),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_449),
.B(n_240),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_456),
.B(n_240),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_409),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_417),
.B(n_231),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_449),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_613),
.B(n_458),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_613),
.B(n_458),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_489),
.B(n_591),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_537),
.B(n_297),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_458),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_537),
.B(n_297),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_400),
.C(n_443),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_258),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_486),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_415),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_615),
.B(n_573),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_534),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_487),
.B(n_202),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_228),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_467),
.B(n_458),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_501),
.B(n_476),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_466),
.B(n_297),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_466),
.B(n_297),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_500),
.Y(n_636)
);

NAND2x1p5_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_241),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_534),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_539),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_466),
.B(n_297),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_539),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_489),
.B(n_416),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

OAI221xp5_ASAP7_75t_L g647 ( 
.A1(n_468),
.A2(n_313),
.B1(n_263),
.B2(n_284),
.C(n_255),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_467),
.B(n_417),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_580),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_502),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_476),
.B(n_241),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_498),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_482),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_591),
.B(n_418),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_482),
.B(n_244),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_469),
.B(n_425),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_572),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_472),
.B(n_473),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_529),
.B(n_443),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_468),
.A2(n_259),
.B1(n_280),
.B2(n_274),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_597),
.A2(n_255),
.B(n_192),
.C(n_198),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_570),
.A2(n_464),
.B1(n_459),
.B2(n_450),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_490),
.B(n_257),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_500),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_473),
.B(n_422),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_466),
.B(n_297),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_490),
.B(n_260),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_479),
.B(n_484),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_580),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_SL g671 ( 
.A(n_561),
.B(n_244),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_518),
.B(n_297),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_484),
.B(n_422),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_597),
.A2(n_284),
.B(n_263),
.C(n_242),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_609),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_492),
.B(n_248),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_483),
.B(n_282),
.C(n_270),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_494),
.B(n_248),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_518),
.B(n_297),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_590),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_518),
.B(n_297),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_494),
.B(n_495),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_572),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_495),
.B(n_250),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_498),
.B(n_423),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_481),
.A2(n_283),
.B1(n_243),
.B2(n_245),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_481),
.A2(n_293),
.B1(n_273),
.B2(n_271),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_529),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_505),
.B(n_432),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_488),
.B(n_287),
.C(n_279),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_505),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_585),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_517),
.B(n_277),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_542),
.B(n_286),
.C(n_301),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_508),
.B(n_509),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_497),
.B(n_285),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_590),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_557),
.B(n_581),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_598),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_599),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_497),
.B(n_288),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_508),
.A2(n_302),
.B1(n_272),
.B2(n_264),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_499),
.B(n_288),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_536),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_499),
.B(n_294),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_533),
.B(n_294),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_530),
.B(n_300),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_599),
.B(n_607),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_607),
.B(n_300),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_475),
.B(n_566),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_518),
.B(n_209),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_554),
.B(n_247),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_549),
.B(n_289),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_578),
.A2(n_168),
.B(n_249),
.C(n_198),
.Y(n_717)
);

OAI221xp5_ASAP7_75t_L g718 ( 
.A1(n_605),
.A2(n_224),
.B1(n_220),
.B2(n_217),
.C(n_216),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_513),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_601),
.B(n_227),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_601),
.B(n_252),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_513),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_475),
.B(n_464),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_471),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_531),
.B(n_445),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_598),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_601),
.B(n_254),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_603),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_550),
.B(n_266),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_531),
.B(n_445),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_556),
.B(n_267),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_603),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_477),
.B(n_295),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_608),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_485),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_608),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_611),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_516),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_531),
.B(n_445),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_522),
.B(n_290),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_569),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_496),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_601),
.B(n_303),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_506),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_559),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_516),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_541),
.B(n_314),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_579),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_531),
.B(n_445),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_582),
.B(n_583),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_441),
.Y(n_751)
);

NAND2x1_ASAP7_75t_L g752 ( 
.A(n_525),
.B(n_526),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_611),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_577),
.B(n_441),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_588),
.B(n_441),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

NOR2x2_ASAP7_75t_L g757 ( 
.A(n_512),
.B(n_11),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_594),
.B(n_441),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_586),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_525),
.B(n_315),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_527),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_600),
.B(n_441),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_614),
.B(n_217),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_544),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_485),
.B(n_220),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_544),
.B(n_441),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_546),
.A2(n_586),
.B1(n_612),
.B2(n_578),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_493),
.B(n_510),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_525),
.B(n_441),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_540),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_503),
.B(n_441),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_546),
.A2(n_308),
.B1(n_305),
.B2(n_299),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_514),
.B(n_249),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_485),
.B(n_292),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_503),
.B(n_401),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_527),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_524),
.B(n_292),
.C(n_296),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_589),
.Y(n_779)
);

NOR2x1p5_ASAP7_75t_L g780 ( 
.A(n_512),
.B(n_296),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_528),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_725),
.A2(n_560),
.B(n_565),
.Y(n_782)
);

AO22x1_ASAP7_75t_L g783 ( 
.A1(n_624),
.A2(n_299),
.B1(n_305),
.B2(n_612),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_SL g784 ( 
.A(n_644),
.B(n_512),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_633),
.B(n_485),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_730),
.A2(n_560),
.B(n_565),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_485),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_697),
.B(n_570),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_689),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_748),
.B(n_606),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_739),
.A2(n_560),
.B(n_565),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_749),
.A2(n_526),
.B(n_521),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_713),
.A2(n_526),
.B(n_521),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_741),
.B(n_512),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_695),
.B(n_512),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_695),
.B(n_630),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_657),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_751),
.A2(n_755),
.B(n_754),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_647),
.A2(n_515),
.B(n_571),
.C(n_602),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_634),
.A2(n_642),
.B(n_635),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_764),
.B(n_559),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_735),
.B(n_515),
.Y(n_802)
);

CKINVDCx11_ASAP7_75t_R g803 ( 
.A(n_700),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_684),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_764),
.Y(n_805)
);

AO22x1_ASAP7_75t_L g806 ( 
.A1(n_624),
.A2(n_612),
.B1(n_546),
.B2(n_515),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_662),
.A2(n_515),
.B1(n_589),
.B2(n_562),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_735),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_630),
.B(n_515),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_616),
.B(n_507),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_684),
.Y(n_811)
);

OAI21xp33_ASAP7_75t_SL g812 ( 
.A1(n_737),
.A2(n_548),
.B(n_547),
.Y(n_812)
);

BUFx12f_ASAP7_75t_L g813 ( 
.A(n_724),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_693),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_618),
.B(n_561),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_634),
.A2(n_507),
.B(n_511),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_631),
.A2(n_584),
.B(n_546),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_686),
.B(n_627),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_693),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_659),
.B(n_540),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_723),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_758),
.A2(n_519),
.B(n_511),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_779),
.B(n_729),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_750),
.A2(n_612),
.B1(n_568),
.B2(n_545),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_653),
.B(n_694),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_694),
.B(n_561),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_617),
.B(n_753),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_628),
.B(n_519),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_631),
.A2(n_523),
.B(n_532),
.C(n_553),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_692),
.B(n_520),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_639),
.B(n_523),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_641),
.B(n_532),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_690),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_653),
.B(n_561),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_740),
.B(n_470),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_645),
.B(n_545),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_629),
.B(n_561),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_756),
.A2(n_610),
.B1(n_553),
.B2(n_568),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_762),
.A2(n_555),
.B(n_551),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_654),
.B(n_612),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_638),
.B(n_470),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_620),
.A2(n_555),
.B(n_551),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_646),
.B(n_563),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_759),
.A2(n_563),
.B1(n_552),
.B2(n_604),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_714),
.A2(n_552),
.B(n_543),
.Y(n_847)
);

OAI321xp33_ASAP7_75t_L g848 ( 
.A1(n_733),
.A2(n_678),
.A3(n_716),
.B1(n_660),
.B2(n_691),
.C(n_718),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_640),
.B(n_543),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_620),
.A2(n_538),
.B(n_528),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_649),
.B(n_592),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_643),
.B(n_538),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_674),
.A2(n_564),
.B(n_470),
.C(n_604),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_700),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_663),
.B(n_561),
.C(n_595),
.Y(n_856)
);

O2A1O1Ixp5_ASAP7_75t_L g857 ( 
.A1(n_622),
.A2(n_592),
.B(n_535),
.C(n_604),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_622),
.A2(n_558),
.B(n_478),
.Y(n_858)
);

OAI321xp33_ASAP7_75t_L g859 ( 
.A1(n_716),
.A2(n_12),
.A3(n_15),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_714),
.A2(n_558),
.B(n_478),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_669),
.B(n_558),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_720),
.A2(n_593),
.B(n_596),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_726),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_670),
.B(n_593),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_774),
.B(n_12),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_674),
.A2(n_596),
.B(n_593),
.C(n_535),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_770),
.A2(n_727),
.B(n_721),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_763),
.A2(n_596),
.B(n_535),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_663),
.B(n_595),
.C(n_496),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_752),
.A2(n_595),
.B(n_496),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_667),
.B(n_595),
.C(n_496),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_681),
.B(n_496),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_768),
.B(n_595),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_675),
.B(n_612),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_770),
.A2(n_612),
.B(n_504),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_702),
.B(n_504),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_766),
.A2(n_595),
.B(n_401),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_667),
.B(n_401),
.C(n_504),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_721),
.A2(n_504),
.B(n_609),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_652),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_764),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_750),
.B(n_401),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_728),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_642),
.A2(n_401),
.B(n_504),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_763),
.B(n_504),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_769),
.B(n_401),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_778),
.B(n_401),
.C(n_19),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_738),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_619),
.B(n_18),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_SL g890 ( 
.A1(n_666),
.A2(n_609),
.B(n_22),
.C(n_27),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_666),
.A2(n_609),
.B(n_65),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_699),
.B(n_747),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_21),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_672),
.A2(n_609),
.B(n_66),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_732),
.Y(n_895)
);

AOI21xp33_ASAP7_75t_L g896 ( 
.A1(n_745),
.A2(n_29),
.B(n_30),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_735),
.B(n_32),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_672),
.A2(n_609),
.B(n_72),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_738),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_619),
.Y(n_900)
);

NAND2x1_ASAP7_75t_L g901 ( 
.A(n_746),
.B(n_777),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_704),
.B(n_33),
.C(n_36),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_652),
.B(n_33),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_680),
.A2(n_682),
.B(n_632),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_R g905 ( 
.A(n_618),
.B(n_69),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_651),
.B(n_36),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_764),
.B(n_73),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_765),
.A2(n_775),
.B1(n_651),
.B2(n_655),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_680),
.A2(n_90),
.B(n_143),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_746),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_712),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_655),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_777),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_781),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_712),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_658),
.B(n_37),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_727),
.A2(n_63),
.B(n_136),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_637),
.A2(n_61),
.B1(n_134),
.B2(n_133),
.Y(n_918)
);

O2A1O1Ixp5_ASAP7_75t_L g919 ( 
.A1(n_709),
.A2(n_150),
.B(n_131),
.C(n_124),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_743),
.A2(n_114),
.B(n_106),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_682),
.A2(n_103),
.B(n_100),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_781),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_668),
.A2(n_40),
.B(n_43),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_696),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_765),
.A2(n_775),
.B(n_710),
.C(n_683),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_742),
.A2(n_46),
.B(n_47),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_736),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_621),
.A2(n_48),
.B(n_52),
.Y(n_929)
);

BUFx4_ASAP7_75t_SL g930 ( 
.A(n_757),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_708),
.A2(n_661),
.B(n_780),
.C(n_656),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_SL g932 ( 
.A1(n_743),
.A2(n_52),
.B(n_54),
.C(n_760),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_637),
.A2(n_54),
.B1(n_744),
.B2(n_767),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_623),
.B(n_773),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_665),
.A2(n_673),
.B(n_760),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_767),
.A2(n_773),
.B1(n_650),
.B2(n_771),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_687),
.B(n_688),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_650),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_677),
.B(n_703),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_648),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_679),
.B(n_705),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_685),
.A2(n_707),
.B1(n_711),
.B2(n_698),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_772),
.A2(n_776),
.B(n_626),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_625),
.A2(n_636),
.B(n_664),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_719),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_722),
.A2(n_761),
.B(n_715),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_717),
.B(n_731),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_676),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_717),
.B(n_676),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_676),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_676),
.B(n_671),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_634),
.A2(n_642),
.B(n_635),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_748),
.A2(n_759),
.B1(n_769),
.B2(n_756),
.Y(n_953)
);

NOR2x1_ASAP7_75t_L g954 ( 
.A(n_653),
.B(n_694),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_657),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_653),
.B(n_694),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_735),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_657),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_633),
.A2(n_697),
.B1(n_624),
.B2(n_750),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_657),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_633),
.B(n_613),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_633),
.A2(n_697),
.B1(n_624),
.B2(n_750),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_657),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_633),
.B(n_613),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_961),
.B(n_964),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_796),
.A2(n_809),
.B(n_848),
.Y(n_966)
);

AOI21x1_ASAP7_75t_SL g967 ( 
.A1(n_795),
.A2(n_947),
.B(n_885),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_808),
.Y(n_968)
);

AO31x2_ASAP7_75t_L g969 ( 
.A1(n_830),
.A2(n_926),
.A3(n_936),
.B(n_933),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_888),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_959),
.B(n_962),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_935),
.A2(n_822),
.B(n_841),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_782),
.A2(n_791),
.B(n_786),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_940),
.B(n_828),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_904),
.A2(n_793),
.B(n_857),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_899),
.Y(n_976)
);

AND3x4_ASAP7_75t_L g977 ( 
.A(n_824),
.B(n_956),
.C(n_954),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_782),
.A2(n_791),
.B(n_786),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_904),
.A2(n_793),
.B(n_787),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_943),
.A2(n_844),
.B(n_851),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_844),
.A2(n_851),
.B(n_858),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_941),
.B(n_908),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_866),
.A2(n_952),
.B(n_800),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_818),
.B(n_939),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_860),
.A2(n_862),
.B(n_884),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_948),
.A2(n_785),
.B(n_810),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_808),
.B(n_957),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_939),
.B(n_823),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_784),
.B(n_934),
.Y(n_989)
);

AO21x1_ASAP7_75t_L g990 ( 
.A1(n_917),
.A2(n_920),
.B(n_937),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_799),
.A2(n_790),
.B(n_882),
.Y(n_991)
);

AOI221x1_ASAP7_75t_L g992 ( 
.A1(n_893),
.A2(n_923),
.B1(n_929),
.B2(n_817),
.C(n_794),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_802),
.A2(n_942),
.B1(n_957),
.B2(n_808),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_837),
.B(n_849),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_834),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_948),
.A2(n_792),
.B(n_870),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_805),
.Y(n_997)
);

OAI21x1_ASAP7_75t_SL g998 ( 
.A1(n_909),
.A2(n_921),
.B(n_854),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_802),
.A2(n_957),
.B1(n_808),
.B2(n_912),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_946),
.A2(n_792),
.B(n_847),
.Y(n_1000)
);

BUFx4f_ASAP7_75t_L g1001 ( 
.A(n_813),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_870),
.A2(n_829),
.B(n_868),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_853),
.B(n_820),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_804),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_788),
.B(n_821),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_946),
.A2(n_877),
.B(n_884),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_855),
.B(n_789),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_878),
.A2(n_869),
.B(n_871),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_916),
.B(n_931),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_877),
.A2(n_901),
.B(n_846),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_957),
.Y(n_1011)
);

AO21x2_ASAP7_75t_L g1012 ( 
.A1(n_879),
.A2(n_825),
.B(n_875),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_900),
.B(n_805),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_826),
.B(n_802),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_826),
.B(n_831),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_807),
.B(n_902),
.C(n_892),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_854),
.A2(n_874),
.B(n_852),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_861),
.A2(n_864),
.B(n_845),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_876),
.A2(n_832),
.B(n_833),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_919),
.A2(n_806),
.B(n_953),
.C(n_783),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_911),
.B(n_915),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_812),
.A2(n_949),
.B(n_838),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_865),
.B(n_911),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_811),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_910),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_906),
.B(n_895),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_863),
.B(n_924),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_889),
.A2(n_896),
.B(n_903),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_842),
.B(n_915),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_894),
.A2(n_909),
.B(n_921),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_840),
.A2(n_960),
.B(n_850),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_883),
.B(n_843),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_928),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_911),
.B(n_915),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_913),
.Y(n_1035)
);

OA22x2_ASAP7_75t_L g1036 ( 
.A1(n_897),
.A2(n_880),
.B1(n_859),
.B2(n_930),
.Y(n_1036)
);

INVx6_ASAP7_75t_L g1037 ( 
.A(n_881),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_814),
.B(n_836),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_938),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_872),
.B(n_905),
.Y(n_1040)
);

OAI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_923),
.A2(n_887),
.B(n_801),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_797),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_914),
.A2(n_922),
.B(n_963),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_819),
.A2(n_958),
.B(n_955),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_891),
.A2(n_898),
.B(n_815),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_945),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_907),
.A2(n_929),
.B(n_927),
.C(n_873),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_897),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_891),
.A2(n_898),
.B(n_815),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_897),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_872),
.B(n_881),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_856),
.A2(n_839),
.B(n_827),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_932),
.B(n_886),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_886),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_886),
.B(n_927),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_886),
.B(n_925),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_835),
.A2(n_950),
.B(n_886),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_918),
.B(n_951),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_890),
.A2(n_752),
.B(n_798),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_803),
.A2(n_935),
.B(n_944),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_961),
.B(n_964),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_813),
.Y(n_1062)
);

OAI22x1_ASAP7_75t_L g1063 ( 
.A1(n_823),
.A2(n_570),
.B1(n_741),
.B2(n_468),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_796),
.B(n_427),
.C(n_741),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_961),
.B(n_964),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_796),
.A2(n_926),
.B(n_904),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_798),
.A2(n_752),
.B(n_867),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_805),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_882),
.A2(n_944),
.B(n_935),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_796),
.A2(n_959),
.B(n_962),
.C(n_817),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_796),
.A2(n_959),
.B(n_962),
.C(n_817),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_961),
.B(n_964),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_796),
.A2(n_926),
.B(n_904),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_804),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_888),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_804),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_808),
.B(n_957),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_796),
.A2(n_926),
.B(n_904),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_789),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_798),
.A2(n_752),
.B(n_867),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_888),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_935),
.A2(n_944),
.B(n_822),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_961),
.B(n_964),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_841),
.A2(n_943),
.B(n_816),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_796),
.A2(n_926),
.B(n_904),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_808),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_808),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_813),
.B(n_498),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_841),
.A2(n_943),
.B(n_816),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_789),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_961),
.B(n_964),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_900),
.B(n_809),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_961),
.B(n_964),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_796),
.A2(n_926),
.B(n_904),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_961),
.B(n_964),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_935),
.A2(n_944),
.B(n_822),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_796),
.B(n_729),
.C(n_443),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_796),
.A2(n_431),
.B(n_630),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_SL g1099 ( 
.A1(n_917),
.A2(n_920),
.B(n_909),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_935),
.A2(n_944),
.B(n_822),
.Y(n_1100)
);

BUFx8_ASAP7_75t_SL g1101 ( 
.A(n_813),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_882),
.A2(n_944),
.B(n_935),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_796),
.A2(n_823),
.B1(n_809),
.B2(n_937),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_823),
.A2(n_570),
.B1(n_741),
.B2(n_468),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_808),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_888),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_804),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_796),
.A2(n_790),
.B(n_431),
.C(n_937),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_813),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_SL g1110 ( 
.A(n_1054),
.B(n_968),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1005),
.B(n_1015),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_988),
.B(n_995),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1098),
.B(n_1064),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_970),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_968),
.Y(n_1115)
);

CKINVDCx8_ASAP7_75t_R g1116 ( 
.A(n_1062),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1023),
.B(n_1063),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1014),
.B(n_1021),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1066),
.A2(n_1078),
.B(n_1073),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1085),
.A2(n_1094),
.B(n_1009),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1079),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_989),
.A2(n_1016),
.B1(n_1103),
.B2(n_1097),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_987),
.B(n_1021),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1021),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1023),
.B(n_1104),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_984),
.B(n_1016),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_982),
.A2(n_974),
.B1(n_989),
.B2(n_971),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_965),
.B(n_1061),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1026),
.B(n_1065),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1036),
.A2(n_990),
.B1(n_1028),
.B2(n_966),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1090),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1108),
.B(n_1088),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_987),
.B(n_1048),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1072),
.B(n_1083),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1001),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1014),
.B(n_1039),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_979),
.A2(n_978),
.B(n_973),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1007),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1001),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1070),
.A2(n_1071),
.B1(n_1095),
.B2(n_1093),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_968),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1003),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_976),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1007),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1091),
.B(n_1070),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1025),
.Y(n_1146)
);

AOI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_977),
.A2(n_1036),
.B(n_1014),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1039),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1092),
.B(n_1050),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1071),
.B(n_994),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_986),
.A2(n_1002),
.B(n_1059),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_968),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1035),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1027),
.B(n_1032),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1013),
.B(n_1034),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_SL g1156 ( 
.A(n_1054),
.B(n_1011),
.Y(n_1156)
);

BUFx4f_ASAP7_75t_L g1157 ( 
.A(n_977),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1040),
.A2(n_1029),
.B1(n_1050),
.B2(n_1041),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1029),
.B(n_1033),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1034),
.B(n_1046),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1099),
.A2(n_1022),
.B1(n_991),
.B2(n_998),
.C(n_1020),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1040),
.B(n_1011),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_992),
.B(n_969),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_1011),
.B(n_1086),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_975),
.A2(n_996),
.B(n_1058),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1037),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1062),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_969),
.B(n_1004),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1075),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1077),
.B(n_1086),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1081),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_969),
.B(n_1024),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1109),
.B(n_1101),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_969),
.B(n_1076),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1077),
.B(n_1087),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1087),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1105),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1101),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1105),
.B(n_1051),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1074),
.B(n_1107),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_997),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1056),
.A2(n_1081),
.B1(n_1106),
.B2(n_1058),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_993),
.A2(n_1055),
.B(n_1020),
.C(n_1047),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1105),
.B(n_1068),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1106),
.B(n_1038),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1109),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_1037),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1054),
.A2(n_1000),
.B(n_1031),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1105),
.B(n_997),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1060),
.B(n_1037),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1060),
.B(n_1068),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_999),
.B(n_1053),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1044),
.Y(n_1196)
);

BUFx12f_ASAP7_75t_L g1197 ( 
.A(n_967),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1019),
.B(n_1018),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1012),
.A2(n_1057),
.B1(n_1052),
.B2(n_1008),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1043),
.B(n_1017),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_983),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1012),
.B(n_1006),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_L g1203 ( 
.A(n_967),
.B(n_1047),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_985),
.B(n_972),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_985),
.B(n_1049),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1082),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1069),
.B(n_1102),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1045),
.B(n_1049),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1096),
.A2(n_1100),
.B(n_980),
.Y(n_1210)
);

OAI21xp33_ASAP7_75t_L g1211 ( 
.A1(n_1030),
.A2(n_1045),
.B(n_981),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1010),
.A2(n_1080),
.B(n_1067),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1030),
.A2(n_796),
.B1(n_823),
.B2(n_741),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_970),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1098),
.A2(n_796),
.B(n_1108),
.C(n_431),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_970),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1079),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1062),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_970),
.Y(n_1219)
);

OR2x2_ASAP7_75t_SL g1220 ( 
.A(n_1097),
.B(n_1064),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_974),
.B(n_1098),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1063),
.A2(n_431),
.B1(n_662),
.B2(n_807),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_966),
.A2(n_796),
.B(n_1103),
.Y(n_1223)
);

NAND2x1_ASAP7_75t_L g1224 ( 
.A(n_987),
.B(n_1037),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1021),
.Y(n_1225)
);

CKINVDCx6p67_ASAP7_75t_R g1226 ( 
.A(n_1039),
.Y(n_1226)
);

CKINVDCx8_ASAP7_75t_R g1227 ( 
.A(n_1062),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_974),
.B(n_1098),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_982),
.A2(n_796),
.B1(n_1103),
.B2(n_962),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_988),
.B(n_471),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_970),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1108),
.A2(n_796),
.B(n_1098),
.C(n_1103),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1070),
.A2(n_1071),
.B(n_1066),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_970),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_968),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_987),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_1015),
.Y(n_1237)
);

CKINVDCx16_ASAP7_75t_R g1238 ( 
.A(n_1015),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1098),
.B(n_741),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1005),
.B(n_788),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1014),
.B(n_1021),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_968),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_974),
.B(n_1098),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_987),
.B(n_808),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1098),
.A2(n_427),
.B1(n_1104),
.B2(n_1063),
.C(n_431),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_970),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1098),
.A2(n_431),
.B(n_427),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_974),
.B(n_1098),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1233),
.B(n_1119),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1168),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1222),
.A2(n_1113),
.B1(n_1247),
.B2(n_1245),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1114),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_1134),
.B1(n_1239),
.B2(n_1122),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1157),
.A2(n_1126),
.B1(n_1228),
.B2(n_1243),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1137),
.A2(n_1151),
.B(n_1165),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1190),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1197),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1116),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1167),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1138),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1173),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1175),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1227),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1210),
.A2(n_1191),
.B(n_1212),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1143),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1121),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1117),
.A2(n_1125),
.B1(n_1127),
.B2(n_1229),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1146),
.Y(n_1268)
);

BUFx2_ASAP7_75t_SL g1269 ( 
.A(n_1115),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1201),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1189),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1145),
.B(n_1163),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1201),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1240),
.A2(n_1248),
.B1(n_1221),
.B2(n_1223),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_L g1275 ( 
.A(n_1164),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1144),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1172),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1198),
.A2(n_1205),
.B(n_1120),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1172),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1158),
.A2(n_1220),
.B1(n_1129),
.B2(n_1154),
.Y(n_1280)
);

AND2x4_ASAP7_75t_SL g1281 ( 
.A(n_1226),
.B(n_1136),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1193),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1214),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1142),
.A2(n_1140),
.B1(n_1130),
.B2(n_1111),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1159),
.B(n_1214),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1219),
.B(n_1231),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1219),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1132),
.A2(n_1157),
.B1(n_1150),
.B2(n_1230),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1232),
.A2(n_1215),
.B1(n_1112),
.B2(n_1213),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1234),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1131),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1162),
.B(n_1118),
.Y(n_1292)
);

CKINVDCx14_ASAP7_75t_R g1293 ( 
.A(n_1181),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1153),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1207),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1147),
.A2(n_1237),
.B1(n_1238),
.B2(n_1149),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1164),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1196),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1195),
.A2(n_1186),
.B(n_1185),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1174),
.A2(n_1162),
.B1(n_1139),
.B2(n_1135),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1161),
.A2(n_1160),
.B1(n_1241),
.B2(n_1118),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1202),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1217),
.B(n_1148),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1160),
.A2(n_1155),
.B1(n_1136),
.B2(n_1179),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1199),
.B(n_1208),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1188),
.B(n_1183),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1166),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1169),
.B(n_1216),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1194),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1184),
.A2(n_1155),
.B1(n_1133),
.B2(n_1123),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1182),
.A2(n_1236),
.B1(n_1133),
.B2(n_1124),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1246),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1115),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1156),
.A2(n_1218),
.B1(n_1141),
.B2(n_1152),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1182),
.A2(n_1224),
.B1(n_1236),
.B2(n_1177),
.Y(n_1315)
);

CKINVDCx6p67_ASAP7_75t_R g1316 ( 
.A(n_1141),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1200),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1225),
.B(n_1187),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1200),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1225),
.B(n_1187),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1204),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1206),
.A2(n_1192),
.B1(n_1209),
.B2(n_1211),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1192),
.B(n_1171),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1206),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1178),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1110),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1170),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1171),
.B(n_1176),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1180),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1176),
.A2(n_1177),
.B1(n_1170),
.B2(n_1180),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1180),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1152),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1152),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1235),
.B(n_1242),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1235),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1242),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1242),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1244),
.A2(n_1222),
.B1(n_784),
.B2(n_796),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1168),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1161),
.B(n_796),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1128),
.A2(n_796),
.B1(n_741),
.B2(n_1134),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1168),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1168),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1121),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1121),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1126),
.B(n_1122),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1138),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1126),
.B(n_1122),
.Y(n_1348)
);

AO21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1130),
.A2(n_1223),
.B(n_1009),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1190),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1222),
.A2(n_443),
.B1(n_400),
.B2(n_823),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1114),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1167),
.Y(n_1353)
);

BUFx2_ASAP7_75t_SL g1354 ( 
.A(n_1115),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1121),
.Y(n_1355)
);

BUFx2_ASAP7_75t_SL g1356 ( 
.A(n_1115),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1222),
.A2(n_1098),
.B1(n_1016),
.B2(n_796),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1222),
.A2(n_1098),
.B1(n_1016),
.B2(n_796),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1168),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1128),
.A2(n_796),
.B1(n_741),
.B2(n_1134),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1114),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1168),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1249),
.B(n_1299),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1270),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1297),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1266),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1298),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1278),
.A2(n_1264),
.B(n_1289),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1344),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1345),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1253),
.B(n_1260),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1273),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1334),
.A2(n_1360),
.B(n_1341),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1355),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1297),
.B(n_1275),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1278),
.A2(n_1305),
.B(n_1280),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1282),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1281),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1295),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1346),
.B(n_1348),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1285),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1302),
.B(n_1321),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1281),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1282),
.B(n_1309),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1302),
.B(n_1321),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1309),
.B(n_1250),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1292),
.B(n_1252),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1285),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1261),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1334),
.A2(n_1249),
.B(n_1313),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1262),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1262),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1297),
.B(n_1275),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1339),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1339),
.B(n_1342),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1258),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1283),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1342),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1297),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1343),
.B(n_1359),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1287),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1357),
.B(n_1358),
.C(n_1251),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1362),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1362),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1276),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1317),
.A2(n_1319),
.B(n_1324),
.Y(n_1406)
);

AO21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1267),
.A2(n_1319),
.B(n_1317),
.Y(n_1407)
);

INVxp67_ASAP7_75t_R g1408 ( 
.A(n_1296),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1256),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1324),
.A2(n_1290),
.B(n_1361),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1265),
.A2(n_1268),
.B(n_1361),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1347),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1272),
.B(n_1340),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1275),
.B(n_1340),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1288),
.A2(n_1351),
.B1(n_1254),
.B2(n_1338),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1274),
.B(n_1306),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1284),
.B(n_1340),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1249),
.B(n_1286),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1349),
.B(n_1277),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1327),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1292),
.B(n_1277),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1255),
.A2(n_1310),
.B(n_1327),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1279),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1352),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1292),
.B(n_1318),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1294),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1322),
.A2(n_1301),
.B(n_1312),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1377),
.B(n_1257),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1413),
.B(n_1349),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1371),
.B(n_1291),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1410),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1410),
.Y(n_1432)
);

INVx3_ASAP7_75t_SL g1433 ( 
.A(n_1396),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1402),
.A2(n_1257),
.B1(n_1354),
.B2(n_1269),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1413),
.B(n_1328),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1396),
.Y(n_1436)
);

INVx4_ASAP7_75t_R g1437 ( 
.A(n_1409),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1304),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1406),
.B(n_1308),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1406),
.B(n_1308),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1372),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1382),
.B(n_1385),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1379),
.Y(n_1444)
);

CKINVDCx6p67_ASAP7_75t_R g1445 ( 
.A(n_1409),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1418),
.B(n_1325),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1389),
.B(n_1326),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1380),
.B(n_1331),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1415),
.A2(n_1300),
.B1(n_1307),
.B2(n_1303),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1375),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1417),
.A2(n_1315),
.B1(n_1316),
.B2(n_1307),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1386),
.B(n_1329),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1381),
.B(n_1323),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1416),
.A2(n_1291),
.B1(n_1353),
.B2(n_1271),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_L g1456 ( 
.A(n_1373),
.B(n_1356),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1391),
.B(n_1335),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1411),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1419),
.B(n_1367),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1388),
.B(n_1320),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1419),
.B(n_1364),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1399),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_1423),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1460),
.B(n_1366),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_1405),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1429),
.A2(n_1363),
.B1(n_1414),
.B2(n_1407),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1450),
.A2(n_1414),
.B1(n_1363),
.B2(n_1408),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1454),
.B(n_1369),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1450),
.A2(n_1414),
.B1(n_1363),
.B2(n_1408),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1454),
.B(n_1370),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1456),
.A2(n_1373),
.B(n_1363),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1433),
.B(n_1412),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_L g1474 ( 
.A(n_1455),
.B(n_1256),
.C(n_1350),
.D(n_1395),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1434),
.B(n_1420),
.C(n_1374),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1476)
);

OAI211xp5_ASAP7_75t_L g1477 ( 
.A1(n_1434),
.A2(n_1376),
.B(n_1314),
.C(n_1390),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1443),
.B(n_1391),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1455),
.A2(n_1375),
.B1(n_1393),
.B2(n_1330),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1459),
.B(n_1387),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1452),
.A2(n_1392),
.B1(n_1394),
.B2(n_1398),
.C(n_1403),
.Y(n_1482)
);

OAI221xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1452),
.A2(n_1390),
.B1(n_1293),
.B2(n_1311),
.C(n_1395),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1403),
.C(n_1394),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1433),
.B(n_1425),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1428),
.B(n_1392),
.C(n_1404),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1433),
.B(n_1387),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1429),
.A2(n_1393),
.B(n_1375),
.Y(n_1488)
);

NOR3xp33_ASAP7_75t_L g1489 ( 
.A(n_1457),
.B(n_1368),
.C(n_1365),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1457),
.B(n_1426),
.C(n_1427),
.Y(n_1491)
);

NAND2xp33_ASAP7_75t_SL g1492 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1421),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1438),
.C(n_1447),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1435),
.B(n_1400),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1463),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1446),
.B(n_1424),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1437),
.A2(n_1393),
.B1(n_1353),
.B2(n_1271),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1445),
.A2(n_1378),
.B1(n_1383),
.B2(n_1337),
.Y(n_1499)
);

NAND4xp25_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1350),
.C(n_1397),
.D(n_1401),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1438),
.A2(n_1407),
.B1(n_1421),
.B2(n_1425),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1451),
.B(n_1425),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1476),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1490),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1490),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1496),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1478),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1479),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1479),
.B(n_1494),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1468),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1481),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1484),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1493),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1491),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1497),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1472),
.B(n_1462),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1464),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1471),
.B(n_1458),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1502),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1487),
.Y(n_1527)
);

AND2x4_ASAP7_75t_SL g1528 ( 
.A(n_1466),
.B(n_1365),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1442),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1488),
.B(n_1432),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1514),
.B(n_1446),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1518),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1530),
.B(n_1516),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1440),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1506),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1526),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1440),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1507),
.B(n_1500),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1521),
.Y(n_1549)
);

INVxp33_ASAP7_75t_L g1550 ( 
.A(n_1523),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1515),
.B(n_1441),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1526),
.Y(n_1553)
);

NOR2x1p5_ASAP7_75t_SL g1554 ( 
.A(n_1512),
.B(n_1432),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1516),
.B(n_1453),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1517),
.A2(n_1475),
.B(n_1474),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1448),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1518),
.A2(n_1483),
.B1(n_1475),
.B2(n_1467),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1521),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1523),
.A2(n_1470),
.B1(n_1477),
.B2(n_1492),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1525),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1525),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1530),
.B(n_1444),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1526),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1533),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1549),
.B(n_1551),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1559),
.B(n_1498),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1565),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1534),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1537),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1526),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1577)
);

INVxp33_ASAP7_75t_L g1578 ( 
.A(n_1541),
.Y(n_1578)
);

OAI32xp33_ASAP7_75t_L g1579 ( 
.A1(n_1557),
.A2(n_1517),
.A3(n_1511),
.B1(n_1510),
.B2(n_1512),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1551),
.B(n_1517),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1540),
.B(n_1511),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1547),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1522),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1539),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1565),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1538),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1522),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1539),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1540),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1565),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1538),
.B(n_1530),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1543),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1538),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1536),
.B(n_1516),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1532),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1522),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1536),
.B(n_1516),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1562),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1565),
.B(n_1522),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1543),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1556),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1556),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1547),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1516),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1560),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_1604),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1554),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

AND3x1_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1465),
.C(n_1527),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1571),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1604),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1604),
.A2(n_1570),
.B1(n_1600),
.B2(n_1578),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1567),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1569),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1259),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1570),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1560),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1595),
.B(n_1561),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1569),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1566),
.B(n_1563),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1579),
.B(n_1563),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1577),
.B(n_1542),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1545),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1561),
.Y(n_1628)
);

CKINVDCx14_ASAP7_75t_R g1629 ( 
.A(n_1570),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1572),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1564),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1570),
.B(n_1531),
.Y(n_1633)
);

AOI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1582),
.A2(n_1529),
.B1(n_1554),
.B2(n_1520),
.C1(n_1528),
.C2(n_1498),
.Y(n_1634)
);

INVx4_ASAP7_75t_L g1635 ( 
.A(n_1608),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1572),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1529),
.C(n_1545),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1574),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1581),
.B(n_1259),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1574),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1573),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1575),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1573),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1611),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1587),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_R g1648 ( 
.A1(n_1619),
.A2(n_1580),
.B1(n_1568),
.B2(n_1603),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1620),
.B(n_1259),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1615),
.A2(n_1568),
.B(n_1580),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1633),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1612),
.B(n_1605),
.C(n_1603),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1629),
.A2(n_1593),
.B(n_1601),
.Y(n_1653)
);

XNOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1632),
.B(n_1492),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1625),
.A2(n_1605),
.B1(n_1591),
.B2(n_1594),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1628),
.A2(n_1528),
.B1(n_1596),
.B2(n_1599),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1632),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1622),
.Y(n_1660)
);

AOI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1634),
.A2(n_1592),
.B(n_1591),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1637),
.A2(n_1602),
.B(n_1594),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1639),
.B(n_1635),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1611),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1665)
);

AOI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1613),
.A2(n_1592),
.B(n_1602),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1621),
.A2(n_1499),
.B(n_1512),
.C(n_1480),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1635),
.A2(n_1528),
.B1(n_1599),
.B2(n_1596),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1635),
.A2(n_1528),
.B1(n_1527),
.B2(n_1445),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1651),
.B(n_1613),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1659),
.B(n_1626),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1646),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1660),
.B(n_1626),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1645),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1663),
.B(n_1610),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1654),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1655),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1644),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1644),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1622),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1663),
.B(n_1631),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1664),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1662),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1631),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1656),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1653),
.B(n_1627),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1610),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1648),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1672),
.B(n_1681),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1685),
.B(n_1661),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1683),
.A2(n_1657),
.B1(n_1652),
.B2(n_1666),
.C(n_1658),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1688),
.A2(n_1668),
.B1(n_1669),
.B2(n_1667),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1670),
.B(n_1686),
.C(n_1679),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1677),
.A2(n_1638),
.B(n_1616),
.C(n_1630),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1684),
.A2(n_1636),
.B(n_1623),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1686),
.A2(n_1610),
.B(n_1665),
.C(n_1627),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1643),
.C(n_1641),
.D(n_1642),
.Y(n_1697)
);

NAND4xp75_ASAP7_75t_L g1698 ( 
.A(n_1681),
.B(n_1643),
.C(n_1641),
.D(n_1642),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1685),
.A2(n_1640),
.B(n_1617),
.Y(n_1699)
);

NAND4xp25_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1640),
.C(n_1617),
.D(n_1589),
.Y(n_1700)
);

XNOR2xp5_ASAP7_75t_L g1701 ( 
.A(n_1692),
.B(n_1678),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_L g1702 ( 
.A(n_1690),
.B(n_1680),
.C(n_1678),
.D(n_1671),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1689),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1694),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1691),
.B(n_1673),
.C(n_1682),
.D(n_1674),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1697),
.B(n_1675),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1700),
.B(n_1687),
.Y(n_1709)
);

NOR4xp25_ASAP7_75t_L g1710 ( 
.A(n_1699),
.B(n_1687),
.C(n_1585),
.D(n_1590),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1703),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1705),
.A2(n_1710),
.B(n_1708),
.C(n_1706),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1701),
.B(n_1696),
.Y(n_1713)
);

NOR4xp25_ASAP7_75t_L g1714 ( 
.A(n_1704),
.B(n_1695),
.C(n_1575),
.D(n_1590),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1707),
.A2(n_1263),
.B(n_1337),
.C(n_1584),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1711),
.B(n_1709),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1712),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1713),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1715),
.B(n_1702),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1714),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1711),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1716),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1717),
.A2(n_1583),
.B1(n_1586),
.B2(n_1585),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1716),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1721),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1720),
.B(n_1583),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1722),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1724),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1725),
.B(n_1719),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1727),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1728),
.B(n_1718),
.C(n_1729),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1726),
.B(n_1723),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1731),
.Y(n_1733)
);

AOI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1726),
.B(n_1586),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1732),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1583),
.B(n_1606),
.Y(n_1736)
);

NAND2x1_ASAP7_75t_L g1737 ( 
.A(n_1734),
.B(n_1606),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1736),
.A2(n_1607),
.B(n_1513),
.Y(n_1738)
);

AOI322xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1737),
.A3(n_1607),
.B1(n_1503),
.B2(n_1520),
.C1(n_1548),
.C2(n_1552),
.Y(n_1739)
);

OAI221xp5_ASAP7_75t_R g1740 ( 
.A1(n_1739),
.A2(n_1316),
.B1(n_1501),
.B2(n_1437),
.C(n_1445),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1332),
.B(n_1333),
.C(n_1336),
.Y(n_1741)
);


endmodule