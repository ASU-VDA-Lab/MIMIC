module fake_jpeg_6510_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_49),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_26),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_55),
.C(n_87),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_58),
.Y(n_111)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_59),
.B(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_19),
.B1(n_16),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_76),
.B1(n_89),
.B2(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_66),
.Y(n_122)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_79),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_78),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_28),
.B1(n_32),
.B2(n_22),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_95),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_37),
.A2(n_35),
.B1(n_18),
.B2(n_14),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_39),
.A2(n_35),
.B1(n_18),
.B2(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_36),
.B(n_13),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_12),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_12),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_40),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_27),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_109),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_0),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_108),
.B(n_15),
.Y(n_165)
);

OR2x4_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_118),
.B(n_133),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_133),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_54),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_73),
.A2(n_30),
.B1(n_25),
.B2(n_15),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_80),
.B1(n_64),
.B2(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_141),
.A2(n_24),
.B1(n_128),
.B2(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_70),
.C(n_71),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_103),
.C(n_27),
.Y(n_192)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_94),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_31),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_82),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_151),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_76),
.A3(n_100),
.B1(n_63),
.B2(n_82),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_155),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_101),
.C(n_68),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_167),
.C(n_113),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_68),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_104),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_160),
.B1(n_121),
.B2(n_105),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_106),
.A2(n_83),
.B1(n_61),
.B2(n_92),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_166),
.B1(n_168),
.B2(n_117),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_75),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_169),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_107),
.A2(n_92),
.B(n_97),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_165),
.B(n_119),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_83),
.B1(n_84),
.B2(n_58),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_84),
.A3(n_15),
.B1(n_25),
.B2(n_30),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_105),
.A2(n_35),
.B1(n_18),
.B2(n_25),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_103),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_185),
.B1(n_141),
.B2(n_136),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_198),
.C(n_200),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_183),
.B(n_167),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_118),
.B(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_116),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_116),
.B1(n_115),
.B2(n_121),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_115),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_196),
.C(n_204),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_134),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_197),
.Y(n_209)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_103),
.C(n_31),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_27),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_27),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_207),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_156),
.B1(n_140),
.B2(n_142),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_24),
.C(n_1),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_0),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_193),
.Y(n_255)
);

AOI221xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_172),
.B1(n_178),
.B2(n_196),
.C(n_207),
.Y(n_241)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_166),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_226),
.B(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

NOR2x1_ASAP7_75t_R g220 ( 
.A(n_183),
.B(n_181),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_202),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_173),
.A2(n_162),
.B1(n_138),
.B2(n_151),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_227),
.B1(n_185),
.B2(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_149),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_231),
.Y(n_246)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_172),
.A2(n_168),
.B(n_146),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_0),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_2),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_24),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_249),
.B1(n_186),
.B2(n_190),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_255),
.Y(n_271)
);

OAI321xp33_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_212),
.A3(n_220),
.B1(n_226),
.B2(n_211),
.C(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_253),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_192),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_250),
.C(n_251),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_216),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_179),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_258),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_214),
.B(n_203),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_223),
.C(n_213),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_217),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_210),
.B(n_187),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_215),
.B1(n_222),
.B2(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_227),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_244),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_219),
.B1(n_234),
.B2(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_269),
.C(n_246),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_210),
.B1(n_190),
.B2(n_199),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_275),
.B(n_242),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_270),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_199),
.B(n_182),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_257),
.B(n_244),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_224),
.C(n_206),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_191),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_273)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_197),
.B1(n_24),
.B2(n_2),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_255),
.C(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_277),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_246),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.C(n_266),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_262),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_284),
.B(n_288),
.Y(n_294)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_275),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_254),
.C(n_256),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_254),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_283),
.B1(n_286),
.B2(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_279),
.C(n_271),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_301),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_280),
.B(n_269),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_299),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_264),
.B(n_262),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_300),
.B(n_294),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_297),
.A2(n_282),
.B1(n_273),
.B2(n_287),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_259),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_278),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_304),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_279),
.C(n_261),
.Y(n_310)
);

AOI221xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_307),
.C(n_4),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_265),
.B(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_4),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_306),
.B(n_310),
.C(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_4),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.C(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_5),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_319),
.Y(n_321)
);


endmodule