module fake_jpeg_25236_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_29),
.B1(n_18),
.B2(n_24),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_42),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_18),
.B1(n_24),
.B2(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_53),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_33),
.Y(n_50)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_22),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_59),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_35),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_30),
.B1(n_25),
.B2(n_20),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_23),
.B1(n_27),
.B2(n_21),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_31),
.B1(n_32),
.B2(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_37),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_16),
.B(n_34),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_37),
.B1(n_18),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_17),
.B1(n_34),
.B2(n_15),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_23),
.Y(n_91)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_93),
.B1(n_104),
.B2(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_44),
.C(n_40),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_72),
.C(n_61),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_46),
.B1(n_32),
.B2(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_92),
.B1(n_77),
.B2(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_86),
.B(n_90),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_16),
.B(n_1),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_99),
.B(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_77),
.B1(n_60),
.B2(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_79),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_16),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_72),
.B1(n_78),
.B2(n_30),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_20),
.CON(n_103),
.SN(n_103)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_105),
.B1(n_21),
.B2(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_30),
.B1(n_25),
.B2(n_34),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_117),
.B1(n_123),
.B2(n_124),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_77),
.B(n_55),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_133),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_118),
.Y(n_144)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_126),
.B1(n_15),
.B2(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_135),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_72),
.B1(n_75),
.B2(n_57),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_107),
.B1(n_84),
.B2(n_27),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_80),
.B1(n_73),
.B2(n_69),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_65),
.B1(n_58),
.B2(n_68),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_65),
.B1(n_68),
.B2(n_15),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_101),
.B1(n_83),
.B2(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_58),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_138),
.A2(n_139),
.B(n_146),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_87),
.B(n_101),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_81),
.B1(n_82),
.B2(n_104),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_99),
.B(n_101),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_129),
.B(n_121),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_148),
.B(n_3),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_92),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_134),
.B1(n_119),
.B2(n_130),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_100),
.B(n_91),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_118),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_100),
.B1(n_102),
.B2(n_97),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_90),
.B1(n_107),
.B2(n_83),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_160),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_88),
.C(n_86),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_158),
.C(n_115),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_15),
.C(n_21),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_23),
.B1(n_15),
.B2(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_165),
.B1(n_112),
.B2(n_117),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_0),
.B(n_2),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_166),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_189),
.B1(n_195),
.B2(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_190),
.Y(n_198)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_177),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_194),
.C(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_145),
.B1(n_153),
.B2(n_151),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_128),
.A3(n_131),
.B1(n_112),
.B2(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_186),
.A2(n_147),
.B1(n_160),
.B2(n_166),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_8),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_136),
.B(n_9),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_10),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_4),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_196),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_171),
.B1(n_182),
.B2(n_181),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_150),
.B1(n_154),
.B2(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_209),
.B1(n_173),
.B2(n_188),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_218),
.C(n_185),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_149),
.B1(n_147),
.B2(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_214),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_137),
.C(n_146),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_172),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_185),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_229),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_235),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_171),
.B1(n_186),
.B2(n_145),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_173),
.B(n_167),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_194),
.C(n_179),
.Y(n_236)
);

XNOR2x2_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_180),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_239),
.A2(n_219),
.B1(n_197),
.B2(n_217),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_197),
.CI(n_211),
.CON(n_243),
.SN(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_201),
.B1(n_202),
.B2(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_249),
.B1(n_215),
.B2(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_237),
.C(n_220),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.C(n_260),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_258),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_183),
.B1(n_243),
.B2(n_240),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_224),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_4),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_236),
.C(n_230),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_200),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_264),
.B1(n_158),
.B2(n_5),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_222),
.C(n_208),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_208),
.C(n_210),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_143),
.B1(n_184),
.B2(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_235),
.B1(n_152),
.B2(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_174),
.B1(n_189),
.B2(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_270),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_247),
.B(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.C(n_274),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_138),
.B(n_139),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_253),
.B1(n_6),
.B2(n_7),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_5),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_274),
.C(n_270),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_279),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_6),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_278),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_286),
.B(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_288),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_269),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_5),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_287),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_6),
.A3(n_7),
.B1(n_280),
.B2(n_291),
.C(n_293),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_6),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);


endmodule