module fake_jpeg_3606_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_49),
.B1(n_46),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_62),
.B1(n_39),
.B2(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_49),
.B1(n_46),
.B2(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_41),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_39),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_47),
.C(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_66),
.C(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_61),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_42),
.B(n_65),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_1),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_63),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_73),
.B(n_79),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_74),
.C(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_109),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_89),
.C(n_81),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_64),
.B1(n_42),
.B2(n_35),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_34),
.C(n_33),
.D(n_32),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_19),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_64),
.B(n_2),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_92),
.B(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_106),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_3),
.B(n_4),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_102),
.B(n_100),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_117),
.C(n_13),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_20),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_5),
.B(n_7),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_131),
.C(n_117),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_95),
.B(n_10),
.C(n_12),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

OAI22x1_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_125),
.B1(n_124),
.B2(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.C(n_14),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_112),
.A3(n_114),
.B1(n_120),
.B2(n_122),
.C(n_16),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_127),
.B1(n_130),
.B2(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_128),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_136),
.B1(n_132),
.B2(n_17),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_14),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_141),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_140),
.B(n_16),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_17),
.Y(n_146)
);


endmodule