module fake_jpeg_4526_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_23),
.B(n_25),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_17),
.Y(n_72)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_30),
.B1(n_20),
.B2(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_22),
.B(n_24),
.Y(n_115)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_77),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_23),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_31),
.B1(n_24),
.B2(n_33),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_49),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_28),
.B1(n_36),
.B2(n_26),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_66),
.B1(n_69),
.B2(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_116),
.B1(n_120),
.B2(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_88),
.C(n_99),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_105),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_40),
.C(n_39),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_69),
.B1(n_31),
.B2(n_73),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_95),
.B1(n_82),
.B2(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_47),
.C(n_44),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_122),
.B(n_27),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_86),
.B(n_25),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_21),
.B1(n_18),
.B2(n_22),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_21),
.B1(n_18),
.B2(n_28),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_40),
.C(n_44),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_28),
.B1(n_26),
.B2(n_36),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_74),
.A2(n_28),
.B1(n_26),
.B2(n_36),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_120),
.B1(n_83),
.B2(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_25),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_144),
.B1(n_157),
.B2(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_149),
.B1(n_153),
.B2(n_156),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_14),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_79),
.B1(n_50),
.B2(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_25),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_149),
.B1(n_155),
.B2(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_124),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_152),
.B(n_154),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_47),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_114),
.B1(n_105),
.B2(n_106),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_156),
.B1(n_100),
.B2(n_111),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_86),
.B(n_25),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_59),
.B1(n_58),
.B2(n_36),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_50),
.B1(n_59),
.B2(n_27),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_111),
.C(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_178),
.C(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_166),
.B(n_176),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_158),
.B(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_100),
.B1(n_128),
.B2(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_126),
.B1(n_117),
.B2(n_113),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_158),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_117),
.B1(n_113),
.B2(n_94),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_27),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_188),
.B1(n_185),
.B2(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_184),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_185),
.B(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_0),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_189),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_209),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_139),
.B(n_142),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_202),
.C(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_148),
.C(n_155),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_10),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_2),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_206),
.B(n_12),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_2),
.B(n_3),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_222),
.B(n_190),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_216),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_219),
.B1(n_221),
.B2(n_167),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_177),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_220),
.B1(n_188),
.B2(n_171),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_169),
.A2(n_4),
.B(n_6),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_205),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_241),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_166),
.B1(n_163),
.B2(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_180),
.B1(n_189),
.B2(n_161),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_238),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_169),
.B(n_192),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_186),
.C(n_173),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_244),
.C(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_186),
.C(n_159),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_218),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_209),
.B1(n_195),
.B2(n_203),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_206),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_199),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_222),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.C(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_204),
.C(n_194),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_213),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_229),
.B(n_242),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_244),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_233),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_225),
.B(n_226),
.Y(n_280)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_257),
.C(n_258),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_241),
.C(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_275),
.C(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_236),
.C(n_227),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_246),
.B1(n_238),
.B2(n_223),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_279),
.B1(n_263),
.B2(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_232),
.B1(n_229),
.B2(n_224),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_285),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_228),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_283),
.B(n_255),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_195),
.C(n_245),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_249),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_260),
.Y(n_290)
);

OAI221xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_259),
.B1(n_265),
.B2(n_250),
.C(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_277),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_278),
.B1(n_247),
.B2(n_218),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_297),
.C(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_265),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_270),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_262),
.C(n_264),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_268),
.C(n_243),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_302),
.C(n_200),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_212),
.C(n_261),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_305),
.B(n_309),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_280),
.B(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_271),
.B(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_299),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_213),
.B(n_248),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.C(n_292),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_214),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_16),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_16),
.C(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_304),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_16),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_313),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_327),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_331),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_324),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_316),
.B(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_319),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_330),
.C(n_334),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_303),
.C(n_307),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_332),
.B(n_311),
.Y(n_340)
);


endmodule