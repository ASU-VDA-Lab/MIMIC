module fake_jpeg_13559_n_364 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_364);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_364;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_58),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_8),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_60),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_9),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_79),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_71),
.Y(n_124)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_83),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_73),
.A2(n_75),
.B1(n_88),
.B2(n_82),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_6),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_76),
.B(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_48),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_9),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_13),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_13),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_86),
.Y(n_138)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_16),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_92),
.Y(n_153)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_32),
.B(n_13),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_15),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_33),
.B(n_0),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_99),
.Y(n_122)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_97),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_35),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_101),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_36),
.B1(n_23),
.B2(n_43),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_103),
.A2(n_112),
.B1(n_121),
.B2(n_127),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_51),
.B1(n_44),
.B2(n_43),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_104),
.A2(n_105),
.B1(n_157),
.B2(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_51),
.B1(n_44),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_122),
.B1(n_110),
.B2(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_111),
.B(n_116),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_55),
.A2(n_36),
.B1(n_25),
.B2(n_40),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_117),
.A2(n_149),
.B1(n_62),
.B2(n_64),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_133),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_61),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_127)
);

AND2x4_ASAP7_75t_SL g129 ( 
.A(n_78),
.B(n_1),
.Y(n_129)
);

OR2x2_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_80),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_107),
.Y(n_190)
);

CKINVDCx12_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx12_ASAP7_75t_R g141 ( 
.A(n_95),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_74),
.A2(n_49),
.B1(n_85),
.B2(n_100),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_74),
.B1(n_146),
.B2(n_135),
.Y(n_189)
);

CKINVDCx12_ASAP7_75t_R g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_59),
.B(n_70),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_67),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_160),
.A2(n_182),
.B1(n_205),
.B2(n_126),
.Y(n_237)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_69),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_191),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_178),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_168),
.B(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

OR2x2_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_122),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_206),
.B(n_207),
.Y(n_233)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_176),
.Y(n_243)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_56),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_128),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_185),
.Y(n_212)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_109),
.B(n_58),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_190),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_188),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_146),
.B1(n_135),
.B2(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_108),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_196),
.Y(n_230)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_198),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_200),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_153),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_132),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_131),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_179),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_104),
.B1(n_129),
.B2(n_155),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_216),
.B1(n_220),
.B2(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_247),
.B1(n_167),
.B2(n_201),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_163),
.A2(n_104),
.B1(n_113),
.B2(n_150),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_119),
.B1(n_125),
.B2(n_150),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_154),
.B1(n_120),
.B2(n_139),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_161),
.Y(n_274)
);

OR2x2_ASAP7_75t_SL g256 ( 
.A(n_228),
.B(n_200),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_239),
.B(n_177),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_160),
.A2(n_125),
.B1(n_119),
.B2(n_154),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_183),
.B1(n_192),
.B2(n_194),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_170),
.A2(n_115),
.B(n_139),
.C(n_131),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_145),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_165),
.A2(n_115),
.B1(n_172),
.B2(n_205),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_168),
.B1(n_171),
.B2(n_174),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_176),
.B(n_188),
.CI(n_166),
.CON(n_248),
.SN(n_248)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_195),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_224),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_251),
.A2(n_256),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_187),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_262),
.C(n_228),
.Y(n_277)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_203),
.C(n_195),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_212),
.B(n_187),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_173),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_211),
.B1(n_228),
.B2(n_216),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_274),
.B(n_276),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_209),
.B(n_196),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_269),
.B(n_239),
.Y(n_282)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_252),
.B1(n_237),
.B2(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_270),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_221),
.A2(n_203),
.B(n_195),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_180),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_236),
.B1(n_243),
.B2(n_222),
.Y(n_288)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_164),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_292),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_279),
.A2(n_273),
.B1(n_250),
.B2(n_266),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_240),
.B(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_290),
.Y(n_304)
);

AOI221xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_221),
.B1(n_217),
.B2(n_241),
.C(n_242),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_258),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_289),
.B1(n_252),
.B2(n_268),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_222),
.B1(n_241),
.B2(n_248),
.Y(n_289)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_230),
.A3(n_210),
.B1(n_222),
.B2(n_246),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_249),
.A2(n_218),
.A3(n_243),
.B1(n_214),
.B2(n_227),
.C1(n_215),
.C2(n_232),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_269),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_215),
.B(n_227),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_214),
.B(n_259),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_302),
.A2(n_307),
.B1(n_283),
.B2(n_282),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_251),
.B1(n_254),
.B2(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_305),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_255),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_315),
.Y(n_319)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_232),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_293),
.B(n_275),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_284),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_303),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_323),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_292),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_308),
.C(n_297),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_304),
.A2(n_279),
.A3(n_287),
.B1(n_297),
.B2(n_291),
.C(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_329),
.B(n_335),
.Y(n_343)
);

NOR4xp25_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_291),
.C(n_300),
.D(n_304),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_336),
.C(n_280),
.Y(n_340)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_333),
.Y(n_346)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_324),
.C(n_319),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_295),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_286),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_321),
.Y(n_337)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_337),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_327),
.A2(n_309),
.B(n_319),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_338),
.A2(n_327),
.B1(n_318),
.B2(n_307),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_340),
.A2(n_347),
.B1(n_335),
.B2(n_312),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_323),
.C(n_318),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_286),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_339),
.A2(n_288),
.B1(n_321),
.B2(n_290),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_345),
.A2(n_331),
.B(n_339),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_349),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_341),
.A2(n_338),
.B(n_335),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_351),
.Y(n_355)
);

AOI322xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_310),
.A3(n_306),
.B1(n_301),
.B2(n_285),
.C1(n_296),
.C2(n_294),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_342),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_356),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_353),
.A2(n_343),
.B1(n_344),
.B2(n_296),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_343),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_358),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_356),
.A2(n_344),
.B1(n_278),
.B2(n_346),
.Y(n_360)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_360),
.A2(n_298),
.A3(n_351),
.B1(n_354),
.B2(n_355),
.C1(n_357),
.C2(n_359),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_362),
.B(n_326),
.CI(n_304),
.CON(n_363),
.SN(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_361),
.Y(n_364)
);


endmodule