module fake_jpeg_7466_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_33),
.B1(n_20),
.B2(n_32),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_57),
.B1(n_63),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_33),
.B1(n_20),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_52),
.B1(n_30),
.B2(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_33),
.B1(n_19),
.B2(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_54),
.Y(n_77)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_20),
.B1(n_22),
.B2(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_32),
.B1(n_22),
.B2(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_76),
.B1(n_83),
.B2(n_89),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_16),
.C(n_29),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_84),
.C(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_30),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_88),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_16),
.C(n_29),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_32),
.B1(n_24),
.B2(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_112),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_13),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_48),
.B1(n_24),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_77),
.B1(n_86),
.B2(n_43),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_48),
.B1(n_62),
.B2(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_18),
.B(n_27),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_106),
.B(n_107),
.C(n_27),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_70),
.B(n_90),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_27),
.B(n_18),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_72),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_59),
.C(n_46),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_116),
.C(n_85),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_18),
.B(n_27),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_64),
.B(n_51),
.C(n_31),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_24),
.B1(n_34),
.B2(n_51),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_43),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_54),
.B1(n_17),
.B2(n_25),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_36),
.C(n_40),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_54),
.B1(n_17),
.B2(n_25),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_88),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_129),
.C(n_144),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_127),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_91),
.B1(n_74),
.B2(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_133),
.B1(n_147),
.B2(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_131),
.Y(n_153)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_107),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_86),
.B1(n_72),
.B2(n_43),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_136),
.B(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_140),
.B1(n_108),
.B2(n_113),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_26),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_10),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_77),
.B1(n_40),
.B2(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_95),
.C(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_10),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_23),
.B1(n_66),
.B2(n_77),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_157),
.B1(n_163),
.B2(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_97),
.B1(n_107),
.B2(n_108),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_106),
.B1(n_100),
.B2(n_116),
.Y(n_160)
);

AOI22x1_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_101),
.B1(n_23),
.B2(n_27),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_67),
.B1(n_115),
.B2(n_2),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_67),
.B1(n_115),
.B2(n_2),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_137),
.B1(n_130),
.B2(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_115),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_172),
.B1(n_145),
.B2(n_127),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_7),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_120),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.C(n_191),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_129),
.C(n_132),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_188),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_132),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_192),
.B(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_198),
.B1(n_177),
.B2(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_122),
.C(n_5),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_4),
.C(n_5),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_203),
.C(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_196),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_204),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_214),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_155),
.B1(n_150),
.B2(n_157),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_185),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_155),
.B1(n_161),
.B2(n_169),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_171),
.B1(n_160),
.B2(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_225),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_181),
.B(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_182),
.C(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_183),
.B(n_189),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_227),
.B(n_229),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_189),
.A2(n_151),
.B(n_149),
.C(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_241),
.B1(n_213),
.B2(n_222),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_179),
.B(n_203),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_244),
.B(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_208),
.C(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_149),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_151),
.B1(n_176),
.B2(n_148),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_205),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_224),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_216),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_231),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_208),
.C(n_210),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_206),
.C(n_217),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_214),
.C(n_227),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_262),
.B(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_220),
.C(n_224),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_248),
.B1(n_249),
.B2(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_256),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_273),
.B(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_239),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_246),
.B(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_240),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_246),
.B1(n_231),
.B2(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_261),
.C(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_252),
.C(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_266),
.C(n_278),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_286),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_264),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_293),
.B(n_9),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_264),
.B(n_234),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_8),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_286),
.B1(n_251),
.B2(n_10),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_191),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_8),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_304),
.B1(n_297),
.B2(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_11),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_306),
.Y(n_309)
);

OAI221xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_305),
.B1(n_298),
.B2(n_13),
.C(n_14),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_11),
.A3(n_12),
.B(n_14),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_11),
.Y(n_312)
);


endmodule