module fake_jpeg_13837_n_499 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_499);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_499;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_0),
.B(n_14),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_53),
.B(n_63),
.Y(n_147)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_97),
.Y(n_120)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_15),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_24),
.B1(n_23),
.B2(n_27),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_102),
.A2(n_84),
.B1(n_76),
.B2(n_79),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_43),
.B1(n_27),
.B2(n_23),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_133),
.B1(n_141),
.B2(n_26),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_52),
.B(n_50),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_135),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_27),
.B1(n_40),
.B2(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_50),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_20),
.B1(n_29),
.B2(n_40),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_144),
.B1(n_26),
.B2(n_21),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_78),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_17),
.B1(n_33),
.B2(n_37),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_21),
.B1(n_47),
.B2(n_37),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_17),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_149),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_70),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_34),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_156),
.B(n_167),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_96),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_165),
.C(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_160),
.Y(n_245)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_163),
.A2(n_180),
.B1(n_202),
.B2(n_45),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_95),
.C(n_94),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_34),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_47),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_173),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_47),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_181),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_103),
.B(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_37),
.B(n_22),
.C(n_21),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_186),
.A2(n_36),
.B(n_48),
.C(n_45),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_26),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_154),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_155),
.B1(n_85),
.B2(n_83),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_22),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_198),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g198 ( 
.A(n_153),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_146),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_108),
.A2(n_57),
.B1(n_71),
.B2(n_54),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_104),
.A2(n_56),
.B1(n_82),
.B2(n_90),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_115),
.B(n_152),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_111),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_105),
.B(n_22),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_32),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_36),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_131),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_211),
.B(n_193),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_163),
.A2(n_102),
.B1(n_87),
.B2(n_73),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_217),
.A2(n_155),
.B1(n_110),
.B2(n_152),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_168),
.Y(n_267)
);

AOI32xp33_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_108),
.A3(n_136),
.B1(n_150),
.B2(n_92),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_219),
.A2(n_203),
.B(n_185),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_226),
.B(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_148),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_244),
.Y(n_255)
);

OA22x2_ASAP7_75t_SL g230 ( 
.A1(n_165),
.A2(n_136),
.B1(n_110),
.B2(n_148),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_243),
.B(n_186),
.C(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_237),
.A2(n_126),
.B1(n_196),
.B2(n_189),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_146),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_246),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_250),
.A2(n_262),
.B(n_215),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_180),
.B(n_157),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_251),
.A2(n_258),
.B(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_275),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_217),
.A2(n_166),
.B1(n_177),
.B2(n_197),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_202),
.B(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_159),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_265),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_261),
.B(n_267),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_221),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_182),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_212),
.B(n_190),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_273),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_277),
.B1(n_242),
.B2(n_241),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_191),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_272),
.B(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_212),
.B(n_192),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_175),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_278),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_276),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_111),
.B1(n_199),
.B2(n_126),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_287),
.B1(n_228),
.B2(n_241),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_227),
.B(n_201),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_215),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_209),
.B(n_183),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_208),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.C(n_229),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_208),
.B(n_164),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_230),
.A2(n_67),
.B1(n_93),
.B2(n_88),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_230),
.A2(n_164),
.B(n_198),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_299),
.B1(n_305),
.B2(n_310),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_255),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_252),
.A2(n_230),
.B1(n_228),
.B2(n_243),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_296),
.B1(n_317),
.B2(n_271),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_267),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_221),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_307),
.C(n_309),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_312),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_251),
.B1(n_250),
.B2(n_253),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_250),
.A2(n_242),
.B1(n_223),
.B2(n_213),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_235),
.C(n_240),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_235),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_213),
.B1(n_223),
.B2(n_240),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_229),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_224),
.B1(n_222),
.B2(n_247),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_254),
.B1(n_266),
.B2(n_259),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_263),
.B(n_262),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_247),
.C(n_225),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_316),
.C(n_282),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_225),
.C(n_222),
.Y(n_316)
);

OAI22x1_ASAP7_75t_SL g317 ( 
.A1(n_263),
.A2(n_224),
.B1(n_249),
.B2(n_233),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_265),
.B(n_233),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_326),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_337),
.C(n_339),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_330),
.B(n_291),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_331),
.B(n_356),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_344),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_288),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_335),
.A2(n_341),
.B(n_358),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_299),
.A2(n_271),
.B1(n_269),
.B2(n_277),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_343),
.B1(n_303),
.B2(n_304),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_255),
.C(n_273),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_346),
.B1(n_349),
.B2(n_354),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_316),
.A2(n_280),
.B(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_276),
.Y(n_342)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_321),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_268),
.C(n_249),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_347),
.C(n_353),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_281),
.B1(n_248),
.B2(n_239),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_239),
.C(n_198),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_293),
.A2(n_317),
.B1(n_320),
.B2(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_351),
.Y(n_380)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_313),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_352),
.B(n_355),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_295),
.B(n_248),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_290),
.A2(n_297),
.B1(n_306),
.B2(n_325),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_176),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_318),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_297),
.A2(n_75),
.B1(n_178),
.B2(n_161),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_311),
.B1(n_308),
.B2(n_303),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_48),
.B(n_45),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_305),
.B1(n_311),
.B2(n_325),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_361),
.A2(n_366),
.B1(n_372),
.B2(n_382),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_315),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_365),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_307),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_335),
.B1(n_354),
.B2(n_342),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_301),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_379),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_369),
.A2(n_326),
.B1(n_351),
.B2(n_348),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_329),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_376),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_373),
.B(n_9),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_381),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_301),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_334),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_336),
.A2(n_333),
.B1(n_337),
.B2(n_358),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_308),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_334),
.A2(n_298),
.B(n_324),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_384),
.A2(n_341),
.B(n_347),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_350),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_360),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_42),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_R g418 ( 
.A(n_389),
.B(n_370),
.C(n_374),
.Y(n_418)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_345),
.C(n_353),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_394),
.C(n_397),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_369),
.A2(n_357),
.B1(n_331),
.B2(n_330),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_403),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_319),
.C(n_204),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_36),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_396),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_48),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_32),
.C(n_42),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_32),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_412),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_7),
.B(n_15),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_410),
.Y(n_427)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_368),
.A2(n_42),
.B1(n_10),
.B2(n_11),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_408),
.A2(n_359),
.B1(n_375),
.B2(n_376),
.Y(n_423)
);

OA21x2_ASAP7_75t_SL g409 ( 
.A1(n_371),
.A2(n_42),
.B(n_6),
.Y(n_409)
);

NOR3xp33_ASAP7_75t_SL g424 ( 
.A(n_409),
.B(n_359),
.C(n_380),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_360),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_387),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_411),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_388),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_413),
.B(n_394),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_377),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_420),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_407),
.A2(n_368),
.B1(n_370),
.B2(n_384),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_424),
.Y(n_449)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_391),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_426),
.Y(n_447)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_382),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_398),
.B(n_366),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_389),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_407),
.A2(n_362),
.B1(n_381),
.B2(n_363),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_432),
.A2(n_431),
.B1(n_399),
.B2(n_427),
.Y(n_445)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_425),
.B(n_412),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_443),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_429),
.C(n_414),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_438),
.C(n_442),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_426),
.C(n_430),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_402),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_420),
.C(n_415),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_401),
.CI(n_392),
.CON(n_443),
.SN(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_401),
.C(n_393),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_448),
.C(n_438),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_445),
.A2(n_446),
.B1(n_408),
.B2(n_6),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_417),
.A2(n_421),
.B1(n_419),
.B2(n_432),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_397),
.C(n_396),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_390),
.C(n_378),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_454),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_413),
.C(n_361),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_460),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_456),
.A2(n_439),
.B1(n_443),
.B2(n_11),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_375),
.C(n_395),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_457),
.B(n_459),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_380),
.B(n_424),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_458),
.A2(n_464),
.B(n_443),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_416),
.C(n_386),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_404),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_448),
.C(n_440),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_463),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_13),
.C(n_12),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_437),
.Y(n_465)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g483 ( 
.A(n_466),
.B(n_467),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_469),
.B(n_0),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_0),
.C(n_1),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_474),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_451),
.A2(n_11),
.B(n_1),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_450),
.A2(n_11),
.B(n_1),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_475),
.A2(n_453),
.B(n_455),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_457),
.C(n_454),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_476),
.B(n_0),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_478),
.Y(n_490)
);

INVx6_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_484),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_485),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_473),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_0),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_479),
.A2(n_468),
.B(n_466),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_486),
.A2(n_489),
.B(n_471),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_476),
.B(n_467),
.Y(n_489)
);

AO21x1_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_465),
.B(n_483),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_493),
.C(n_2),
.Y(n_495)
);

O2A1O1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_487),
.A2(n_483),
.B(n_490),
.C(n_473),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_481),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_494),
.A2(n_495),
.B(n_3),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_496),
.A2(n_3),
.B(n_4),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_4),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_4),
.Y(n_499)
);


endmodule