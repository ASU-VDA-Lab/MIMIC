module real_aes_6596_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g546 ( .A1(n_0), .A2(n_153), .B(n_547), .C(n_550), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_1), .B(n_491), .Y(n_551) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g187 ( .A(n_3), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_4), .B(n_145), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_5), .A2(n_460), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_6), .A2(n_130), .B(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_7), .A2(n_35), .B1(n_139), .B2(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_8), .B(n_130), .Y(n_156) );
AND2x6_ASAP7_75t_L g154 ( .A(n_9), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_10), .A2(n_154), .B(n_450), .C(n_452), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_11), .B(n_36), .Y(n_110) );
INVx1_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
INVx1_ASAP7_75t_L g180 ( .A(n_13), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_14), .B(n_143), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_15), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_16), .B(n_145), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_17), .B(n_131), .Y(n_192) );
AO32x2_ASAP7_75t_L g214 ( .A1(n_18), .A2(n_130), .A3(n_160), .B1(n_171), .B2(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_19), .B(n_139), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_20), .B(n_131), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_21), .A2(n_53), .B1(n_139), .B2(n_217), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_22), .A2(n_80), .B1(n_139), .B2(n_143), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_23), .B(n_139), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_24), .A2(n_171), .B(n_450), .C(n_511), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_25), .A2(n_171), .B(n_450), .C(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_26), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_27), .B(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_28), .A2(n_460), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_29), .B(n_173), .Y(n_211) );
INVx2_ASAP7_75t_L g141 ( .A(n_30), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_31), .A2(n_462), .B(n_470), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_32), .B(n_139), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_33), .B(n_173), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_34), .B(n_225), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_37), .B(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_38), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_39), .A2(n_77), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_39), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_40), .B(n_145), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_41), .B(n_460), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_42), .A2(n_78), .B1(n_433), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_42), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_43), .A2(n_462), .B(n_464), .C(n_470), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_44), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g548 ( .A(n_45), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_46), .A2(n_89), .B1(n_217), .B2(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g465 ( .A(n_47), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_48), .B(n_139), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_49), .B(n_139), .Y(n_182) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_50), .A2(n_102), .B1(n_114), .B2(n_734), .C(n_740), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_50), .B(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_50), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_51), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_52), .B(n_151), .Y(n_150) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_54), .A2(n_58), .B1(n_139), .B2(n_143), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_55), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_56), .B(n_139), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_57), .B(n_139), .Y(n_222) );
INVx1_ASAP7_75t_L g155 ( .A(n_59), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_60), .B(n_460), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_61), .B(n_491), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_62), .A2(n_151), .B(n_183), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_63), .B(n_139), .Y(n_188) );
INVx1_ASAP7_75t_L g134 ( .A(n_64), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_65), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_66), .B(n_145), .Y(n_501) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_67), .A2(n_130), .A3(n_171), .B1(n_236), .B2(n_240), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_68), .B(n_146), .Y(n_453) );
INVx1_ASAP7_75t_L g166 ( .A(n_69), .Y(n_166) );
INVx1_ASAP7_75t_L g206 ( .A(n_70), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_71), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_72), .B(n_467), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_73), .A2(n_450), .B(n_470), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_74), .B(n_143), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_75), .Y(n_486) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_77), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_78), .A2(n_122), .B1(n_432), .B2(n_433), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_78), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_79), .B(n_466), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_81), .B(n_217), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_82), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_83), .B(n_143), .Y(n_210) );
INVx2_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_85), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_86), .B(n_170), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_87), .B(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g436 ( .A(n_88), .B(n_108), .Y(n_436) );
INVx2_ASAP7_75t_L g724 ( .A(n_88), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_90), .A2(n_100), .B1(n_143), .B2(n_144), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_91), .B(n_460), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_92), .Y(n_731) );
INVx1_ASAP7_75t_L g500 ( .A(n_93), .Y(n_500) );
INVxp67_ASAP7_75t_L g489 ( .A(n_94), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_95), .B(n_143), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g446 ( .A(n_97), .Y(n_446) );
INVx1_ASAP7_75t_L g524 ( .A(n_98), .Y(n_524) );
AND2x2_ASAP7_75t_L g472 ( .A(n_99), .B(n_173), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_105), .B(n_111), .Y(n_103) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_104), .B(n_112), .Y(n_737) );
INVx1_ASAP7_75t_L g758 ( .A(n_104), .Y(n_758) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g739 ( .A(n_106), .Y(n_739) );
INVx1_ASAP7_75t_SL g751 ( .A(n_106), .Y(n_751) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_107), .B(n_724), .Y(n_733) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g723 ( .A(n_108), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g756 ( .A(n_111), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OAI222xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_118), .B1(n_725), .B2(n_726), .C1(n_731), .C2(n_732), .Y(n_114) );
INVx1_ASAP7_75t_L g725 ( .A(n_115), .Y(n_725) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_434), .B1(n_437), .B2(n_721), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_121), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
INVx2_ASAP7_75t_L g432 ( .A(n_122), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_122), .A2(n_432), .B1(n_745), .B2(n_746), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g122 ( .A(n_123), .B(n_356), .Y(n_122) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_314), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_254), .C(n_290), .D(n_304), .Y(n_124) );
OAI221xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_198), .B1(n_230), .B2(n_241), .C(n_245), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_126), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_174), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_157), .Y(n_128) );
AND2x2_ASAP7_75t_L g251 ( .A(n_129), .B(n_158), .Y(n_251) );
INVx3_ASAP7_75t_L g259 ( .A(n_129), .Y(n_259) );
AND2x2_ASAP7_75t_L g313 ( .A(n_129), .B(n_177), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_129), .B(n_176), .Y(n_349) );
AND2x2_ASAP7_75t_L g407 ( .A(n_129), .B(n_269), .Y(n_407) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_136), .B(n_156), .Y(n_129) );
INVx4_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_130), .A2(n_477), .B(n_478), .Y(n_476) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_130), .Y(n_483) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_132), .B(n_133), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_148), .B(n_154), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_145), .Y(n_137) );
INVx3_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_139), .Y(n_526) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
BUFx3_ASAP7_75t_L g238 ( .A(n_140), .Y(n_238) );
AND2x6_ASAP7_75t_L g450 ( .A(n_140), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx1_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx2_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_145), .A2(n_163), .B(n_164), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_SL g204 ( .A1(n_145), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_145), .B(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g236 ( .A1(n_146), .A2(n_170), .B1(n_237), .B2(n_239), .Y(n_236) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
AND2x2_ASAP7_75t_L g448 ( .A(n_147), .B(n_152), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_147), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_153), .Y(n_148) );
INVx2_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_167), .B(n_187), .C(n_188), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_153), .A2(n_170), .B1(n_195), .B2(n_196), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_153), .A2(n_170), .B1(n_216), .B2(n_218), .Y(n_215) );
BUFx3_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_154), .A2(n_179), .B(n_186), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_154), .A2(n_204), .B(n_208), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_221), .B(n_226), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_154), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g460 ( .A(n_154), .B(n_448), .Y(n_460) );
INVx4_ASAP7_75t_SL g471 ( .A(n_154), .Y(n_471) );
AND2x2_ASAP7_75t_L g242 ( .A(n_157), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g256 ( .A(n_157), .B(n_177), .Y(n_256) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_158), .B(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_158), .B(n_259), .Y(n_283) );
OR2x2_ASAP7_75t_L g285 ( .A(n_158), .B(n_243), .Y(n_285) );
AND2x2_ASAP7_75t_L g320 ( .A(n_158), .B(n_243), .Y(n_320) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_158), .Y(n_365) );
INVx1_ASAP7_75t_L g373 ( .A(n_158), .Y(n_373) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_172), .Y(n_158) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_178), .B(n_189), .Y(n_177) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_160), .B(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_171), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_169), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_167), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g549 ( .A(n_170), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_171), .B(n_194), .C(n_197), .Y(n_193) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_173), .A2(n_203), .B(n_211), .Y(n_202) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_173), .A2(n_220), .B(n_229), .Y(n_219) );
INVx2_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_173), .A2(n_459), .B(n_461), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_173), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g517 ( .A(n_173), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_174), .A2(n_291), .B1(n_295), .B2(n_299), .C(n_300), .Y(n_290) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g250 ( .A(n_175), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_190), .Y(n_175) );
INVx2_ASAP7_75t_L g249 ( .A(n_176), .Y(n_249) );
AND2x2_ASAP7_75t_L g302 ( .A(n_176), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_176), .B(n_259), .Y(n_321) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g384 ( .A(n_177), .B(n_259), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_183), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_181), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_181), .A2(n_480), .B(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_183), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_184), .A2(n_209), .B(n_210), .Y(n_208) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g467 ( .A(n_185), .Y(n_467) );
AND2x2_ASAP7_75t_L g306 ( .A(n_190), .B(n_251), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g374 ( .A1(n_190), .A2(n_330), .A3(n_375), .B1(n_377), .B2(n_380), .C1(n_382), .C2(n_386), .Y(n_374) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_191), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
AND2x2_ASAP7_75t_L g379 ( .A(n_191), .B(n_259), .Y(n_379) );
AND2x2_ASAP7_75t_L g411 ( .A(n_191), .B(n_283), .Y(n_411) );
OR2x2_ASAP7_75t_L g414 ( .A(n_191), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g244 ( .A(n_192), .Y(n_244) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_197), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_197), .A2(n_445), .B(n_455), .Y(n_444) );
INVx3_ASAP7_75t_L g491 ( .A(n_197), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_197), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_197), .A2(n_521), .B(n_528), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_197), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_212), .Y(n_199) );
INVx1_ASAP7_75t_L g427 ( .A(n_200), .Y(n_427) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g232 ( .A(n_201), .B(n_219), .Y(n_232) );
INVx2_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g289 ( .A(n_202), .Y(n_289) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
OR2x2_ASAP7_75t_L g421 ( .A(n_202), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g246 ( .A(n_212), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g286 ( .A(n_212), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g338 ( .A(n_212), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_219), .Y(n_212) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_234), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_213), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g347 ( .A(n_213), .B(n_235), .Y(n_347) );
OR2x2_ASAP7_75t_L g355 ( .A(n_213), .B(n_289), .Y(n_355) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx2_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g298 ( .A(n_214), .B(n_219), .Y(n_298) );
AND2x2_ASAP7_75t_L g362 ( .A(n_214), .B(n_235), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_219), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
INVx1_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_219), .Y(n_370) );
INVx1_ASAP7_75t_L g422 ( .A(n_219), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g399 ( .A(n_231), .B(n_308), .Y(n_399) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g326 ( .A(n_233), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g425 ( .A(n_233), .B(n_360), .Y(n_425) );
INVx1_ASAP7_75t_L g247 ( .A(n_234), .Y(n_247) );
AND2x2_ASAP7_75t_L g273 ( .A(n_234), .B(n_267), .Y(n_273) );
BUFx2_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
INVx1_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_238), .Y(n_469) );
INVx2_ASAP7_75t_L g550 ( .A(n_238), .Y(n_550) );
INVx1_ASAP7_75t_L g514 ( .A(n_240), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_241), .B(n_248), .Y(n_401) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI32xp33_ASAP7_75t_L g245 ( .A1(n_242), .A2(n_246), .A3(n_248), .B1(n_250), .B2(n_252), .Y(n_245) );
AND2x2_ASAP7_75t_L g385 ( .A(n_242), .B(n_258), .Y(n_385) );
AND2x2_ASAP7_75t_L g423 ( .A(n_242), .B(n_321), .Y(n_423) );
INVx1_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_247), .B(n_309), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_248), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_248), .B(n_251), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_248), .B(n_320), .Y(n_402) );
OR2x2_ASAP7_75t_L g416 ( .A(n_248), .B(n_285), .Y(n_416) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g343 ( .A(n_249), .B(n_251), .Y(n_343) );
OR2x2_ASAP7_75t_L g352 ( .A(n_249), .B(n_339), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_251), .B(n_302), .Y(n_324) );
INVx2_ASAP7_75t_L g339 ( .A(n_253), .Y(n_339) );
OR2x2_ASAP7_75t_L g354 ( .A(n_253), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g369 ( .A(n_253), .B(n_370), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_253), .A2(n_346), .B(n_427), .C(n_428), .Y(n_426) );
OAI321xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_260), .A3(n_265), .B1(n_268), .B2(n_272), .C(n_276), .Y(n_254) );
INVx1_ASAP7_75t_L g367 ( .A(n_255), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g378 ( .A(n_256), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g330 ( .A(n_258), .Y(n_330) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_259), .B(n_373), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_260), .A2(n_398), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g335 ( .A(n_262), .B(n_309), .Y(n_335) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_263), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_265), .A2(n_306), .B(n_351), .C(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g317 ( .A(n_267), .B(n_274), .Y(n_317) );
BUFx2_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
INVx1_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OR2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g431 ( .A(n_270), .Y(n_431) );
INVx1_ASAP7_75t_L g424 ( .A(n_271), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g277 ( .A(n_273), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g381 ( .A(n_273), .B(n_298), .Y(n_381) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_284), .B2(n_286), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g346 ( .A(n_279), .B(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_280), .B(n_289), .Y(n_309) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g311 ( .A(n_285), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_288), .A2(n_406), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g294 ( .A(n_289), .Y(n_294) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_289), .Y(n_360) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_292), .B(n_411), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_293), .A2(n_298), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_296), .B(n_306), .Y(n_403) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g372 ( .A(n_297), .Y(n_372) );
AND2x2_ASAP7_75t_L g331 ( .A(n_298), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g420 ( .A(n_298), .Y(n_420) );
INVx1_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
INVx1_ASAP7_75t_L g391 ( .A(n_302), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_310), .B2(n_311), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_308), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_309), .B(n_347), .Y(n_413) );
OR2x2_ASAP7_75t_L g386 ( .A(n_310), .B(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g325 ( .A(n_311), .Y(n_325) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_313), .B(n_364), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_333), .C(n_344), .Y(n_314) );
OAI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B(n_322), .C(n_328), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_317), .A2(n_388), .B1(n_392), .B2(n_395), .C(n_397), .Y(n_387) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_320), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g383 ( .A(n_320), .B(n_384), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_321), .A2(n_369), .B(n_371), .C(n_373), .Y(n_368) );
INVx2_ASAP7_75t_L g415 ( .A(n_321), .Y(n_415) );
OAI21xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_325), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g394 ( .A(n_327), .B(n_347), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B(n_337), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_343), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_338), .B(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_343), .B(n_430), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B(n_350), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g371 ( .A(n_347), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND4x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_387), .C(n_404), .D(n_426), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_374), .Y(n_357) );
OAI211xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_363), .B(n_366), .C(n_368), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_362), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_373), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx2_ASAP7_75t_SL g396 ( .A(n_384), .Y(n_396) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g409 ( .A(n_394), .Y(n_409) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_412), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_417), .C(n_418), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g728 ( .A(n_435), .Y(n_728) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g729 ( .A(n_437), .Y(n_729) );
OR3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_619), .C(n_684), .Y(n_437) );
NAND4xp25_ASAP7_75t_SL g438 ( .A(n_439), .B(n_560), .C(n_586), .D(n_609), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_492), .B1(n_530), .B2(n_537), .C(n_552), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_441), .A2(n_553), .B1(n_577), .B2(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_473), .Y(n_441) );
INVx1_ASAP7_75t_SL g613 ( .A(n_442), .Y(n_613) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_457), .Y(n_442) );
OR2x2_ASAP7_75t_L g535 ( .A(n_443), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g555 ( .A(n_443), .B(n_474), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_443), .B(n_482), .Y(n_568) );
AND2x2_ASAP7_75t_L g585 ( .A(n_443), .B(n_457), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_443), .B(n_533), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_443), .B(n_584), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_443), .B(n_473), .Y(n_706) );
AOI211xp5_ASAP7_75t_SL g717 ( .A1(n_443), .A2(n_623), .B(n_718), .C(n_719), .Y(n_717) );
INVx5_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_444), .B(n_474), .Y(n_589) );
AND2x2_ASAP7_75t_L g592 ( .A(n_444), .B(n_475), .Y(n_592) );
OR2x2_ASAP7_75t_L g637 ( .A(n_444), .B(n_474), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_444), .B(n_482), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
INVx5_ASAP7_75t_L g463 ( .A(n_450), .Y(n_463) );
INVx5_ASAP7_75t_SL g536 ( .A(n_457), .Y(n_536) );
AND2x2_ASAP7_75t_L g554 ( .A(n_457), .B(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_457), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_457), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g672 ( .A(n_457), .B(n_482), .Y(n_672) );
OR2x2_ASAP7_75t_L g678 ( .A(n_457), .B(n_568), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_457), .B(n_628), .Y(n_687) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
BUFx2_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_463), .A2(n_471), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_463), .A2(n_471), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_468), .C(n_469), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_466), .A2(n_469), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
AND2x2_ASAP7_75t_L g569 ( .A(n_474), .B(n_536), .Y(n_569) );
INVx1_ASAP7_75t_SL g582 ( .A(n_474), .Y(n_582) );
OR2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g623 ( .A(n_474), .B(n_482), .Y(n_623) );
AND2x2_ASAP7_75t_L g681 ( .A(n_474), .B(n_533), .Y(n_681) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_475), .B(n_536), .Y(n_608) );
INVx3_ASAP7_75t_L g533 ( .A(n_482), .Y(n_533) );
OR2x2_ASAP7_75t_L g574 ( .A(n_482), .B(n_536), .Y(n_574) );
AND2x2_ASAP7_75t_L g584 ( .A(n_482), .B(n_582), .Y(n_584) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_482), .Y(n_632) );
AND2x2_ASAP7_75t_L g641 ( .A(n_482), .B(n_555), .Y(n_641) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_490), .Y(n_482) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_491), .A2(n_543), .B(n_551), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_492), .A2(n_658), .B1(n_660), .B2(n_662), .C(n_665), .Y(n_657) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
AND2x2_ASAP7_75t_L g631 ( .A(n_494), .B(n_612), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_494), .B(n_690), .Y(n_694) );
OR2x2_ASAP7_75t_L g715 ( .A(n_494), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_494), .B(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx5_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
AND2x2_ASAP7_75t_L g639 ( .A(n_495), .B(n_506), .Y(n_639) );
AND2x2_ASAP7_75t_L g700 ( .A(n_495), .B(n_579), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_495), .B(n_533), .Y(n_713) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_518), .Y(n_504) );
AND2x4_ASAP7_75t_L g540 ( .A(n_505), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
AND2x2_ASAP7_75t_L g634 ( .A(n_505), .B(n_612), .Y(n_634) );
AND2x2_ASAP7_75t_L g644 ( .A(n_505), .B(n_562), .Y(n_644) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_505), .Y(n_652) );
AND2x2_ASAP7_75t_L g664 ( .A(n_505), .B(n_542), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_505), .B(n_596), .Y(n_668) );
AND2x2_ASAP7_75t_L g705 ( .A(n_505), .B(n_700), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_505), .B(n_579), .Y(n_716) );
OR2x2_ASAP7_75t_L g718 ( .A(n_505), .B(n_654), .Y(n_718) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g604 ( .A(n_506), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g614 ( .A(n_506), .B(n_559), .Y(n_614) );
AND2x2_ASAP7_75t_L g626 ( .A(n_506), .B(n_542), .Y(n_626) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_506), .Y(n_656) );
AND2x4_ASAP7_75t_L g690 ( .A(n_506), .B(n_541), .Y(n_690) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_510), .B(n_514), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
BUFx2_ASAP7_75t_L g539 ( .A(n_518), .Y(n_539) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
AND2x2_ASAP7_75t_L g612 ( .A(n_519), .B(n_542), .Y(n_612) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g559 ( .A(n_520), .B(n_542), .Y(n_559) );
BUFx2_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_532), .B(n_613), .Y(n_692) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_533), .B(n_555), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_533), .B(n_536), .Y(n_594) );
AND2x2_ASAP7_75t_L g649 ( .A(n_533), .B(n_585), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g586 ( .A1(n_534), .A2(n_587), .B1(n_595), .B2(n_597), .C(n_601), .Y(n_586) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g581 ( .A(n_535), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g622 ( .A(n_535), .B(n_623), .Y(n_622) );
OAI321xp33_ASAP7_75t_L g629 ( .A1(n_535), .A2(n_588), .A3(n_630), .B1(n_632), .B2(n_633), .C(n_635), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_536), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_539), .B(n_690), .Y(n_708) );
AND2x2_ASAP7_75t_L g595 ( .A(n_540), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_540), .B(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_541), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_541), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_541), .B(n_653), .Y(n_683) );
INVx1_ASAP7_75t_L g720 ( .A(n_541), .Y(n_720) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_557), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_554), .A2(n_664), .B(n_713), .C(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_555), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_555), .B(n_593), .Y(n_659) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_559), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_559), .B(n_562), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_559), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_559), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B1(n_575), .B2(n_580), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g576 ( .A(n_562), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g599 ( .A(n_562), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_562), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_605), .Y(n_647) );
OR2x2_ASAP7_75t_L g654 ( .A(n_562), .B(n_579), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_562), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g704 ( .A(n_562), .B(n_690), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_570), .B2(n_572), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g610 ( .A(n_565), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_568), .A2(n_583), .B1(n_651), .B2(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g698 ( .A(n_569), .Y(n_698) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_573), .A2(n_610), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_609) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g588 ( .A(n_574), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_578), .B(n_644), .Y(n_676) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_579), .Y(n_596) );
INVx1_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g618 ( .A(n_585), .Y(n_618) );
AND2x2_ASAP7_75t_L g627 ( .A(n_585), .B(n_628), .Y(n_627) );
NAND2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g671 ( .A(n_592), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_595), .A2(n_621), .B1(n_624), .B2(n_627), .C(n_629), .Y(n_620) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_599), .B(n_656), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_603), .B(n_606), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_606), .Y(n_703) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g666 ( .A(n_611), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_611), .B(n_671), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_614), .B(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_638), .C(n_657), .D(n_670), .Y(n_619) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g628 ( .A(n_623), .Y(n_628) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g661 ( .A(n_632), .B(n_637), .Y(n_661) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_642), .C(n_650), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_640), .A2(n_682), .B(n_710), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_SL g669 ( .A(n_641), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g673 ( .A(n_647), .Y(n_673) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_653), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_653), .B(n_664), .Y(n_697) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g674 ( .A(n_664), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B(n_669), .Y(n_665) );
INVxp33_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .A3(n_674), .B1(n_675), .B2(n_677), .C1(n_679), .C2(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_685), .B(n_702), .C(n_709), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g701 ( .A(n_690), .Y(n_701) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .C(n_707), .Y(n_702) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g730 ( .A(n_722), .Y(n_730) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_738), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
AOI21xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_752), .B(n_755), .Y(n_740) );
INVxp33_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_748), .C(n_751), .Y(n_742) );
INVx1_ASAP7_75t_L g750 ( .A(n_744), .Y(n_750) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
endmodule