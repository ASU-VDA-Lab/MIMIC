module fake_netlist_6_1564_n_979 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_979);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_979;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_923;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_608;
wire n_683;
wire n_620;
wire n_420;
wire n_261;
wire n_630;
wire n_394;
wire n_312;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_231;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_882;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_651;
wire n_271;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_385;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_649;
wire n_855;
wire n_283;

INVx2_ASAP7_75t_SL g195 ( 
.A(n_24),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_35),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_64),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_21),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_71),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_60),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_154),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_47),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_33),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_126),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_141),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_161),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_103),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_7),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_151),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_36),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_75),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_100),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_5),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_73),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_107),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_24),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_109),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_83),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_112),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_12),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_69),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_119),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_169),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_62),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_108),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_187),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_3),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_147),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_48),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_172),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_97),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_80),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_135),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_28),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_78),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_105),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_98),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_118),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_21),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_59),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_193),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_176),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_122),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_153),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_174),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_3),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_95),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_58),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_179),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_181),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_214),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_204),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_230),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_246),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_260),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_278),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_285),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_196),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_219),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_199),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_197),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_211),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_212),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_227),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_198),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_226),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_238),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_240),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_241),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_244),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_250),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_201),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_249),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_252),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_258),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_222),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_236),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_242),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_268),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_202),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_266),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_270),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_276),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_273),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_287),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_302),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_228),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_206),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_291),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_291),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_218),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_373),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_374),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_377),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_229),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_379),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_359),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_217),
.B(n_259),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_308),
.A2(n_203),
.B1(n_223),
.B2(n_232),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_308),
.A2(n_305),
.B1(n_207),
.B2(n_303),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_208),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_310),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_209),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_210),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_315),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_300),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_304),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

CKINVDCx6p67_ASAP7_75t_R g414 ( 
.A(n_366),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_361),
.A2(n_262),
.B1(n_299),
.B2(n_298),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_316),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_213),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_321),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

CKINVDCx11_ASAP7_75t_R g423 ( 
.A(n_331),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_343),
.B(n_304),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_215),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_359),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_341),
.B(n_304),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_354),
.A2(n_220),
.B(n_216),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_344),
.B(n_221),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_423),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_414),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_432),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_432),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_404),
.B(n_304),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_386),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_R g456 ( 
.A(n_391),
.B(n_362),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_431),
.B(n_362),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_400),
.B(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_408),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_395),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_350),
.Y(n_466)
);

NOR2x1p5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_352),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_421),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_395),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_426),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_416),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_403),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_399),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_419),
.B(n_325),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_405),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_407),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_402),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_383),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_R g482 ( 
.A(n_441),
.B(n_375),
.Y(n_482)
);

NOR2x1p5_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_352),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_410),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_427),
.B(n_326),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_399),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_398),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_434),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_404),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_404),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_404),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_404),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_404),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_387),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_387),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_387),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_387),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_411),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_411),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_415),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_388),
.B(n_311),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_508),
.B(n_438),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_496),
.B(n_331),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_L g516 ( 
.A(n_476),
.B(n_320),
.C(n_319),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_466),
.B(n_412),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_311),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_509),
.B(n_396),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_449),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_504),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_460),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_412),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_461),
.B(n_312),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_483),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_480),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_319),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_489),
.A2(n_438),
.B1(n_396),
.B2(n_349),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_471),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_468),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_469),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_477),
.B(n_388),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_500),
.B(n_312),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_388),
.Y(n_551)
);

NAND3x1_ASAP7_75t_L g552 ( 
.A(n_475),
.B(n_357),
.C(n_356),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_320),
.C(n_381),
.Y(n_553)
);

NAND3x1_ASAP7_75t_L g554 ( 
.A(n_475),
.B(n_357),
.C(n_356),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_487),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_505),
.B(n_360),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_506),
.B(n_388),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_442),
.B(n_445),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_346),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_486),
.A2(n_438),
.B1(n_297),
.B2(n_259),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_493),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_507),
.B(n_412),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_457),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_473),
.B(n_259),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_448),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_452),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

OR2x2_ASAP7_75t_SL g573 ( 
.A(n_458),
.B(n_438),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_454),
.B(n_415),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_462),
.B(n_413),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_454),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_464),
.B(n_413),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_317),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_490),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_496),
.B(n_317),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_526),
.A2(n_481),
.B(n_501),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_549),
.B(n_497),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_535),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_549),
.B(n_464),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_517),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_535),
.B(n_450),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_551),
.B(n_582),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_465),
.Y(n_594)
);

INVx8_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_551),
.B(n_494),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_534),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_529),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_574),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_470),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_550),
.B(n_323),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_569),
.A2(n_491),
.B1(n_472),
.B2(n_478),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_576),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_557),
.B(n_495),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_557),
.B(n_459),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_569),
.A2(n_491),
.B1(n_498),
.B2(n_497),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_538),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_467),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_532),
.B(n_482),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_514),
.B(n_472),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_545),
.B(n_498),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_547),
.B(n_478),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_534),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_548),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_514),
.A2(n_323),
.B1(n_451),
.B2(n_501),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_501),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_561),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_501),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_524),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_566),
.Y(n_627)
);

OAI221xp5_ASAP7_75t_L g628 ( 
.A1(n_563),
.A2(n_365),
.B1(n_369),
.B2(n_370),
.C(n_422),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_559),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_519),
.B(n_527),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_519),
.B(n_413),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_527),
.B(n_418),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_524),
.A2(n_451),
.B1(n_439),
.B2(n_428),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_539),
.B(n_418),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_540),
.B(n_444),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_515),
.A2(n_445),
.B1(n_440),
.B2(n_418),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_575),
.B(n_440),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_530),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_575),
.B(n_440),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_577),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_539),
.B(n_428),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_613),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_588),
.B(n_516),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_641),
.A2(n_556),
.B(n_571),
.C(n_570),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_589),
.A2(n_526),
.B(n_520),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_589),
.A2(n_546),
.B(n_520),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_599),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_592),
.B(n_584),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_629),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_605),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_615),
.A2(n_546),
.B(n_520),
.Y(n_656)
);

OAI321xp33_ASAP7_75t_L g657 ( 
.A1(n_603),
.A2(n_563),
.A3(n_584),
.B1(n_542),
.B2(n_553),
.C(n_583),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_601),
.B(n_515),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_607),
.B(n_559),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_615),
.A2(n_546),
.B(n_520),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_630),
.A2(n_585),
.B(n_546),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_594),
.B(n_558),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_643),
.B(n_581),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_593),
.B(n_581),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_586),
.A2(n_585),
.B(n_568),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_610),
.B(n_581),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_626),
.A2(n_585),
.B(n_568),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_614),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_638),
.B(n_536),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_596),
.A2(n_585),
.B(n_542),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_606),
.A2(n_577),
.B(n_530),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_619),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_608),
.A2(n_573),
.B1(n_554),
.B2(n_552),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_623),
.A2(n_624),
.B(n_627),
.C(n_587),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_631),
.A2(n_521),
.B(n_518),
.Y(n_675)
);

AOI21xp33_ASAP7_75t_L g676 ( 
.A1(n_591),
.A2(n_537),
.B(n_528),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_634),
.A2(n_642),
.B(n_639),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_620),
.A2(n_572),
.B(n_579),
.C(n_543),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_597),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_639),
.A2(n_579),
.B(n_543),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_616),
.B(n_541),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_604),
.B(n_524),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_642),
.A2(n_524),
.B(n_533),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_598),
.B(n_533),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_567),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_597),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_644),
.A2(n_567),
.B(n_425),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_602),
.A2(n_533),
.B1(n_567),
.B2(n_297),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_609),
.B(n_560),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_612),
.A2(n_412),
.B(n_425),
.C(n_420),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_632),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_622),
.A2(n_567),
.B(n_425),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_611),
.B(n_533),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_621),
.B(n_224),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_650),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_677),
.A2(n_625),
.B(n_595),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_645),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_646),
.B(n_618),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_683),
.A2(n_595),
.B(n_636),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_653),
.B(n_618),
.Y(n_700)
);

OAI22x1_ASAP7_75t_L g701 ( 
.A1(n_658),
.A2(n_637),
.B1(n_621),
.B2(n_635),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_672),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_668),
.A2(n_633),
.B1(n_618),
.B2(n_617),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_662),
.B(n_633),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_655),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_654),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_669),
.A2(n_628),
.B(n_420),
.C(n_422),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_657),
.A2(n_430),
.B(n_389),
.C(n_382),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_633),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_674),
.B(n_640),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_664),
.B(n_567),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_673),
.B(n_610),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_673),
.B(n_430),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_683),
.A2(n_595),
.B(n_425),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_686),
.B(n_409),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_SL g716 ( 
.A(n_657),
.B(n_681),
.C(n_659),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_647),
.B(n_610),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_652),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_689),
.B(n_541),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_691),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_682),
.B(n_409),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_676),
.B(n_382),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_685),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_648),
.Y(n_724)
);

BUFx4f_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_666),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_666),
.B(n_225),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_648),
.B(n_389),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_679),
.Y(n_729)
);

NOR2x1_ASAP7_75t_L g730 ( 
.A(n_686),
.B(n_390),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_679),
.B(n_231),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_678),
.A2(n_281),
.B1(n_234),
.B2(n_237),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_685),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_671),
.B(n_390),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_670),
.A2(n_282),
.B(n_247),
.C(n_248),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_693),
.A2(n_684),
.B1(n_688),
.B2(n_692),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_694),
.B(n_233),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_698),
.B(n_680),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_717),
.A2(n_704),
.B(n_713),
.C(n_700),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_721),
.A2(n_690),
.B(n_687),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_696),
.A2(n_649),
.B(n_667),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_696),
.A2(n_665),
.B(n_651),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_695),
.B(n_697),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_736),
.A2(n_660),
.A3(n_656),
.B(n_675),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_709),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_734),
.A2(n_661),
.B(n_429),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_699),
.A2(n_392),
.B(n_401),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_725),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_712),
.B(n_718),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_699),
.A2(n_259),
.A3(n_297),
.B(n_2),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_702),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_714),
.A2(n_392),
.B(n_401),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_723),
.B(n_428),
.Y(n_753)
);

NOR4xp25_ASAP7_75t_L g754 ( 
.A(n_735),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_720),
.B(n_253),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_714),
.A2(n_433),
.B(n_429),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_706),
.Y(n_758)
);

AOI21x1_ASAP7_75t_SL g759 ( 
.A1(n_737),
.A2(n_255),
.B(n_254),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_711),
.A2(n_433),
.B(n_429),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_716),
.A2(n_289),
.B(n_261),
.C(n_263),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_SL g762 ( 
.A1(n_719),
.A2(n_726),
.B(n_732),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_731),
.B(n_257),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_SL g764 ( 
.A1(n_703),
.A2(n_392),
.B(n_297),
.C(n_6),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_721),
.A2(n_297),
.A3(n_5),
.B(n_8),
.Y(n_765)
);

AND2x2_ASAP7_75t_SL g766 ( 
.A(n_725),
.B(n_429),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_727),
.B(n_264),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_297),
.B(n_383),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_716),
.A2(n_284),
.B(n_269),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_SL g770 ( 
.A1(n_707),
.A2(n_439),
.B(n_436),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_708),
.A2(n_383),
.B(n_384),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_SL g772 ( 
.A(n_722),
.B(n_265),
.C(n_271),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_723),
.B(n_272),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_707),
.A2(n_383),
.B(n_384),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_705),
.B(n_279),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_701),
.A2(n_439),
.B(n_436),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_729),
.B(n_280),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_715),
.A2(n_730),
.B(n_724),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_SL g779 ( 
.A(n_733),
.B(n_283),
.C(n_290),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_715),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_728),
.A2(n_294),
.B(n_296),
.C(n_733),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_728),
.A2(n_383),
.B(n_384),
.Y(n_782)
);

OAI22x1_ASAP7_75t_L g783 ( 
.A1(n_717),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_714),
.A2(n_439),
.B(n_436),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_700),
.B(n_429),
.Y(n_785)
);

NOR4xp25_ASAP7_75t_L g786 ( 
.A(n_717),
.B(n_4),
.C(n_9),
.D(n_10),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_721),
.A2(n_439),
.B(n_436),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_749),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_741),
.A2(n_385),
.B(n_384),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_762),
.B(n_739),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_783),
.A2(n_436),
.B1(n_433),
.B2(n_397),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_763),
.A2(n_433),
.B1(n_11),
.B2(n_12),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_748),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_769),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_742),
.A2(n_385),
.B(n_384),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_740),
.A2(n_433),
.B(n_385),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_751),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_750),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_774),
.A2(n_397),
.B(n_385),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_745),
.B(n_748),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_748),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_743),
.B(n_13),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_786),
.B(n_15),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_755),
.B(n_385),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_755),
.B(n_397),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_766),
.B(n_397),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_738),
.B(n_15),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_784),
.A2(n_397),
.B(n_124),
.Y(n_808)
);

CKINVDCx6p67_ASAP7_75t_R g809 ( 
.A(n_777),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_770),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_747),
.A2(n_121),
.B(n_190),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_758),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_761),
.A2(n_16),
.B(n_17),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_750),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_785),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_778),
.B(n_39),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_752),
.A2(n_125),
.B(n_189),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_750),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_772),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_771),
.A2(n_20),
.B(n_22),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_765),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_764),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_775),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_781),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_780),
.B(n_40),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_815),
.B(n_765),
.Y(n_826)
);

AO31x2_ASAP7_75t_L g827 ( 
.A1(n_798),
.A2(n_776),
.A3(n_757),
.B(n_760),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_814),
.Y(n_828)
);

AO21x2_ASAP7_75t_L g829 ( 
.A1(n_796),
.A2(n_787),
.B(n_746),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_797),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_797),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_812),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_790),
.B(n_754),
.Y(n_833)
);

AO21x2_ASAP7_75t_L g834 ( 
.A1(n_818),
.A2(n_768),
.B(n_782),
.Y(n_834)
);

OA21x2_ASAP7_75t_L g835 ( 
.A1(n_789),
.A2(n_773),
.B(n_756),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_821),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_810),
.A2(n_767),
.B(n_759),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_814),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_816),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_809),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_815),
.B(n_765),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_788),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_790),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_789),
.Y(n_844)
);

NOR2x1_ASAP7_75t_SL g845 ( 
.A(n_807),
.B(n_753),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_800),
.B(n_744),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_810),
.A2(n_753),
.B(n_744),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_800),
.B(n_744),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_800),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_813),
.A2(n_753),
.B(n_779),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_823),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_795),
.A2(n_753),
.B(n_130),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_795),
.A2(n_129),
.B(n_188),
.Y(n_853)
);

INVx8_ASAP7_75t_L g854 ( 
.A(n_825),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_820),
.Y(n_855)
);

AND3x2_ASAP7_75t_L g856 ( 
.A(n_802),
.B(n_26),
.C(n_27),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_830),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_831),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_836),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_848),
.B(n_820),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_855),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_838),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

AO21x2_ASAP7_75t_L g864 ( 
.A1(n_855),
.A2(n_808),
.B(n_822),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_846),
.B(n_820),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_828),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_828),
.B(n_802),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_826),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_826),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_826),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_841),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_841),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_854),
.Y(n_873)
);

CKINVDCx6p67_ASAP7_75t_R g874 ( 
.A(n_873),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_867),
.A2(n_803),
.B1(n_833),
.B2(n_843),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_866),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_867),
.B(n_841),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_870),
.A2(n_803),
.B1(n_850),
.B2(n_819),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_873),
.Y(n_879)
);

CKINVDCx11_ASAP7_75t_R g880 ( 
.A(n_873),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_864),
.A2(n_794),
.B1(n_840),
.B2(n_842),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_873),
.A2(n_819),
.B1(n_791),
.B2(n_840),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_873),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_864),
.A2(n_792),
.B1(n_856),
.B2(n_824),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_877),
.B(n_870),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_876),
.B(n_862),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_883),
.B(n_872),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_879),
.B(n_872),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_874),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_880),
.B(n_868),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_886),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_885),
.B(n_868),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_887),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_SL g894 ( 
.A1(n_889),
.A2(n_882),
.B1(n_845),
.B2(n_854),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_886),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_890),
.B(n_869),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_887),
.B(n_875),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_893),
.B(n_888),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_897),
.B(n_878),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_896),
.B(n_869),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_895),
.B(n_881),
.Y(n_901)
);

AOI331xp33_ASAP7_75t_L g902 ( 
.A1(n_891),
.A2(n_884),
.A3(n_859),
.B1(n_791),
.B2(n_858),
.B3(n_881),
.C1(n_847),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_892),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_898),
.B(n_897),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_903),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_901),
.B(n_894),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_899),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_904),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_907),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_904),
.B(n_902),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_906),
.A2(n_901),
.B1(n_884),
.B2(n_842),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_905),
.B(n_900),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_910),
.A2(n_908),
.B(n_911),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_909),
.A2(n_851),
.B1(n_839),
.B2(n_860),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_912),
.B(n_832),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_911),
.A2(n_851),
.B1(n_839),
.B2(n_860),
.Y(n_916)
);

AO22x1_ASAP7_75t_L g917 ( 
.A1(n_908),
.A2(n_793),
.B1(n_801),
.B2(n_825),
.Y(n_917)
);

OAI32xp33_ASAP7_75t_L g918 ( 
.A1(n_910),
.A2(n_865),
.A3(n_871),
.B1(n_863),
.B2(n_793),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_909),
.B(n_871),
.Y(n_919)
);

NOR2x1_ASAP7_75t_L g920 ( 
.A(n_913),
.B(n_801),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_915),
.B(n_865),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_919),
.B(n_857),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_916),
.A2(n_854),
.B1(n_864),
.B2(n_837),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_914),
.B(n_27),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_917),
.B(n_29),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_918),
.B(n_863),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_915),
.B(n_29),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_913),
.A2(n_863),
.B(n_816),
.C(n_825),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_927),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_925),
.Y(n_930)
);

NAND4xp25_ASAP7_75t_L g931 ( 
.A(n_920),
.B(n_816),
.C(n_849),
.D(n_848),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_924),
.A2(n_848),
.B1(n_861),
.B2(n_857),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_928),
.B(n_926),
.Y(n_933)
);

AOI322xp5_ASAP7_75t_L g934 ( 
.A1(n_923),
.A2(n_861),
.A3(n_32),
.B1(n_30),
.B2(n_844),
.C1(n_829),
.C2(n_827),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_921),
.B(n_30),
.Y(n_935)
);

OAI221xp5_ASAP7_75t_L g936 ( 
.A1(n_922),
.A2(n_806),
.B1(n_835),
.B2(n_804),
.C(n_805),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_924),
.A2(n_835),
.B1(n_829),
.B2(n_806),
.Y(n_937)
);

AOI33xp33_ASAP7_75t_L g938 ( 
.A1(n_923),
.A2(n_32),
.A3(n_844),
.B1(n_43),
.B2(n_45),
.B3(n_51),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_930),
.A2(n_835),
.B1(n_852),
.B2(n_853),
.Y(n_939)
);

AOI221x1_ASAP7_75t_L g940 ( 
.A1(n_929),
.A2(n_935),
.B1(n_933),
.B2(n_931),
.C(n_938),
.Y(n_940)
);

OAI221xp5_ASAP7_75t_L g941 ( 
.A1(n_932),
.A2(n_805),
.B1(n_804),
.B2(n_799),
.C(n_57),
.Y(n_941)
);

AOI32xp33_ASAP7_75t_L g942 ( 
.A1(n_936),
.A2(n_817),
.A3(n_808),
.B1(n_811),
.B2(n_827),
.Y(n_942)
);

AOI221xp5_ASAP7_75t_L g943 ( 
.A1(n_937),
.A2(n_834),
.B1(n_52),
.B2(n_56),
.C(n_61),
.Y(n_943)
);

NOR4xp25_ASAP7_75t_L g944 ( 
.A(n_934),
.B(n_42),
.C(n_63),
.D(n_65),
.Y(n_944)
);

AOI21xp33_ASAP7_75t_SL g945 ( 
.A1(n_930),
.A2(n_66),
.B(n_67),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_930),
.A2(n_68),
.B(n_74),
.C(n_76),
.Y(n_946)
);

OAI221xp5_ASAP7_75t_L g947 ( 
.A1(n_930),
.A2(n_799),
.B1(n_81),
.B2(n_82),
.C(n_85),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_940),
.A2(n_799),
.B(n_87),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_945),
.Y(n_949)
);

OAI222xp33_ASAP7_75t_L g950 ( 
.A1(n_941),
.A2(n_827),
.B1(n_88),
.B2(n_89),
.C1(n_90),
.C2(n_91),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_943),
.A2(n_834),
.B1(n_827),
.B2(n_93),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_947),
.C(n_944),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_939),
.A2(n_79),
.B1(n_92),
.B2(n_101),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_942),
.A2(n_106),
.B1(n_111),
.B2(n_114),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_949),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_948),
.A2(n_952),
.B(n_954),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_953),
.B(n_115),
.Y(n_957)
);

OAI221xp5_ASAP7_75t_L g958 ( 
.A1(n_955),
.A2(n_951),
.B1(n_950),
.B2(n_120),
.C(n_127),
.Y(n_958)
);

NAND2x1_ASAP7_75t_L g959 ( 
.A(n_956),
.B(n_116),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_L g960 ( 
.A(n_957),
.B(n_117),
.C(n_128),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_959),
.A2(n_960),
.B(n_958),
.C(n_134),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_959),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_962),
.B(n_131),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_961),
.Y(n_964)
);

OAI211xp5_ASAP7_75t_SL g965 ( 
.A1(n_964),
.A2(n_133),
.B(n_138),
.C(n_139),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_963),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_966),
.B(n_146),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_965),
.B(n_148),
.Y(n_968)
);

XNOR2xp5_ASAP7_75t_L g969 ( 
.A(n_968),
.B(n_149),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_969),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_970),
.B(n_967),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_971),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_972),
.B(n_152),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_973),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_974),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_SL g976 ( 
.A1(n_975),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_976),
.A2(n_192),
.B(n_164),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_977),
.A2(n_160),
.B1(n_167),
.B2(n_168),
.Y(n_978)
);

AOI211xp5_ASAP7_75t_L g979 ( 
.A1(n_978),
.A2(n_173),
.B(n_177),
.C(n_178),
.Y(n_979)
);


endmodule