module fake_netlist_5_2119_n_793 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_793);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_793;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_728;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

BUFx2_ASAP7_75t_L g158 ( 
.A(n_26),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_71),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_20),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_59),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_13),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_18),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_60),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_82),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_53),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_64),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_17),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_23),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_58),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_102),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_77),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_22),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_0),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_27),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_194),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_29),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_1),
.B(n_2),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_251)
);

BUFx8_ASAP7_75t_SL g252 ( 
.A(n_171),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_173),
.B(n_174),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_255),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_187),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_187),
.Y(n_266)
);

CKINVDCx6p67_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_255),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

NOR2x1p5_ASAP7_75t_L g277 ( 
.A(n_222),
.B(n_162),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_224),
.B(n_207),
.C(n_210),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_231),
.B(n_190),
.Y(n_289)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_211),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_L g298 ( 
.A(n_215),
.B(n_207),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_255),
.B(n_190),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_244),
.B(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_243),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_247),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_247),
.Y(n_311)
);

NAND2x1p5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_216),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_244),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g314 ( 
.A(n_259),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_247),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_238),
.C(n_254),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_289),
.A2(n_249),
.B(n_221),
.C(n_216),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_215),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_263),
.B(n_242),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_242),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_267),
.B(n_245),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_282),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_216),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_221),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_282),
.B(n_221),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_277),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_295),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_229),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_259),
.B(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_219),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_260),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_253),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_253),
.C(n_256),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_235),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_275),
.B(n_215),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_275),
.B(n_215),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_227),
.Y(n_347)
);

OAI221xp5_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_234),
.B1(n_236),
.B2(n_217),
.C(n_226),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_220),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_220),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_249),
.B(n_248),
.C(n_241),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_267),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_220),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_241),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_220),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_L g359 ( 
.A(n_301),
.B(n_210),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_239),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_159),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_280),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_271),
.B(n_160),
.Y(n_364)
);

INVx8_ASAP7_75t_L g365 ( 
.A(n_280),
.Y(n_365)
);

NOR3xp33_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_191),
.C(n_213),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_239),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_246),
.B(n_248),
.C(n_209),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_261),
.B(n_258),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_307),
.B(n_269),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_325),
.A2(n_276),
.B(n_265),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_269),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_272),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_288),
.B(n_278),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_272),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_363),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_318),
.A2(n_246),
.B(n_226),
.C(n_283),
.Y(n_379)
);

INVx11_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_279),
.B(n_281),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_262),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_306),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_311),
.A2(n_286),
.B(n_284),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_322),
.B(n_334),
.Y(n_386)
);

BUFx4f_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_317),
.A2(n_204),
.B1(n_176),
.B2(n_178),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_316),
.A2(n_286),
.B(n_284),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_352),
.A2(n_274),
.B(n_262),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_338),
.A2(n_324),
.B(n_344),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_346),
.A2(n_274),
.B(n_268),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_335),
.A2(n_200),
.B1(n_181),
.B2(n_183),
.Y(n_399)
);

AO21x1_ASAP7_75t_L g400 ( 
.A1(n_317),
.A2(n_366),
.B(n_313),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_335),
.A2(n_268),
.B(n_251),
.C(n_239),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_336),
.B(n_239),
.Y(n_402)
);

NAND2x1p5_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_271),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_336),
.B(n_271),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_252),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_354),
.B(n_351),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_271),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_366),
.A2(n_167),
.B1(n_188),
.B2(n_192),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_341),
.B(n_193),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_340),
.B(n_202),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_252),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_339),
.B(n_205),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_330),
.A2(n_212),
.B(n_88),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_312),
.A2(n_87),
.B(n_151),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_312),
.A2(n_86),
.B(n_150),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_319),
.A2(n_85),
.B(n_149),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_358),
.A2(n_356),
.B(n_343),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_345),
.A2(n_360),
.B(n_367),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_309),
.B(n_30),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_365),
.A2(n_84),
.B(n_147),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_315),
.A2(n_83),
.B(n_145),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_347),
.B(n_364),
.Y(n_429)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_359),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_323),
.B(n_353),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_362),
.A2(n_90),
.B(n_144),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_348),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_331),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_357),
.A2(n_91),
.B(n_143),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_357),
.A2(n_81),
.B(n_142),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_331),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_307),
.B(n_32),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_357),
.A2(n_93),
.B(n_141),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_14),
.C(n_16),
.Y(n_441)
);

NOR3xp33_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_14),
.C(n_16),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_393),
.A2(n_33),
.B(n_34),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_379),
.A2(n_35),
.B(n_36),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_400),
.B(n_37),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_387),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_372),
.A2(n_38),
.B(n_39),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_40),
.B(n_41),
.Y(n_449)
);

OAI21x1_ASAP7_75t_SL g450 ( 
.A1(n_427),
.A2(n_42),
.B(n_43),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_46),
.Y(n_451)
);

OA22x2_ASAP7_75t_L g452 ( 
.A1(n_390),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_409),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_424),
.A2(n_51),
.B(n_52),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_378),
.B(n_388),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_423),
.A2(n_54),
.B(n_55),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_402),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_389),
.B(n_57),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_382),
.B(n_61),
.Y(n_460)
);

NAND2x1p5_ASAP7_75t_L g461 ( 
.A(n_410),
.B(n_395),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_380),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_66),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_397),
.A2(n_439),
.B(n_408),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_67),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_68),
.Y(n_469)
);

AOI21xp33_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_69),
.B(n_70),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_377),
.B(n_72),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_73),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_74),
.A3(n_75),
.B(n_76),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_398),
.A2(n_92),
.B(n_94),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_387),
.Y(n_476)
);

AO21x2_ASAP7_75t_L g477 ( 
.A1(n_422),
.A2(n_391),
.B(n_384),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_95),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_373),
.A2(n_155),
.B(n_97),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_376),
.A2(n_139),
.B(n_99),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_374),
.A2(n_96),
.B(n_100),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_411),
.B(n_101),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_375),
.A2(n_104),
.B(n_105),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_410),
.B(n_106),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_401),
.A2(n_107),
.B(n_109),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_381),
.A2(n_138),
.B(n_112),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_110),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_371),
.A2(n_113),
.B(n_115),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_395),
.A2(n_117),
.B(n_118),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_411),
.A2(n_120),
.B(n_121),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_418),
.B(n_122),
.Y(n_492)
);

AOI21x1_ASAP7_75t_SL g493 ( 
.A1(n_425),
.A2(n_123),
.B(n_124),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_410),
.B(n_126),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_127),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_438),
.A2(n_128),
.B(n_133),
.C(n_134),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_399),
.B(n_135),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_428),
.B(n_136),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_392),
.A2(n_394),
.B(n_404),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_403),
.B(n_432),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_462),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_466),
.A2(n_463),
.B(n_488),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_421),
.B(n_420),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_454),
.A2(n_440),
.B(n_437),
.Y(n_505)
);

INVx3_ASAP7_75t_SL g506 ( 
.A(n_476),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_471),
.A2(n_436),
.B(n_417),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_492),
.A2(n_406),
.B(n_426),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_457),
.B(n_433),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_419),
.B(n_433),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_475),
.A2(n_456),
.B(n_493),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_480),
.A2(n_481),
.B(n_489),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_465),
.B(n_453),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_461),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_471),
.A2(n_469),
.B(n_460),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_468),
.A2(n_483),
.B1(n_478),
.B2(n_455),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_467),
.B(n_451),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_464),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_458),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_443),
.A2(n_446),
.B(n_444),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_473),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_450),
.A2(n_444),
.B(n_443),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_497),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_485),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_460),
.A2(n_490),
.B(n_448),
.Y(n_533)
);

AOI22x1_ASAP7_75t_L g534 ( 
.A1(n_486),
.A2(n_484),
.B1(n_491),
.B2(n_449),
.Y(n_534)
);

AO31x2_ASAP7_75t_L g535 ( 
.A1(n_496),
.A2(n_472),
.A3(n_482),
.B(n_470),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_442),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_474),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_470),
.A2(n_484),
.B(n_486),
.Y(n_539)
);

OAI21x1_ASAP7_75t_SL g540 ( 
.A1(n_491),
.A2(n_449),
.B(n_452),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_452),
.A2(n_477),
.B(n_474),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_477),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_424),
.B(n_393),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_468),
.A2(n_483),
.B1(n_331),
.B2(n_322),
.Y(n_546)
);

AO21x1_ASAP7_75t_L g547 ( 
.A1(n_518),
.A2(n_541),
.B(n_525),
.Y(n_547)
);

AOI21xp33_ASAP7_75t_L g548 ( 
.A1(n_546),
.A2(n_529),
.B(n_534),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_513),
.B(n_517),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_520),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_503),
.Y(n_551)
);

BUFx2_ASAP7_75t_SL g552 ( 
.A(n_513),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_530),
.Y(n_553)
);

AO21x1_ASAP7_75t_L g554 ( 
.A1(n_525),
.A2(n_543),
.B(n_526),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_527),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_508),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_545),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_511),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_521),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_524),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_546),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_502),
.A2(n_526),
.B(n_540),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_514),
.A2(n_515),
.B(n_544),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_517),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_501),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_538),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_509),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_511),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_519),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_522),
.B(n_523),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_519),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_519),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_515),
.A2(n_507),
.B(n_514),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_506),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_512),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_531),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_500),
.A2(n_504),
.B(n_505),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_531),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_539),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_523),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_566),
.B(n_542),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_557),
.B(n_542),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_553),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_572),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_536),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_533),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_569),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_559),
.B(n_539),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_571),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_556),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_562),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_559),
.B(n_539),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_573),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_583),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_579),
.B(n_528),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_560),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_550),
.B(n_506),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_561),
.B(n_535),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_550),
.B(n_535),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_565),
.B(n_535),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_549),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_547),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_565),
.B(n_535),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_563),
.B(n_505),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_585),
.B(n_501),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_548),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_587),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_587),
.B(n_570),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_551),
.B(n_555),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_547),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_567),
.B(n_554),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_571),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_576),
.B(n_569),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_554),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_576),
.B(n_569),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_576),
.A2(n_549),
.B1(n_578),
.B2(n_577),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_576),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_597),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_600),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_584),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_582),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_622),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_622),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_604),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_591),
.B(n_607),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_611),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_589),
.B(n_582),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_608),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_591),
.A2(n_576),
.B1(n_571),
.B2(n_581),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_589),
.B(n_582),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_608),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_580),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_632),
.B(n_575),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_612),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_612),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_SL g654 ( 
.A(n_621),
.B(n_552),
.Y(n_654)
);

OR2x6_ASAP7_75t_SL g655 ( 
.A(n_607),
.B(n_552),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_595),
.B(n_549),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_594),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_613),
.B(n_568),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_575),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_593),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_592),
.A2(n_575),
.B1(n_586),
.B2(n_568),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_610),
.B(n_618),
.Y(n_664)
);

NOR2x1_ASAP7_75t_L g665 ( 
.A(n_599),
.B(n_629),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_606),
.A2(n_609),
.B1(n_601),
.B2(n_615),
.C(n_630),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_603),
.Y(n_667)
);

AND2x4_ASAP7_75t_SL g668 ( 
.A(n_620),
.B(n_632),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_625),
.B(n_588),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_588),
.B(n_628),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_610),
.B(n_614),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_621),
.B(n_628),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_670),
.B(n_627),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_657),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_651),
.B(n_596),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_638),
.B(n_626),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_638),
.B(n_626),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_643),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_657),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_669),
.B(n_627),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

NAND4xp25_ASAP7_75t_L g685 ( 
.A(n_666),
.B(n_617),
.C(n_629),
.D(n_599),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_661),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_662),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_645),
.B(n_617),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_614),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_665),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_658),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_636),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_648),
.B(n_602),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_674),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_658),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_664),
.B(n_602),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_642),
.B(n_611),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_664),
.B(n_598),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_673),
.B(n_631),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_667),
.Y(n_700)
);

AND2x4_ASAP7_75t_SL g701 ( 
.A(n_635),
.B(n_620),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_641),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_693),
.B(n_689),
.Y(n_703)
);

INVx3_ASAP7_75t_SL g704 ( 
.A(n_690),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_693),
.B(n_689),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_691),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_694),
.B(n_637),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_700),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_697),
.B(n_620),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_686),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_676),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_687),
.B(n_637),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_677),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_692),
.B(n_656),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_677),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_682),
.B(n_659),
.Y(n_716)
);

NOR2x1p5_ASAP7_75t_L g717 ( 
.A(n_685),
.B(n_599),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_676),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_681),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_713),
.Y(n_720)
);

AOI33xp33_ASAP7_75t_L g721 ( 
.A1(n_708),
.A2(n_647),
.A3(n_679),
.B1(n_678),
.B2(n_688),
.B3(n_699),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_620),
.B1(n_677),
.B2(n_710),
.Y(n_722)
);

AOI21xp33_ASAP7_75t_L g723 ( 
.A1(n_714),
.A2(n_690),
.B(n_683),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_711),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_718),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_703),
.B(n_698),
.Y(n_726)
);

OAI221xp5_ASAP7_75t_L g727 ( 
.A1(n_704),
.A2(n_647),
.B1(n_629),
.B2(n_707),
.C(n_712),
.Y(n_727)
);

AOI32xp33_ASAP7_75t_L g728 ( 
.A1(n_703),
.A2(n_699),
.A3(n_679),
.B1(n_678),
.B2(n_688),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_716),
.A2(n_655),
.B1(n_668),
.B2(n_701),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_706),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_724),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_722),
.A2(n_655),
.B1(n_704),
.B2(n_713),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_725),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_720),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_729),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_733),
.B(n_727),
.Y(n_737)
);

AOI221xp5_ASAP7_75t_L g738 ( 
.A1(n_732),
.A2(n_723),
.B1(n_727),
.B2(n_728),
.C(n_730),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_736),
.A2(n_723),
.B(n_633),
.Y(n_739)
);

AOI221xp5_ASAP7_75t_L g740 ( 
.A1(n_734),
.A2(n_731),
.B1(n_680),
.B2(n_654),
.C(n_726),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_737),
.B(n_721),
.C(n_663),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_739),
.B(n_720),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_738),
.B(n_705),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_742),
.Y(n_744)
);

OAI21xp33_ASAP7_75t_L g745 ( 
.A1(n_743),
.A2(n_740),
.B(n_682),
.Y(n_745)
);

NAND4xp75_ASAP7_75t_L g746 ( 
.A(n_744),
.B(n_741),
.C(n_624),
.D(n_623),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_745),
.A2(n_668),
.B1(n_715),
.B2(n_713),
.Y(n_747)
);

NOR4xp25_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_735),
.C(n_597),
.D(n_706),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_746),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_747),
.Y(n_750)
);

NAND4xp75_ASAP7_75t_L g751 ( 
.A(n_748),
.B(n_624),
.C(n_705),
.D(n_623),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_747),
.B(n_735),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_746),
.Y(n_753)
);

XNOR2xp5_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_654),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

XNOR2x1_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_715),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_752),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_753),
.Y(n_758)
);

XNOR2x1_ASAP7_75t_L g759 ( 
.A(n_753),
.B(n_715),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_754),
.B(n_716),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_757),
.B(n_751),
.Y(n_761)
);

AND4x1_ASAP7_75t_L g762 ( 
.A(n_758),
.B(n_709),
.C(n_663),
.D(n_631),
.Y(n_762)
);

AOI22x1_ASAP7_75t_L g763 ( 
.A1(n_755),
.A2(n_634),
.B1(n_597),
.B2(n_684),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_760),
.A2(n_759),
.B1(n_756),
.B2(n_684),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_758),
.B(n_696),
.Y(n_765)
);

XNOR2xp5_ASAP7_75t_L g766 ( 
.A(n_756),
.B(n_701),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_R g767 ( 
.A(n_761),
.B(n_684),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_675),
.B1(n_695),
.B2(n_681),
.Y(n_768)
);

AO22x1_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_702),
.B1(n_650),
.B2(n_635),
.Y(n_769)
);

AOI21xp33_ASAP7_75t_L g770 ( 
.A1(n_764),
.A2(n_763),
.B(n_762),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_764),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_765),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_765),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_765),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_765),
.Y(n_775)
);

AO22x2_ASAP7_75t_L g776 ( 
.A1(n_771),
.A2(n_650),
.B1(n_695),
.B2(n_691),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_772),
.A2(n_675),
.B1(n_672),
.B2(n_671),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_773),
.A2(n_650),
.B(n_698),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_767),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_774),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_775),
.A2(n_660),
.B1(n_651),
.B2(n_596),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_768),
.A2(n_644),
.B1(n_652),
.B2(n_653),
.Y(n_782)
);

AOI21xp33_ASAP7_75t_L g783 ( 
.A1(n_770),
.A2(n_596),
.B(n_639),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_780),
.A2(n_769),
.B(n_596),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_779),
.A2(n_619),
.B(n_640),
.Y(n_785)
);

AO21x2_ASAP7_75t_L g786 ( 
.A1(n_783),
.A2(n_605),
.B(n_616),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_778),
.A2(n_651),
.B1(n_660),
.B2(n_616),
.Y(n_787)
);

OA22x2_ASAP7_75t_L g788 ( 
.A1(n_781),
.A2(n_646),
.B1(n_649),
.B2(n_641),
.Y(n_788)
);

AND3x1_ASAP7_75t_L g789 ( 
.A(n_784),
.B(n_785),
.C(n_787),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_SL g790 ( 
.A1(n_788),
.A2(n_776),
.B(n_782),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_789),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_791),
.B(n_790),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_792),
.A2(n_786),
.B1(n_777),
.B2(n_660),
.Y(n_793)
);


endmodule