module real_jpeg_15284_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_0),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_0),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_1),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_2),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_3),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_3),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_145),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_4),
.A2(n_9),
.B1(n_37),
.B2(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_4),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_4),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_4),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_4),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_5),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_5),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_5),
.B(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_5),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_5),
.B(n_354),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

NAND2x1p5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_39),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_7),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_69),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_7),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_7),
.B(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_9),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_10),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_10),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_11),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_11),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_11),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_11),
.B(n_89),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_11),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_11),
.B(n_340),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_215),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_R g17 ( 
.A(n_18),
.B(n_212),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_163),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_19),
.B(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_96),
.C(n_136),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_20),
.A2(n_21),
.B1(n_97),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_60),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_22),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.C(n_45),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_23),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_28),
.C(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_30),
.Y(n_357)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_32),
.B(n_194),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_34),
.B(n_194),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_35),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_378)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_36),
.A2(n_255),
.B(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_42),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_44),
.Y(n_259)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_56),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_47),
.B(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_49),
.Y(n_338)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_50),
.Y(n_284)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_50),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_51),
.B(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_59),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_73),
.B1(n_94),
.B2(n_95),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_71),
.B2(n_72),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_70),
.C(n_72),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_69),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_69),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_78),
.B(n_80),
.C(n_91),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_78),
.B1(n_92),
.B2(n_93),
.Y(n_162)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_80),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_88),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_81),
.A2(n_88),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_81),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_84),
.B(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_88),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_88),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_97),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_122),
.C(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_99),
.B(n_104),
.C(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_109),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_122),
.B1(n_134),
.B2(n_135),
.Y(n_110)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_116),
.C(n_121),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_113),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_113),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_116),
.A2(n_117),
.B1(n_142),
.B2(n_143),
.Y(n_230)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_120),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_120),
.A2(n_121),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_120),
.B(n_283),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_121),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.C(n_132),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_132),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_127),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_129),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_136),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_155),
.C(n_160),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_137),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_147),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_138),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_140),
.A2(n_141),
.B1(n_147),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_146),
.Y(n_342)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_148),
.A2(n_154),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_153),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_156),
.B(n_161),
.Y(n_375)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_187),
.B1(n_210),
.B2(n_211),
.Y(n_168)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_186),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_185),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_175),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_198),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_209),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_R g215 ( 
.A1(n_216),
.A2(n_370),
.B(n_385),
.Y(n_215)
);

OAI21x1_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_285),
.B(n_369),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_269),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_218),
.B(n_269),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_243),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_220),
.B(n_225),
.C(n_243),
.Y(n_372)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.C(n_231),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_231),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_239),
.Y(n_317)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_236),
.B(n_317),
.Y(n_316)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_244),
.B(n_254),
.C(n_265),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.C(n_249),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_270),
.A2(n_271),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_273),
.B(n_275),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.C(n_282),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_282),
.B(n_319),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_363),
.B(n_368),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_321),
.B(n_362),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_313),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_288),
.B(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_304),
.C(n_311),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_289),
.A2(n_290),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_297),
.C(n_300),
.Y(n_315)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_304),
.A2(n_311),
.B1(n_312),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_324)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_316),
.C(n_318),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_332),
.B(n_361),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_323),
.B(n_328),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.C(n_327),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_327),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_329),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_346),
.B(n_360),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_343),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_334),
.B(n_343),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_339),
.Y(n_351)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_352),
.B(n_359),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_348),
.B(n_351),
.Y(n_359)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_358),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_365),
.Y(n_368)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_380),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_373),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_377),
.C(n_379),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_382),
.Y(n_387)
);


endmodule