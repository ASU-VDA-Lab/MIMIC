module real_aes_6656_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_0), .A2(n_177), .B(n_180), .C(n_184), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_1), .B(n_168), .Y(n_187) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_3), .B(n_178), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_4), .A2(n_141), .B(n_144), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_136), .B(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_6), .A2(n_136), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_7), .B(n_168), .Y(n_553) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_8), .A2(n_170), .B(n_242), .Y(n_241) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_9), .A2(n_457), .B1(n_744), .B2(n_745), .C1(n_748), .C2(n_751), .Y(n_456) );
AND2x6_ASAP7_75t_L g141 ( .A(n_10), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_11), .A2(n_141), .B(n_144), .C(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g513 ( .A(n_12), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_13), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_13), .B(n_40), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_14), .B(n_183), .Y(n_524) );
INVx1_ASAP7_75t_L g162 ( .A(n_15), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_16), .B(n_178), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_17), .B(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_18), .A2(n_179), .B(n_533), .C(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_19), .B(n_168), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_20), .B(n_156), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_21), .A2(n_144), .B(n_147), .C(n_155), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_22), .A2(n_182), .B(n_250), .C(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_23), .B(n_183), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_24), .B(n_183), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_25), .Y(n_494) );
INVx1_ASAP7_75t_L g474 ( .A(n_26), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_27), .A2(n_144), .B(n_155), .C(n_245), .Y(n_244) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_29), .Y(n_520) );
INVx1_ASAP7_75t_L g488 ( .A(n_30), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_31), .A2(n_136), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_33), .A2(n_194), .B(n_195), .C(n_199), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_34), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_35), .A2(n_182), .B(n_550), .C(n_552), .Y(n_549) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_37), .B(n_247), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_38), .A2(n_144), .B(n_155), .C(n_473), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g548 ( .A(n_39), .Y(n_548) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_184), .B(n_511), .C(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_42), .B(n_135), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_43), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_44), .B(n_178), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_45), .B(n_136), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_46), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_48), .A2(n_194), .B(n_199), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g181 ( .A(n_49), .Y(n_181) );
INVx1_ASAP7_75t_L g225 ( .A(n_50), .Y(n_225) );
INVx1_ASAP7_75t_L g561 ( .A(n_51), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_52), .A2(n_102), .B1(n_112), .B2(n_755), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_53), .B(n_136), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_54), .Y(n_164) );
CKINVDCx14_ASAP7_75t_R g509 ( .A(n_55), .Y(n_509) );
INVx1_ASAP7_75t_L g142 ( .A(n_56), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_57), .B(n_136), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_58), .B(n_168), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_59), .A2(n_154), .B(n_210), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g161 ( .A(n_60), .Y(n_161) );
INVx1_ASAP7_75t_SL g551 ( .A(n_61), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_62), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_63), .B(n_178), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_64), .B(n_168), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_65), .B(n_179), .Y(n_260) );
INVx1_ASAP7_75t_L g497 ( .A(n_66), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_67), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_68), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_69), .A2(n_144), .B(n_199), .C(n_208), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_70), .Y(n_234) );
INVx1_ASAP7_75t_L g109 ( .A(n_71), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_72), .A2(n_136), .B(n_508), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_73), .A2(n_93), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_73), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_74), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_75), .A2(n_136), .B(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_76), .A2(n_100), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_76), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_77), .A2(n_135), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_78), .Y(n_471) );
INVx1_ASAP7_75t_L g531 ( .A(n_79), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_80), .B(n_152), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_81), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_82), .A2(n_136), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g534 ( .A(n_83), .Y(n_534) );
INVx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g523 ( .A(n_85), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_86), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_87), .B(n_183), .Y(n_261) );
INVx2_ASAP7_75t_L g106 ( .A(n_88), .Y(n_106) );
OR2x2_ASAP7_75t_L g448 ( .A(n_88), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g460 ( .A(n_88), .B(n_450), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_89), .A2(n_144), .B(n_199), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_90), .B(n_136), .Y(n_192) );
INVx1_ASAP7_75t_L g196 ( .A(n_91), .Y(n_196) );
INVxp67_ASAP7_75t_L g237 ( .A(n_92), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_93), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_94), .B(n_170), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_95), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g209 ( .A(n_96), .Y(n_209) );
INVx1_ASAP7_75t_L g256 ( .A(n_97), .Y(n_256) );
INVx2_ASAP7_75t_L g564 ( .A(n_98), .Y(n_564) );
AND2x2_ASAP7_75t_L g227 ( .A(n_99), .B(n_158), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_100), .Y(n_746) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g756 ( .A(n_103), .Y(n_756) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_110), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_106), .C(n_107), .Y(n_104) );
AND2x2_ASAP7_75t_L g450 ( .A(n_105), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g463 ( .A(n_106), .B(n_450), .Y(n_463) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_106), .B(n_449), .Y(n_750) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_455), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g754 ( .A(n_114), .Y(n_754) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_446), .B(n_452), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B1(n_123), .B2(n_124), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_123), .A2(n_458), .B1(n_461), .B2(n_464), .Y(n_457) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_124), .A2(n_458), .B1(n_752), .B2(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_401), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_336), .Y(n_125) );
NAND4xp25_ASAP7_75t_SL g126 ( .A(n_127), .B(n_281), .C(n_305), .D(n_328), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_218), .B1(n_252), .B2(n_265), .C(n_268), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_188), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_130), .A2(n_166), .B1(n_219), .B2(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_130), .B(n_189), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_130), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_130), .B(n_342), .Y(n_428) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
AND2x2_ASAP7_75t_L g296 ( .A(n_131), .B(n_189), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_131), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g319 ( .A(n_131), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g324 ( .A(n_131), .B(n_167), .Y(n_324) );
INVx2_ASAP7_75t_L g356 ( .A(n_131), .Y(n_356) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_131), .Y(n_400) );
AND2x2_ASAP7_75t_L g417 ( .A(n_131), .B(n_294), .Y(n_417) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g335 ( .A(n_132), .B(n_294), .Y(n_335) );
AND2x4_ASAP7_75t_L g349 ( .A(n_132), .B(n_166), .Y(n_349) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_132), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_132), .B(n_288), .Y(n_373) );
AND2x2_ASAP7_75t_L g423 ( .A(n_132), .B(n_190), .Y(n_423) );
AND2x2_ASAP7_75t_L g433 ( .A(n_132), .B(n_167), .Y(n_433) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_163), .Y(n_132) );
AOI21xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_143), .B(n_156), .Y(n_133) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_137), .B(n_141), .Y(n_257) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g251 ( .A(n_139), .Y(n_251) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx3_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx1_ASAP7_75t_L g247 ( .A(n_140), .Y(n_247) );
BUFx3_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
INVx4_ASAP7_75t_SL g186 ( .A(n_141), .Y(n_186) );
INVx5_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_153), .Y(n_147) );
INVx2_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_152), .A2(n_196), .B(n_197), .C(n_198), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_152), .A2(n_198), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_152), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_499), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_153), .A2(n_178), .B(n_474), .C(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_154), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_157), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_158), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_158), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_158), .A2(n_257), .B(n_471), .C(n_472), .Y(n_470) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_158), .A2(n_507), .B(n_514), .Y(n_506) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g171 ( .A(n_159), .B(n_160), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_165), .A2(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g289 ( .A(n_166), .B(n_189), .Y(n_289) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_166), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_166), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g379 ( .A(n_166), .Y(n_379) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g267 ( .A(n_167), .B(n_204), .Y(n_267) );
AND2x2_ASAP7_75t_L g294 ( .A(n_167), .B(n_205), .Y(n_294) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_187), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_169), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_169), .A2(n_206), .B(n_216), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_169), .B(n_217), .Y(n_216) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_169), .A2(n_255), .B(n_262), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_169), .B(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_169), .A2(n_493), .B(n_500), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_169), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_170), .A2(n_243), .B(n_244), .Y(n_242) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g264 ( .A(n_171), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_186), .Y(n_173) );
INVx2_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_175), .A2(n_186), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_175), .A2(n_186), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_175), .A2(n_186), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_175), .A2(n_186), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_175), .A2(n_186), .B(n_548), .C(n_549), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_SL g560 ( .A1(n_175), .A2(n_186), .B(n_561), .C(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_178), .B(n_237), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_178), .A2(n_211), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_179), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_182), .B(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g511 ( .A(n_183), .Y(n_511) );
INVx2_ASAP7_75t_L g499 ( .A(n_184), .Y(n_499) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_185), .Y(n_198) );
INVx1_ASAP7_75t_L g535 ( .A(n_185), .Y(n_535) );
INVx1_ASAP7_75t_L g199 ( .A(n_186), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_188), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_202), .Y(n_188) );
OR2x2_ASAP7_75t_L g320 ( .A(n_189), .B(n_203), .Y(n_320) );
AND2x2_ASAP7_75t_L g357 ( .A(n_189), .B(n_267), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_189), .B(n_288), .Y(n_368) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_189), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_189), .B(n_324), .Y(n_441) );
INVx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
AND2x2_ASAP7_75t_L g275 ( .A(n_190), .B(n_203), .Y(n_275) );
AND2x2_ASAP7_75t_L g391 ( .A(n_190), .B(n_286), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_190), .B(n_324), .Y(n_413) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_203), .Y(n_359) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_204), .Y(n_311) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g288 ( .A(n_205), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_212), .C(n_213), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_211), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_211), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g552 ( .A(n_214), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_219), .B(n_301), .Y(n_420) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_220), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g272 ( .A(n_220), .B(n_273), .Y(n_272) );
INVx5_ASAP7_75t_SL g280 ( .A(n_220), .Y(n_280) );
OR2x2_ASAP7_75t_L g303 ( .A(n_220), .B(n_273), .Y(n_303) );
OR2x2_ASAP7_75t_L g313 ( .A(n_220), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g376 ( .A(n_220), .B(n_230), .Y(n_376) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_220), .B(n_229), .Y(n_414) );
NOR4xp25_ASAP7_75t_L g435 ( .A(n_220), .B(n_356), .C(n_436), .D(n_437), .Y(n_435) );
AND2x2_ASAP7_75t_L g445 ( .A(n_220), .B(n_277), .Y(n_445) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g270 ( .A(n_229), .B(n_266), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_229), .B(n_272), .Y(n_439) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_239), .Y(n_229) );
OR2x2_ASAP7_75t_L g279 ( .A(n_230), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g286 ( .A(n_230), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_230), .B(n_254), .Y(n_298) );
INVxp67_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_230), .B(n_273), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_230), .B(n_240), .Y(n_367) );
AND2x2_ASAP7_75t_L g382 ( .A(n_230), .B(n_277), .Y(n_382) );
OR2x2_ASAP7_75t_L g411 ( .A(n_230), .B(n_240), .Y(n_411) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_238), .Y(n_230) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_231), .A2(n_529), .B(n_536), .Y(n_528) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_231), .A2(n_546), .B(n_553), .Y(n_545) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_231), .A2(n_559), .B(n_565), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_239), .B(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_239), .B(n_280), .Y(n_419) );
OR2x2_ASAP7_75t_L g440 ( .A(n_239), .B(n_317), .Y(n_440) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g253 ( .A(n_240), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g277 ( .A(n_240), .B(n_273), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_240), .B(n_254), .Y(n_292) );
AND2x2_ASAP7_75t_L g362 ( .A(n_240), .B(n_286), .Y(n_362) );
AND2x2_ASAP7_75t_L g396 ( .A(n_240), .B(n_280), .Y(n_396) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_241), .B(n_280), .Y(n_299) );
AND2x2_ASAP7_75t_L g327 ( .A(n_241), .B(n_254), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_248), .B(n_249), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_249), .A2(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_252), .B(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_253), .A2(n_342), .B1(n_378), .B2(n_395), .C(n_397), .Y(n_394) );
INVx5_ASAP7_75t_SL g273 ( .A(n_254), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_258), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_257), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_257), .A2(n_520), .B(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g482 ( .A(n_264), .Y(n_482) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OAI33xp33_ASAP7_75t_L g293 ( .A1(n_266), .A2(n_294), .A3(n_295), .B1(n_297), .B2(n_300), .B3(n_304), .Y(n_293) );
OR2x2_ASAP7_75t_L g309 ( .A(n_266), .B(n_310), .Y(n_309) );
AOI322xp5_ASAP7_75t_L g418 ( .A1(n_266), .A2(n_335), .A3(n_342), .B1(n_419), .B2(n_420), .C1(n_421), .C2(n_424), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_266), .B(n_294), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_SL g442 ( .A1(n_266), .A2(n_294), .B(n_443), .C(n_445), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_267), .A2(n_282), .B1(n_287), .B2(n_290), .C(n_293), .Y(n_281) );
INVx1_ASAP7_75t_L g374 ( .A(n_267), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_267), .B(n_423), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B1(n_274), .B2(n_276), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g351 ( .A(n_272), .B(n_286), .Y(n_351) );
AND2x2_ASAP7_75t_L g409 ( .A(n_272), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_280), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_273), .B(n_286), .Y(n_345) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_275), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_275), .B(n_353), .Y(n_407) );
OAI321xp33_ASAP7_75t_L g426 ( .A1(n_275), .A2(n_348), .A3(n_427), .B1(n_428), .B2(n_429), .C(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g393 ( .A(n_276), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_277), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g332 ( .A(n_277), .B(n_280), .Y(n_332) );
AOI321xp33_ASAP7_75t_L g390 ( .A1(n_277), .A2(n_294), .A3(n_391), .B1(n_392), .B2(n_393), .C(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g307 ( .A(n_279), .B(n_292), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_280), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_280), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_280), .B(n_366), .Y(n_403) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g326 ( .A(n_284), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g291 ( .A(n_285), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g399 ( .A(n_286), .Y(n_399) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_296), .B(n_331), .Y(n_380) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g344 ( .A(n_299), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g389 ( .A(n_299), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g444 ( .A(n_303), .B(n_367), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B1(n_312), .B2(n_318), .C(n_321), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_SL g388 ( .A(n_314), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_316), .B(n_366), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_316), .A2(n_384), .B(n_386), .Y(n_383) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g429 ( .A(n_317), .B(n_411), .Y(n_429) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g331 ( .A(n_320), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g375 ( .A(n_327), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g437 ( .A(n_327), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B(n_333), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_331), .B(n_349), .Y(n_385) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g406 ( .A(n_335), .Y(n_406) );
NAND5xp2_ASAP7_75t_L g336 ( .A(n_337), .B(n_354), .C(n_363), .D(n_383), .E(n_390), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_343), .C(n_346), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g378 ( .A(n_342), .Y(n_378) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_350), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_358), .B(n_360), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_355), .A2(n_409), .B1(n_412), .B2(n_414), .C(n_415), .Y(n_408) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AOI321xp33_ASAP7_75t_L g363 ( .A1(n_356), .A2(n_364), .A3(n_368), .B1(n_369), .B2(n_375), .C(n_377), .Y(n_363) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g434 ( .A(n_368), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g386 ( .A(n_371), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NOR2xp67_ASAP7_75t_SL g398 ( .A(n_372), .B(n_379), .Y(n_398) );
AOI321xp33_ASAP7_75t_SL g430 ( .A1(n_375), .A2(n_431), .A3(n_432), .B1(n_433), .B2(n_434), .C(n_435), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_380), .C(n_381), .Y(n_377) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_388), .B(n_396), .Y(n_425) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .C(n_400), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_426), .C(n_438), .Y(n_401) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B(n_408), .C(n_418), .Y(n_402) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_407), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_439), .B1(n_440), .B2(n_441), .C(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g431 ( .A(n_429), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g454 ( .A(n_448), .Y(n_454) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_452), .A2(n_456), .B(n_754), .Y(n_455) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g753 ( .A(n_462), .Y(n_753) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g752 ( .A(n_464), .Y(n_752) );
OR4x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_634), .C(n_681), .D(n_721), .Y(n_464) );
NAND3xp33_ASAP7_75t_SL g465 ( .A(n_466), .B(n_580), .C(n_609), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_502), .B(n_537), .C(n_573), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_467), .A2(n_593), .B(n_610), .C(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_469), .B(n_572), .Y(n_571) );
INVx3_ASAP7_75t_SL g576 ( .A(n_469), .Y(n_576) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_469), .Y(n_588) );
AND2x4_ASAP7_75t_L g592 ( .A(n_469), .B(n_544), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_469), .B(n_492), .Y(n_603) );
OR2x2_ASAP7_75t_L g627 ( .A(n_469), .B(n_540), .Y(n_627) );
AND2x2_ASAP7_75t_L g640 ( .A(n_469), .B(n_545), .Y(n_640) );
AND2x2_ASAP7_75t_L g680 ( .A(n_469), .B(n_666), .Y(n_680) );
AND2x2_ASAP7_75t_L g687 ( .A(n_469), .B(n_650), .Y(n_687) );
AND2x2_ASAP7_75t_L g717 ( .A(n_469), .B(n_479), .Y(n_717) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_478), .B(n_644), .Y(n_656) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_479), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g594 ( .A(n_479), .B(n_491), .Y(n_594) );
BUFx3_ASAP7_75t_L g602 ( .A(n_479), .Y(n_602) );
OR2x2_ASAP7_75t_L g623 ( .A(n_479), .B(n_505), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_479), .B(n_644), .Y(n_734) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_481), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_490), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_491), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g587 ( .A(n_491), .Y(n_587) );
AND2x2_ASAP7_75t_L g650 ( .A(n_491), .B(n_545), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_491), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_652) );
AND2x2_ASAP7_75t_L g666 ( .A(n_491), .B(n_540), .Y(n_666) );
AND2x2_ASAP7_75t_L g692 ( .A(n_491), .B(n_576), .Y(n_692) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g572 ( .A(n_492), .B(n_545), .Y(n_572) );
BUFx2_ASAP7_75t_L g706 ( .A(n_492), .Y(n_706) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI32xp33_ASAP7_75t_L g672 ( .A1(n_503), .A2(n_633), .A3(n_647), .B1(n_673), .B2(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
AND2x2_ASAP7_75t_L g613 ( .A(n_504), .B(n_557), .Y(n_613) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_505), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g667 ( .A(n_505), .B(n_557), .Y(n_667) );
AND2x2_ASAP7_75t_L g678 ( .A(n_505), .B(n_570), .Y(n_678) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g579 ( .A(n_506), .B(n_558), .Y(n_579) );
AND2x2_ASAP7_75t_L g583 ( .A(n_506), .B(n_558), .Y(n_583) );
AND2x2_ASAP7_75t_L g618 ( .A(n_506), .B(n_569), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_506), .B(n_527), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_506), .A2(n_576), .B(n_587), .C(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g684 ( .A(n_506), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_506), .B(n_517), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_515), .B(n_567), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_515), .B(n_583), .Y(n_673) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g578 ( .A(n_516), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
AND2x2_ASAP7_75t_L g570 ( .A(n_517), .B(n_528), .Y(n_570) );
OR2x2_ASAP7_75t_L g585 ( .A(n_517), .B(n_528), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_517), .B(n_569), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_517), .Y(n_612) );
AND2x2_ASAP7_75t_L g631 ( .A(n_517), .B(n_568), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_517), .A2(n_596), .B1(n_642), .B2(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_517), .B(n_684), .Y(n_708) );
AND2x2_ASAP7_75t_L g723 ( .A(n_517), .B(n_583), .Y(n_723) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g555 ( .A(n_518), .Y(n_555) );
AND2x2_ASAP7_75t_L g597 ( .A(n_518), .B(n_528), .Y(n_597) );
AND2x2_ASAP7_75t_L g599 ( .A(n_518), .B(n_557), .Y(n_599) );
AND3x2_ASAP7_75t_L g661 ( .A(n_518), .B(n_625), .C(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g696 ( .A(n_527), .B(n_568), .Y(n_696) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_528), .B(n_567), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_528), .B(n_608), .C(n_684), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_554), .B1(n_566), .B2(n_571), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_540), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g648 ( .A(n_540), .Y(n_648) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_543), .A2(n_665), .A3(n_666), .B(n_667), .Y(n_664) );
AND2x2_ASAP7_75t_L g689 ( .A(n_543), .B(n_576), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_543), .B(n_602), .Y(n_735) );
AND2x2_ASAP7_75t_L g644 ( .A(n_544), .B(n_576), .Y(n_644) );
AND2x2_ASAP7_75t_L g705 ( .A(n_544), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g575 ( .A(n_545), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g633 ( .A(n_545), .Y(n_633) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g654 ( .A(n_555), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_556), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AOI221x1_ASAP7_75t_SL g621 ( .A1(n_557), .A2(n_622), .B1(n_624), .B2(n_626), .C(n_628), .Y(n_621) );
INVx2_ASAP7_75t_L g569 ( .A(n_558), .Y(n_569) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
INVx1_ASAP7_75t_L g651 ( .A(n_566), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_567), .B(n_584), .Y(n_676) );
INVx1_ASAP7_75t_SL g739 ( .A(n_567), .Y(n_739) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g657 ( .A(n_570), .B(n_583), .Y(n_657) );
INVx1_ASAP7_75t_L g725 ( .A(n_571), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_571), .B(n_654), .Y(n_738) );
INVx2_ASAP7_75t_SL g577 ( .A(n_572), .Y(n_577) );
AND2x2_ASAP7_75t_L g620 ( .A(n_572), .B(n_576), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_572), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_572), .B(n_647), .Y(n_674) );
AOI21xp33_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_577), .B(n_578), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_575), .B(n_647), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_575), .B(n_602), .Y(n_743) );
OR2x2_ASAP7_75t_L g615 ( .A(n_576), .B(n_594), .Y(n_615) );
AND2x2_ASAP7_75t_L g714 ( .A(n_576), .B(n_705), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_577), .A2(n_590), .B1(n_595), .B2(n_598), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_577), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g637 ( .A(n_579), .B(n_585), .Y(n_637) );
INVx1_ASAP7_75t_L g701 ( .A(n_579), .Y(n_701) );
AOI311xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_586), .A3(n_588), .B(n_589), .C(n_600), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_584), .A2(n_716), .B1(n_728), .B2(n_731), .C(n_733), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_584), .B(n_739), .Y(n_741) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g638 ( .A(n_586), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_629), .B(n_630), .C(n_632), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_591), .A2(n_593), .B(n_698), .C(n_699), .Y(n_697) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_592), .B(n_666), .Y(n_732) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_595), .A2(n_615), .B1(n_616), .B2(n_619), .C(n_621), .Y(n_614) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g617 ( .A(n_597), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g700 ( .A(n_597), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_601), .A2(n_659), .B(n_660), .C(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_602), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_602), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g624 ( .A(n_608), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_612), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g726 ( .A(n_615), .Y(n_726) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_618), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g653 ( .A(n_618), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g730 ( .A(n_618), .Y(n_730) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g671 ( .A(n_620), .B(n_647), .Y(n_671) );
INVx1_ASAP7_75t_SL g665 ( .A(n_627), .Y(n_665) );
INVx1_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_652), .C(n_668), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .A3(n_639), .B1(n_641), .B2(n_645), .C1(n_649), .C2(n_651), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_636), .A2(n_689), .B(n_690), .C(n_697), .Y(n_688) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_639), .A2(n_660), .B1(n_691), .B2(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g649 ( .A(n_647), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g686 ( .A(n_647), .B(n_687), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_738), .A3(n_739), .B1(n_740), .B2(n_742), .Y(n_737) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g659 ( .A(n_650), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_650), .A2(n_703), .B1(n_707), .B2(n_709), .C(n_712), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_650), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g719 ( .A(n_654), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g729 ( .A(n_654), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g720 ( .A(n_663), .B(n_684), .Y(n_720) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_685), .B(n_688), .C(n_702), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_696), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g711 ( .A(n_708), .Y(n_711) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_718), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_724), .B(n_727), .C(n_737), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
endmodule