module fake_netlist_5_2297_n_3103 (n_137, n_294, n_318, n_380, n_419, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_409, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_3103);

input n_137;
input n_294;
input n_318;
input n_380;
input n_419;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_3103;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_2771;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_3086;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_3036;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_3010;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_3048;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2959;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1749;
wire n_1097;
wire n_696;
wire n_550;
wire n_3101;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_436;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_422;
wire n_475;
wire n_777;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_2915;
wire n_1239;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_2682;
wire n_901;
wire n_553;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_2932;
wire n_2753;
wire n_464;
wire n_2980;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_1585;
wire n_571;
wire n_461;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3025;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_2622;
wire n_1278;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_586;
wire n_838;
wire n_2784;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_1276;
wire n_702;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_931;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_870;
wire n_1481;
wire n_2626;
wire n_3042;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_568;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3003;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_3030;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3075;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_3031;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_457;
wire n_514;
wire n_2093;
wire n_2339;
wire n_2320;
wire n_2038;
wire n_2473;
wire n_1208;
wire n_1045;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3045;
wire n_1870;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_504;
wire n_511;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_513;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_560;
wire n_2288;
wire n_2240;
wire n_2696;
wire n_1351;
wire n_1044;
wire n_2436;
wire n_1205;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_2953;
wire n_824;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_3059;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_1630;
wire n_716;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_531;
wire n_3020;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_1346;
wire n_3053;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_515;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1644;
wire n_1283;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_455;
wire n_2993;
wire n_1719;
wire n_1048;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3041;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1668;
wire n_1301;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_3067;
wire n_1932;
wire n_2755;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_540;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_3099;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_2971;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1998;
wire n_1105;
wire n_1019;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_458;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_2988;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_487;
wire n_3035;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_427;
wire n_1399;
wire n_1991;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_500;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_435;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_2692;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_2184;
wire n_1184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2430;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_3070;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_2748;
wire n_518;
wire n_505;
wire n_2057;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_428;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3017;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_3054;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_3050;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_2957;
wire n_839;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_608;
wire n_1367;
wire n_928;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_2961;
wire n_2702;
wire n_2570;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_2612;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_465;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_3004;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_453;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_3057;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_2938;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_2975;
wire n_438;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1827;
wire n_1180;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g420 ( 
.A(n_202),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_21),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_324),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_144),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_58),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_111),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_23),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_132),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_44),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_58),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_397),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_46),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_203),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_373),
.Y(n_435)
);

BUFx8_ASAP7_75t_SL g436 ( 
.A(n_39),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_200),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_358),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_344),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_75),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_36),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_409),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_141),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_368),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_246),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_31),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_127),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_417),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_89),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_348),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_26),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_13),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_107),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_357),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_294),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_124),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_46),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_53),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_135),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_153),
.Y(n_460)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_116),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_220),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_333),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_263),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_280),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_129),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_364),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_327),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_315),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_241),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_190),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_274),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_189),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_355),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_141),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_70),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_293),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_63),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_232),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_114),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_273),
.Y(n_481)
);

BUFx8_ASAP7_75t_SL g482 ( 
.A(n_262),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_212),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_272),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_212),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_86),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_309),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_345),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_334),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_38),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_361),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_224),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_67),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_319),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_45),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_88),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_171),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_404),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_115),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_220),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_41),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_145),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_36),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_275),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_342),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_148),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_395),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_377),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_140),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_158),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_9),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_28),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_63),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_282),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_103),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_314),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_288),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_351),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_302),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_128),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_250),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_298),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_208),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_130),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_123),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_156),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_388),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_38),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_401),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_73),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_151),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_384),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_230),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_144),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_322),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_97),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_30),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_248),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_150),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_374),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_64),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_89),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_106),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_132),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_249),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_149),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_112),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_60),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_84),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_225),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_283),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_114),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_222),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_347),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_33),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_235),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_161),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_22),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_353),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_140),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_93),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_150),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_74),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_135),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_202),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_224),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_154),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_138),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_271),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_329),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_268),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_238),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_231),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_164),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_71),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_195),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_85),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_120),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_81),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_16),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_332),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_408),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_299),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_174),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_205),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_405),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_162),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_161),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_32),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_331),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_242),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_27),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_20),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_214),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_152),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_413),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_18),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_102),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_29),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_296),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_407),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_326),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_199),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_106),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_69),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_25),
.Y(n_607)
);

INVxp33_ASAP7_75t_R g608 ( 
.A(n_51),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_257),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_138),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_372),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_244),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_68),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_359),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_100),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_68),
.Y(n_616)
);

BUFx5_ASAP7_75t_L g617 ( 
.A(n_143),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_276),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_366),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_34),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_306),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_186),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_108),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_411),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_182),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_60),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_52),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_316),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_0),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_287),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_410),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_360),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_183),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_69),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_349),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_85),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_369),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_166),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_217),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_206),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_318),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_142),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_37),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_330),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_41),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_304),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_211),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_78),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_148),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_156),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_290),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_33),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_13),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_321),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_160),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_102),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_155),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_54),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_402),
.Y(n_659)
);

CKINVDCx16_ASAP7_75t_R g660 ( 
.A(n_62),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_363),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_70),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_163),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_254),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_176),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_34),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_168),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_0),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_365),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_258),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_97),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_107),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_87),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_375),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_157),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_28),
.Y(n_676)
);

BUFx8_ASAP7_75t_SL g677 ( 
.A(n_270),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_25),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_66),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_200),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_199),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_115),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_182),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_35),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_179),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_226),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_92),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_370),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_176),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_312),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_301),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_32),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_169),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_284),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_178),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_399),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_111),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_234),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_267),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_103),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_154),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_82),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_51),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_320),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_184),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_387),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_175),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_256),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_54),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_104),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_48),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_59),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_76),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_247),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_378),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_143),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_216),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_190),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_91),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_305),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_303),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_88),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_341),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_165),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_116),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_264),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_461),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_541),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_461),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_436),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_580),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_461),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_453),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_541),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_461),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_453),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_461),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_461),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_678),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_461),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_461),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_461),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_617),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_546),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_678),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_617),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_617),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_617),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_707),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_617),
.Y(n_751)
);

CKINVDCx16_ASAP7_75t_R g752 ( 
.A(n_660),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_617),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_660),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_451),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_451),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_617),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_451),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_540),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_451),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_451),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_662),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_451),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_546),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_486),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_540),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_486),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_486),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_420),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_420),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_662),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_486),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_486),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_486),
.Y(n_775)
);

BUFx2_ASAP7_75t_SL g776 ( 
.A(n_469),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_496),
.B(n_1),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_463),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_421),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_421),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_481),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_445),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_522),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_445),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_426),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_422),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_470),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_470),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_424),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_472),
.B(n_1),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_426),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_696),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_472),
.Y(n_793)
);

INVxp33_ASAP7_75t_SL g794 ( 
.A(n_427),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_474),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_696),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_429),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_474),
.B(n_2),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_484),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_484),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_494),
.B(n_2),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_699),
.Y(n_802)
);

INVxp33_ASAP7_75t_L g803 ( 
.A(n_434),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_494),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_606),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_606),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_431),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_433),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_498),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_498),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_518),
.Y(n_811)
);

INVxp33_ASAP7_75t_SL g812 ( 
.A(n_437),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_518),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_434),
.Y(n_814)
);

INVxp33_ASAP7_75t_SL g815 ( 
.A(n_441),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_606),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_699),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_519),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_440),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_606),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_519),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_532),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_623),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_532),
.Y(n_824)
);

INVx4_ASAP7_75t_R g825 ( 
.A(n_708),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_533),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_533),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_708),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_552),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_552),
.Y(n_830)
);

INVxp33_ASAP7_75t_SL g831 ( 
.A(n_443),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_440),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_517),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_606),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_570),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_606),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_463),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_522),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_570),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_573),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_573),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_583),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_543),
.Y(n_843)
);

INVxp33_ASAP7_75t_SL g844 ( 
.A(n_447),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_674),
.Y(n_845)
);

INVxp33_ASAP7_75t_L g846 ( 
.A(n_446),
.Y(n_846)
);

INVxp67_ASAP7_75t_SL g847 ( 
.A(n_655),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_456),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_582),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_655),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_655),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_655),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_423),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_655),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_655),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_691),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_462),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_482),
.Y(n_858)
);

INVxp33_ASAP7_75t_SL g859 ( 
.A(n_457),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_462),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_490),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_490),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_512),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_623),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_680),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_512),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_781),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_864),
.B(n_680),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_757),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_778),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_757),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_761),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_778),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_767),
.B(n_602),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_778),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_778),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_792),
.B(n_602),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_736),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_776),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_865),
.B(n_796),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_757),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_802),
.B(n_632),
.Y(n_883)
);

OA21x2_ASAP7_75t_L g884 ( 
.A1(n_759),
.A2(n_854),
.B(n_851),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_730),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_736),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_817),
.B(n_632),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_828),
.B(n_654),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_776),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_805),
.Y(n_890)
);

OA21x2_ASAP7_75t_L g891 ( 
.A1(n_759),
.A2(n_584),
.B(n_582),
.Y(n_891)
);

INVxp33_ASAP7_75t_SL g892 ( 
.A(n_730),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_745),
.A2(n_459),
.B1(n_460),
.B2(n_458),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_778),
.B(n_463),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_834),
.B(n_654),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_762),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_837),
.Y(n_897)
);

CKINVDCx14_ASAP7_75t_R g898 ( 
.A(n_858),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_805),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_837),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_760),
.B(n_510),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_762),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_765),
.B(n_859),
.Y(n_903)
);

BUFx8_ASAP7_75t_L g904 ( 
.A(n_746),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_790),
.B(n_463),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_836),
.B(n_425),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_760),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_837),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_847),
.B(n_432),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_783),
.A2(n_838),
.B1(n_752),
.B2(n_733),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_833),
.Y(n_912)
);

OA21x2_ASAP7_75t_L g913 ( 
.A1(n_764),
.A2(n_601),
.B(n_584),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_766),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_823),
.B(n_510),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_728),
.A2(n_476),
.B1(n_483),
.B2(n_473),
.Y(n_916)
);

CKINVDCx11_ASAP7_75t_R g917 ( 
.A(n_842),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_837),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_845),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_766),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_768),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_768),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_737),
.A2(n_611),
.B(n_601),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_806),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_734),
.A2(n_430),
.B1(n_449),
.B2(n_428),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_806),
.B(n_816),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_769),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_837),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_816),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_843),
.B(n_435),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_769),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_820),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_754),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_820),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_755),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_773),
.A2(n_612),
.B(n_611),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_755),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_754),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_856),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_852),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_852),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_755),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_823),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_737),
.A2(n_618),
.B(n_612),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_739),
.A2(n_485),
.B1(n_495),
.B2(n_493),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_779),
.B(n_618),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_773),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_774),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_438),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_SL g950 ( 
.A1(n_763),
.A2(n_478),
.B1(n_480),
.B2(n_466),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_780),
.Y(n_951)
);

AND2x4_ASAP7_75t_SL g952 ( 
.A(n_782),
.B(n_543),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_853),
.B(n_439),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_794),
.B(n_812),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_774),
.Y(n_955)
);

CKINVDCx16_ASAP7_75t_R g956 ( 
.A(n_746),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_775),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_775),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_786),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_784),
.B(n_630),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_850),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_850),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_851),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_854),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_787),
.B(n_788),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_794),
.B(n_448),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_855),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_793),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_795),
.B(n_630),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_812),
.B(n_555),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_855),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_729),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_815),
.B(n_624),
.Y(n_973)
);

OA21x2_ASAP7_75t_L g974 ( 
.A1(n_729),
.A2(n_646),
.B(n_641),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_732),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_732),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_799),
.B(n_641),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_743),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_770),
.B(n_803),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_727),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_735),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_763),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_731),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_738),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_740),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_772),
.A2(n_509),
.B1(n_530),
.B2(n_524),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_743),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_744),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_744),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_849),
.B(n_442),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_923),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_923),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_966),
.B(n_815),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_906),
.B(n_849),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_979),
.B(n_831),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_944),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_979),
.B(n_831),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_943),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_944),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_873),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_956),
.B(n_772),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_926),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_926),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_975),
.B(n_463),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_926),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_946),
.B(n_646),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_943),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_926),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_975),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_907),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_873),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_976),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_873),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_907),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_976),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_978),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_872),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_978),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_877),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_987),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_987),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_873),
.Y(n_1024)
);

AND2x2_ASAP7_75t_SL g1025 ( 
.A(n_905),
.B(n_974),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_988),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_877),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_956),
.B(n_750),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_946),
.B(n_659),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_SL g1031 ( 
.A(n_905),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_988),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_989),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_901),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_989),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_972),
.Y(n_1036)
);

XNOR2xp5_ASAP7_75t_L g1037 ( 
.A(n_925),
.B(n_547),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_875),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_890),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_875),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_972),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_972),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_899),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_980),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_875),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_899),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_875),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_924),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_980),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_924),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_875),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_990),
.A2(n_742),
.B(n_741),
.Y(n_1052)
);

AND2x2_ASAP7_75t_SL g1053 ( 
.A(n_905),
.B(n_463),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_909),
.B(n_849),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_984),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_984),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_896),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_901),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_934),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_869),
.A2(n_748),
.B(n_747),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_869),
.A2(n_748),
.B(n_747),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_897),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_896),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_902),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_902),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_897),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_897),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_946),
.B(n_659),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_910),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_934),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_940),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_910),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_914),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_940),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_881),
.B(n_800),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_914),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_920),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_920),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_970),
.B(n_844),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_941),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_897),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_921),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_908),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_935),
.B(n_849),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_941),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_955),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_915),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_922),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_922),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_927),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_962),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_927),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_917),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_915),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_962),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_931),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_931),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_948),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_908),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_964),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_948),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_961),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_904),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_967),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_967),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_971),
.Y(n_1109)
);

BUFx8_ASAP7_75t_L g1110 ( 
.A(n_885),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_964),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_971),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_929),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_871),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_929),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_935),
.B(n_849),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_871),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_882),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_908),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_879),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_973),
.B(n_844),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_895),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_886),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_882),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_884),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_881),
.B(n_804),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_933),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_884),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_929),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_868),
.B(n_809),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_965),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_868),
.B(n_810),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_908),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_908),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_965),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_903),
.B(n_859),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_965),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_904),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_929),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_935),
.B(n_849),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_938),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_884),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_884),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_982),
.B(n_786),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_981),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_981),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_929),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_946),
.B(n_811),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_981),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_982),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_981),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_981),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_912),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_952),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_985),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1122),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1122),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1112),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1095),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1053),
.A2(n_974),
.B1(n_913),
.B2(n_936),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1122),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1112),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1128),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1128),
.B(n_960),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1031),
.A2(n_556),
.B1(n_639),
.B2(n_525),
.Y(n_1166)
);

NOR2x1p5_ASAP7_75t_L g1167 ( 
.A(n_1028),
.B(n_731),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1053),
.B(n_952),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1132),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1060),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1053),
.B(n_880),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1010),
.B(n_895),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_993),
.B(n_959),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1132),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1136),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1136),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1138),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1138),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1079),
.A2(n_925),
.B1(n_911),
.B2(n_889),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1001),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1003),
.Y(n_1181)
);

AND2x6_ASAP7_75t_L g1182 ( 
.A(n_1125),
.B(n_664),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1003),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1060),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1004),
.Y(n_1185)
);

AND2x6_ASAP7_75t_L g1186 ( 
.A(n_1125),
.B(n_664),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1025),
.B(n_880),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_998),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1012),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1060),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1001),
.Y(n_1191)
);

AND2x6_ASAP7_75t_L g1192 ( 
.A(n_1125),
.B(n_720),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1028),
.B(n_1002),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1004),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1137),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1001),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1006),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1121),
.B(n_954),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1037),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1006),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_L g1201 ( 
.A(n_995),
.B(n_950),
.C(n_916),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1010),
.B(n_895),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_997),
.B(n_953),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_1155),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1060),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1008),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1014),
.B(n_895),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1061),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1014),
.B(n_942),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1061),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1001),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1009),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_1120),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1031),
.A2(n_974),
.B1(n_913),
.B2(n_936),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1089),
.B(n_930),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1031),
.A2(n_1025),
.B1(n_1129),
.B2(n_1143),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1105),
.B(n_885),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1009),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1114),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1110),
.Y(n_1220)
);

INVx6_ASAP7_75t_L g1221 ( 
.A(n_1110),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1154),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1114),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1149),
.B(n_960),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1117),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1117),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1118),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1016),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1031),
.A2(n_974),
.B1(n_913),
.B2(n_936),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1118),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1149),
.B(n_960),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1025),
.B(n_889),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1155),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1075),
.A2(n_949),
.B1(n_874),
.B2(n_883),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1007),
.B(n_960),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1002),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1061),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1124),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1061),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1096),
.B(n_789),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1124),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1017),
.B(n_942),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1105),
.A2(n_904),
.B1(n_577),
.B2(n_600),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1131),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1034),
.B(n_789),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1058),
.B(n_797),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1011),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1017),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1129),
.A2(n_913),
.B1(n_936),
.B2(n_891),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1075),
.B(n_797),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1057),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1126),
.A2(n_986),
.B1(n_887),
.B2(n_888),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1018),
.B(n_1020),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1131),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1133),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1057),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1001),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1126),
.B(n_807),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1151),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1133),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1018),
.B(n_985),
.Y(n_1261)
);

BUFx10_ASAP7_75t_L g1262 ( 
.A(n_1007),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1063),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1063),
.Y(n_1264)
);

AND2x6_ASAP7_75t_L g1265 ( 
.A(n_1129),
.B(n_720),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1020),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1011),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1022),
.B(n_807),
.Y(n_1268)
);

NOR2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1110),
.B(n_983),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1064),
.Y(n_1270)
);

INVx4_ASAP7_75t_L g1271 ( 
.A(n_1001),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1022),
.A2(n_1023),
.B1(n_1032),
.B2(n_1026),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1007),
.B(n_969),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1023),
.B(n_985),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1026),
.B(n_808),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1085),
.B(n_985),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1064),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1013),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1013),
.Y(n_1279)
);

AO22x2_ASAP7_75t_L g1280 ( 
.A1(n_1007),
.A2(n_556),
.B1(n_639),
.B2(n_525),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1065),
.Y(n_1281)
);

OAI21xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1143),
.A2(n_801),
.B(n_798),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1032),
.B(n_985),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1065),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1069),
.Y(n_1285)
);

AND2x2_ASAP7_75t_SL g1286 ( 
.A(n_1030),
.B(n_721),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1116),
.B(n_937),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1069),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1033),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1033),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1144),
.A2(n_891),
.B1(n_977),
.B2(n_969),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1123),
.B(n_808),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1145),
.B(n_848),
.C(n_893),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1072),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1013),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1146),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1035),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1035),
.B(n_848),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1141),
.B(n_937),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1127),
.B(n_814),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1144),
.A2(n_891),
.B1(n_977),
.B2(n_969),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1036),
.B(n_937),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1072),
.B(n_878),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1005),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_L g1305 ( 
.A(n_1139),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1030),
.A2(n_891),
.B1(n_977),
.B2(n_969),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1073),
.B(n_945),
.Y(n_1307)
);

AND2x6_ASAP7_75t_L g1308 ( 
.A(n_991),
.B(n_726),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1030),
.A2(n_977),
.B1(n_567),
.B2(n_711),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1027),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1073),
.B(n_951),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1030),
.A2(n_690),
.B1(n_670),
.B2(n_651),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1076),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1068),
.A2(n_992),
.B1(n_996),
.B2(n_991),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1076),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1068),
.A2(n_567),
.B1(n_711),
.B2(n_565),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1077),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1077),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1068),
.A2(n_565),
.B1(n_446),
.B2(n_471),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1078),
.B(n_951),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1078),
.B(n_968),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1082),
.Y(n_1322)
);

INVxp33_ASAP7_75t_SL g1323 ( 
.A(n_1037),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1142),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1036),
.B(n_937),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1082),
.B(n_968),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_1139),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1013),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1068),
.B(n_819),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1083),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1083),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1090),
.B(n_892),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1090),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1110),
.B(n_723),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1091),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1091),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1092),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1041),
.B(n_937),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_992),
.A2(n_471),
.B1(n_492),
.B2(n_452),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1041),
.B(n_937),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1013),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1092),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1094),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1094),
.B(n_475),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1042),
.B(n_721),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1098),
.B(n_726),
.Y(n_1346)
);

INVx5_ASAP7_75t_L g1347 ( 
.A(n_1005),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1098),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1099),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1099),
.Y(n_1350)
);

INVx5_ASAP7_75t_L g1351 ( 
.A(n_1005),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1100),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1181),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1300),
.B(n_912),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1244),
.B(n_919),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1221),
.B(n_723),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1244),
.B(n_904),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1185),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1173),
.B(n_986),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1183),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1193),
.B(n_919),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1234),
.B(n_1100),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1255),
.B(n_1260),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1197),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1173),
.B(n_1103),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1200),
.Y(n_1366)
);

AND2x6_ASAP7_75t_L g1367 ( 
.A(n_1170),
.B(n_996),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1222),
.B(n_939),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1259),
.B(n_939),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1212),
.B(n_1103),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1255),
.B(n_1104),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1218),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1240),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1176),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1198),
.B(n_1104),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1198),
.B(n_1106),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1303),
.B(n_1106),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1176),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1216),
.B(n_1042),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1164),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1169),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1160),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_SL g1383 ( 
.A(n_1217),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1189),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1215),
.B(n_1107),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1215),
.B(n_1107),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1185),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1171),
.A2(n_1109),
.B(n_1108),
.C(n_1049),
.Y(n_1388)
);

BUFx8_ASAP7_75t_L g1389 ( 
.A(n_1324),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1260),
.B(n_1108),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_L g1391 ( 
.A(n_1216),
.B(n_1109),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1188),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1206),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1266),
.B(n_994),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1194),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1266),
.B(n_1054),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1297),
.B(n_1044),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1297),
.B(n_1044),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1250),
.B(n_846),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1187),
.A2(n_1147),
.B1(n_1150),
.B2(n_1146),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1330),
.B(n_1049),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1174),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1250),
.B(n_983),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1257),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1258),
.B(n_608),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1282),
.A2(n_1000),
.B1(n_492),
.B2(n_497),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1337),
.B(n_867),
.Y(n_1407)
);

AND2x2_ASAP7_75t_SL g1408 ( 
.A(n_1286),
.B(n_721),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1213),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1330),
.B(n_1055),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1175),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1337),
.B(n_1168),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1258),
.B(n_1147),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1177),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1240),
.B(n_1275),
.C(n_1268),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1350),
.B(n_1055),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1337),
.B(n_1056),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1178),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1254),
.B(n_1203),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1171),
.A2(n_1056),
.B(n_701),
.C(n_1000),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1203),
.B(n_698),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1187),
.A2(n_1150),
.B1(n_1153),
.B2(n_1152),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1194),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1332),
.B(n_1152),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1286),
.B(n_1158),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1158),
.B(n_1153),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1213),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1179),
.A2(n_629),
.B1(n_681),
.B2(n_562),
.C(n_515),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1232),
.A2(n_1156),
.B1(n_1052),
.B2(n_1115),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1350),
.B(n_1156),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1189),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1195),
.B(n_575),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1248),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1332),
.B(n_444),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1195),
.B(n_450),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1352),
.B(n_1148),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1232),
.A2(n_1052),
.B1(n_1115),
.B2(n_1113),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1252),
.A2(n_813),
.B(n_821),
.C(n_818),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1195),
.B(n_581),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1268),
.B(n_454),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1248),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1275),
.B(n_626),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1314),
.A2(n_1130),
.B1(n_1140),
.B2(n_1113),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1257),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1298),
.B(n_455),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1298),
.B(n_464),
.Y(n_1446)
);

NOR2xp67_ASAP7_75t_SL g1447 ( 
.A(n_1304),
.B(n_1347),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1352),
.B(n_1130),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1293),
.B(n_898),
.C(n_692),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1329),
.B(n_465),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1245),
.B(n_663),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1311),
.B(n_1140),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1289),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1246),
.B(n_1344),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1307),
.B(n_1236),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1199),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1289),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_1148),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1290),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1307),
.B(n_777),
.C(n_502),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1326),
.B(n_999),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1290),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1344),
.B(n_675),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1228),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1235),
.B(n_1013),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1201),
.B(n_503),
.C(n_501),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1235),
.B(n_1015),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1326),
.B(n_999),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1224),
.B(n_467),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1251),
.B(n_999),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1292),
.B(n_771),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1256),
.B(n_999),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1220),
.B(n_785),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1263),
.B(n_1038),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1317),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1228),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1339),
.A2(n_832),
.B1(n_791),
.B2(n_499),
.C(n_500),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1335),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1264),
.B(n_1348),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1224),
.B(n_468),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1335),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1336),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1314),
.A2(n_684),
.B1(n_703),
.B2(n_676),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1204),
.B(n_534),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1270),
.B(n_718),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1277),
.B(n_1038),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1224),
.A2(n_1111),
.B(n_1102),
.C(n_824),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1281),
.B(n_1038),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1312),
.B(n_513),
.C(n_511),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1336),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1284),
.B(n_1038),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1235),
.B(n_1015),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1257),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1306),
.A2(n_1111),
.B1(n_1102),
.B2(n_1088),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1339),
.A2(n_497),
.B1(n_499),
.B2(n_452),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1182),
.A2(n_506),
.B1(n_520),
.B2(n_500),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1204),
.B(n_534),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1285),
.B(n_1062),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1199),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1288),
.B(n_1062),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1257),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_SL g1503 ( 
.A(n_1217),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1231),
.A2(n_1066),
.B1(n_1067),
.B2(n_1062),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1365),
.B(n_1349),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1365),
.B(n_1294),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1382),
.Y(n_1507)
);

INVx8_ASAP7_75t_L g1508 ( 
.A(n_1367),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1404),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1384),
.B(n_1231),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1467),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1359),
.A2(n_1231),
.B1(n_1165),
.B2(n_1273),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1404),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1483),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1399),
.B(n_1305),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1404),
.B(n_1273),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1374),
.B(n_1157),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1491),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1393),
.Y(n_1519)
);

OR2x2_ASAP7_75t_SL g1520 ( 
.A(n_1415),
.B(n_1327),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1456),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1375),
.B(n_1313),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1378),
.B(n_1162),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1433),
.Y(n_1524)
);

BUFx4f_ASAP7_75t_L g1525 ( 
.A(n_1356),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1389),
.Y(n_1526)
);

NAND2xp33_ASAP7_75t_SL g1527 ( 
.A(n_1447),
.B(n_1269),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1375),
.B(n_1315),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1376),
.B(n_1342),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1441),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1356),
.B(n_1363),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1385),
.B(n_1170),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1453),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1376),
.B(n_1342),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1457),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1356),
.B(n_1221),
.Y(n_1536)
);

AND2x6_ASAP7_75t_SL g1537 ( 
.A(n_1359),
.B(n_1217),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1459),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1462),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1442),
.A2(n_1318),
.B(n_1331),
.C(n_1322),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1355),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1380),
.B(n_1273),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1463),
.B(n_1323),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1386),
.B(n_1333),
.Y(n_1545)
);

INVx5_ASAP7_75t_L g1546 ( 
.A(n_1367),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1479),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1482),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1381),
.B(n_1165),
.Y(n_1549)
);

BUFx12f_ASAP7_75t_L g1550 ( 
.A(n_1389),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1413),
.B(n_1253),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1358),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1408),
.B(n_1305),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1402),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1411),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1442),
.A2(n_1165),
.B1(n_1346),
.B2(n_1343),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1408),
.B(n_1343),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1413),
.B(n_1219),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1393),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1404),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1387),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1377),
.B(n_1223),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1444),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1395),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1463),
.A2(n_1242),
.B1(n_1209),
.B2(n_1320),
.Y(n_1565)
);

BUFx4f_ASAP7_75t_SL g1566 ( 
.A(n_1392),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1414),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1354),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1367),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1444),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1383),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1423),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1472),
.B(n_1454),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1455),
.B(n_1480),
.Y(n_1574)
);

NAND2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1444),
.B(n_1328),
.Y(n_1575)
);

NOR2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1369),
.B(n_1221),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1418),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1455),
.B(n_1225),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1362),
.B(n_1262),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1353),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1360),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1364),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1361),
.B(n_1500),
.Y(n_1583)
);

BUFx12f_ASAP7_75t_SL g1584 ( 
.A(n_1485),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1403),
.A2(n_1321),
.B1(n_1172),
.B2(n_1207),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1373),
.B(n_1394),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1366),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1372),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1383),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1397),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1367),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1368),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1573),
.B(n_1403),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1574),
.B(n_1451),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1549),
.B(n_1431),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1515),
.B(n_1568),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1544),
.B(n_1451),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1507),
.B(n_1576),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1544),
.B(n_1243),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1541),
.B(n_1559),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1553),
.B(n_1464),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1553),
.B(n_1486),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1578),
.B(n_1421),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1507),
.B(n_1486),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_SL g1605 ( 
.A(n_1551),
.B(n_1494),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1512),
.B(n_1432),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1525),
.B(n_1432),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1510),
.B(n_1405),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1525),
.B(n_1439),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1519),
.B(n_1439),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1592),
.B(n_1405),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1510),
.B(n_1498),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1505),
.B(n_1419),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1583),
.B(n_1477),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1506),
.B(n_1484),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1522),
.B(n_1502),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1542),
.B(n_1204),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1542),
.B(n_1233),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1542),
.B(n_1233),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1549),
.B(n_1510),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1549),
.B(n_1233),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1562),
.B(n_1480),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1528),
.B(n_1409),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1565),
.B(n_1427),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1566),
.B(n_1449),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1558),
.B(n_1591),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1440),
.Y(n_1627)
);

NAND2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1591),
.B(n_1494),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1545),
.B(n_1474),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1586),
.B(n_1445),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1556),
.B(n_1407),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1585),
.B(n_1466),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1446),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1581),
.B(n_1428),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1581),
.B(n_1357),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1582),
.B(n_1434),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1571),
.B(n_1503),
.Y(n_1637)
);

NAND2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1569),
.B(n_1502),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1582),
.B(n_1460),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1546),
.B(n_1412),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1554),
.B(n_1370),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1546),
.B(n_1417),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1555),
.B(n_1371),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1546),
.B(n_1262),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_SL g1645 ( 
.A(n_1571),
.B(n_1503),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1615),
.B(n_1533),
.Y(n_1646)
);

NAND2x1_ASAP7_75t_L g1647 ( 
.A(n_1630),
.B(n_1569),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1594),
.B(n_1533),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1626),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1626),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1632),
.A2(n_1540),
.B(n_1534),
.Y(n_1651)
);

AO21x1_ASAP7_75t_L g1652 ( 
.A1(n_1616),
.A2(n_1532),
.B(n_1579),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1622),
.B(n_1529),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

BUFx4f_ASAP7_75t_L g1655 ( 
.A(n_1612),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1643),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1639),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1599),
.A2(n_1531),
.B1(n_1390),
.B2(n_1424),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_L g1659 ( 
.A(n_1608),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1640),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1606),
.A2(n_1584),
.B1(n_1490),
.B2(n_1531),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1642),
.B(n_1546),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1613),
.B(n_1529),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1641),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1595),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1635),
.A2(n_1437),
.B(n_1579),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1603),
.B(n_1534),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1602),
.A2(n_1540),
.B(n_1406),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1597),
.B(n_1546),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1633),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1598),
.Y(n_1671)
);

AND3x1_ASAP7_75t_SL g1672 ( 
.A(n_1604),
.B(n_1167),
.C(n_568),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1637),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1634),
.A2(n_1496),
.B1(n_1406),
.B2(n_1536),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1593),
.B(n_1511),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1601),
.B(n_1538),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1538),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1631),
.B(n_1539),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1605),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1624),
.B(n_1514),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1595),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1605),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1616),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1629),
.B(n_1518),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1628),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1645),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1614),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1620),
.B(n_1539),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1595),
.B(n_1548),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1596),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1611),
.A2(n_1531),
.B1(n_1166),
.B2(n_1523),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1600),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1628),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1651),
.A2(n_1429),
.B(n_1557),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1666),
.A2(n_1591),
.B(n_1569),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1647),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1666),
.A2(n_1388),
.B(n_1443),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1670),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1666),
.A2(n_1458),
.B(n_1452),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1692),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1670),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1649),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1609),
.Y(n_1706)
);

AO21x2_ASAP7_75t_L g1707 ( 
.A1(n_1651),
.A2(n_1668),
.B(n_1652),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1649),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1607),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_SL g1710 ( 
.A1(n_1652),
.A2(n_1420),
.B(n_1401),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1650),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1647),
.A2(n_1272),
.B(n_1400),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1659),
.B(n_1610),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1654),
.B(n_1617),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1654),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1650),
.A2(n_1422),
.B(n_1495),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1660),
.B(n_1508),
.Y(n_1717)
);

CKINVDCx16_ASAP7_75t_R g1718 ( 
.A(n_1671),
.Y(n_1718)
);

AOI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1657),
.A2(n_1619),
.B(n_1618),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1646),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1646),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1654),
.Y(n_1722)
);

INVx8_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1684),
.A2(n_1469),
.B(n_1461),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1664),
.B(n_1567),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1692),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1678),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1654),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_L g1729 ( 
.A(n_1673),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1684),
.A2(n_1426),
.B(n_1379),
.Y(n_1731)
);

BUFx10_ASAP7_75t_L g1732 ( 
.A(n_1656),
.Y(n_1732)
);

INVx5_ASAP7_75t_L g1733 ( 
.A(n_1654),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1654),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1678),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1680),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1683),
.Y(n_1737)
);

BUFx12f_ASAP7_75t_L g1738 ( 
.A(n_1687),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1692),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1694),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1683),
.A2(n_1426),
.B(n_1379),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1668),
.A2(n_1532),
.B(n_1391),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1678),
.Y(n_1743)
);

NAND2x1_ASAP7_75t_L g1744 ( 
.A(n_1686),
.B(n_1367),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1679),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1686),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1679),
.Y(n_1747)
);

AO21x2_ASAP7_75t_L g1748 ( 
.A1(n_1695),
.A2(n_1425),
.B(n_1488),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1660),
.B(n_1621),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1648),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1695),
.A2(n_1669),
.B(n_1667),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1664),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1677),
.B(n_1166),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1648),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1662),
.A2(n_1473),
.B(n_1471),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1660),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1667),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1662),
.A2(n_1499),
.B(n_1475),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1656),
.B(n_1577),
.Y(n_1759)
);

INVx5_ASAP7_75t_L g1760 ( 
.A(n_1676),
.Y(n_1760)
);

BUFx2_ASAP7_75t_SL g1761 ( 
.A(n_1694),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1659),
.B(n_1509),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1662),
.A2(n_1501),
.B(n_1448),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1689),
.B(n_1584),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1688),
.A2(n_826),
.B(n_822),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1665),
.Y(n_1766)
);

OAI21x1_ASAP7_75t_L g1767 ( 
.A1(n_1663),
.A2(n_1436),
.B(n_1274),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1694),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1663),
.A2(n_1283),
.B(n_1261),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1682),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1676),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1688),
.A2(n_1276),
.B(n_1430),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1665),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1653),
.A2(n_1276),
.B(n_1575),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1682),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1682),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1653),
.A2(n_1425),
.B(n_1438),
.Y(n_1777)
);

CKINVDCx16_ASAP7_75t_R g1778 ( 
.A(n_1693),
.Y(n_1778)
);

BUFx2_ASAP7_75t_R g1779 ( 
.A(n_1675),
.Y(n_1779)
);

AO21x2_ASAP7_75t_L g1780 ( 
.A1(n_1658),
.A2(n_1396),
.B(n_1398),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1677),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1730),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1727),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1730),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1778),
.A2(n_1674),
.B1(n_1166),
.B2(n_534),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1727),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1740),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1718),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1729),
.Y(n_1789)
);

BUFx12f_ASAP7_75t_L g1790 ( 
.A(n_1729),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1718),
.A2(n_1520),
.B1(n_1521),
.B2(n_1334),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1723),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1727),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1736),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1735),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1778),
.A2(n_1674),
.B1(n_534),
.B2(n_520),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1707),
.A2(n_1742),
.B1(n_1659),
.B2(n_1761),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1703),
.Y(n_1798)
);

CKINVDCx6p67_ASAP7_75t_R g1799 ( 
.A(n_1729),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1757),
.B(n_1685),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1707),
.A2(n_1659),
.B1(n_1655),
.B2(n_1685),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1753),
.A2(n_523),
.B1(n_537),
.B2(n_506),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1740),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1761),
.A2(n_1521),
.B1(n_1589),
.B2(n_1526),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1736),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1737),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1738),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1738),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1709),
.A2(n_1658),
.B(n_1435),
.Y(n_1809)
);

BUFx12f_ASAP7_75t_L g1810 ( 
.A(n_1738),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1737),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1779),
.A2(n_1693),
.B1(n_1661),
.B2(n_1655),
.Y(n_1812)
);

CKINVDCx11_ASAP7_75t_R g1813 ( 
.A(n_1723),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1768),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1735),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1735),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1723),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1705),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1753),
.A2(n_537),
.B1(n_539),
.B2(n_523),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1771),
.B(n_1655),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1705),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1708),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1728),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1708),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1754),
.B(n_1768),
.Y(n_1825)
);

CKINVDCx12_ASAP7_75t_R g1826 ( 
.A(n_1717),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1707),
.A2(n_561),
.B1(n_568),
.B2(n_539),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1713),
.A2(n_1655),
.B1(n_1536),
.B2(n_1531),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1711),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1711),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1743),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1743),
.Y(n_1832)
);

BUFx12f_ASAP7_75t_L g1833 ( 
.A(n_1766),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1707),
.A2(n_561),
.B1(n_576),
.B2(n_569),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1780),
.A2(n_1681),
.B1(n_1675),
.B2(n_1280),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1723),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1780),
.A2(n_1681),
.B1(n_1280),
.B2(n_1536),
.Y(n_1837)
);

BUFx10_ASAP7_75t_L g1838 ( 
.A(n_1764),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1709),
.A2(n_1625),
.B(n_1496),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1754),
.Y(n_1840)
);

BUFx10_ASAP7_75t_L g1841 ( 
.A(n_1728),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1703),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1752),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1754),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1780),
.A2(n_569),
.B1(n_579),
.B2(n_576),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1728),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1703),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1757),
.B(n_1690),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1752),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1700),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1706),
.B(n_1690),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1706),
.A2(n_1536),
.B1(n_1334),
.B2(n_1589),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1752),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1726),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1780),
.A2(n_579),
.B1(n_590),
.B2(n_586),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1726),
.A2(n_1334),
.B1(n_1526),
.B2(n_1497),
.Y(n_1856)
);

CKINVDCx6p67_ASAP7_75t_R g1857 ( 
.A(n_1723),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1696),
.A2(n_586),
.B1(n_595),
.B2(n_590),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1714),
.A2(n_1672),
.B1(n_1527),
.B2(n_1450),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1726),
.A2(n_1497),
.B1(n_1587),
.B2(n_1580),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1696),
.A2(n_595),
.B1(n_607),
.B2(n_598),
.Y(n_1861)
);

BUFx8_ASAP7_75t_L g1862 ( 
.A(n_1728),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1739),
.B(n_1691),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1747),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1696),
.A2(n_598),
.B1(n_610),
.B2(n_607),
.Y(n_1865)
);

INVx6_ASAP7_75t_L g1866 ( 
.A(n_1733),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1696),
.A2(n_610),
.B1(n_625),
.B2(n_622),
.Y(n_1867)
);

CKINVDCx11_ASAP7_75t_R g1868 ( 
.A(n_1728),
.Y(n_1868)
);

INVxp67_ASAP7_75t_SL g1869 ( 
.A(n_1756),
.Y(n_1869)
);

BUFx12f_ASAP7_75t_L g1870 ( 
.A(n_1766),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1700),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1739),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1759),
.A2(n_625),
.B1(n_633),
.B2(n_622),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1714),
.A2(n_1280),
.B1(n_543),
.B2(n_1691),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1747),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1714),
.A2(n_543),
.B1(n_1550),
.B2(n_1508),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1701),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1701),
.Y(n_1878)
);

CKINVDCx11_ASAP7_75t_R g1879 ( 
.A(n_1728),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1781),
.B(n_1537),
.Y(n_1880)
);

INVx6_ASAP7_75t_L g1881 ( 
.A(n_1733),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_1739),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1747),
.Y(n_1883)
);

INVx6_ASAP7_75t_L g1884 ( 
.A(n_1733),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1721),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1704),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1733),
.A2(n_643),
.B1(n_647),
.B2(n_633),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1704),
.Y(n_1888)
);

INVx11_ASAP7_75t_L g1889 ( 
.A(n_1770),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1714),
.A2(n_1478),
.B(n_647),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1721),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1750),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1770),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1750),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1749),
.A2(n_1588),
.B1(n_1550),
.B2(n_1523),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1765),
.A2(n_1638),
.B(n_1508),
.Y(n_1896)
);

INVx5_ASAP7_75t_L g1897 ( 
.A(n_1732),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1721),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1777),
.A2(n_653),
.B1(n_667),
.B2(n_643),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1715),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1746),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1746),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1746),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1770),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1746),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1777),
.A2(n_667),
.B1(n_671),
.B2(n_653),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1751),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1749),
.A2(n_1523),
.B1(n_1517),
.B2(n_1481),
.Y(n_1908)
);

BUFx12f_ASAP7_75t_L g1909 ( 
.A(n_1766),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1781),
.B(n_1524),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1756),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1756),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1776),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1749),
.A2(n_1517),
.B1(n_1470),
.B2(n_1410),
.Y(n_1914)
);

BUFx12f_ASAP7_75t_L g1915 ( 
.A(n_1766),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1745),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1720),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1722),
.B(n_671),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1720),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1722),
.B(n_679),
.Y(n_1920)
);

INVx8_ASAP7_75t_L g1921 ( 
.A(n_1717),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1922)
);

BUFx12f_ASAP7_75t_L g1923 ( 
.A(n_1773),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1733),
.A2(n_1508),
.B1(n_682),
.B2(n_683),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_1776),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1777),
.A2(n_682),
.B1(n_683),
.B2(n_679),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1733),
.A2(n_1773),
.B1(n_1760),
.B2(n_1715),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1777),
.A2(n_689),
.B1(n_697),
.B2(n_687),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1751),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_SL g1930 ( 
.A1(n_1773),
.A2(n_689),
.B1(n_697),
.B2(n_687),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1776),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1751),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1751),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1889),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1796),
.A2(n_1710),
.B(n_1638),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1917),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1796),
.A2(n_713),
.B1(n_716),
.B2(n_705),
.C(n_702),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1825),
.B(n_1760),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1782),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1809),
.B(n_1773),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1790),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1838),
.B(n_1880),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1873),
.A2(n_713),
.B1(n_716),
.B2(n_705),
.C(n_702),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1784),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1845),
.A2(n_1772),
.B(n_1724),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1933),
.A2(n_1932),
.B(n_1929),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1794),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1921),
.B(n_1717),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1851),
.B(n_1722),
.Y(n_1950)
);

OA21x2_ASAP7_75t_L g1951 ( 
.A1(n_1929),
.A2(n_1724),
.B(n_1772),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1917),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1953)
);

AOI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1852),
.A2(n_1719),
.B(n_1744),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1805),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1813),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1785),
.A2(n_725),
.B(n_724),
.Y(n_1957)
);

AO31x2_ASAP7_75t_L g1958 ( 
.A1(n_1896),
.A2(n_1715),
.A3(n_1765),
.B(n_725),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1845),
.A2(n_1710),
.B(n_1765),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1806),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1932),
.A2(n_1774),
.B(n_1699),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1907),
.A2(n_1855),
.B(n_1899),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1907),
.A2(n_1774),
.B(n_1697),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1811),
.Y(n_1964)
);

O2A1O1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1839),
.A2(n_724),
.B(n_1734),
.C(n_829),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1818),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1855),
.A2(n_1719),
.B(n_1765),
.Y(n_1967)
);

NAND2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1897),
.B(n_1760),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1785),
.A2(n_1699),
.B(n_1712),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1790),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1838),
.B(n_1715),
.Y(n_1971)
);

AO21x2_ASAP7_75t_L g1972 ( 
.A1(n_1887),
.A2(n_1697),
.B(n_1702),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1854),
.B(n_1760),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1821),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1788),
.B(n_1722),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1913),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1899),
.A2(n_1717),
.B(n_1744),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1810),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1824),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1827),
.A2(n_1834),
.B1(n_1819),
.B2(n_1802),
.Y(n_1980)
);

A2O1A1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1890),
.A2(n_1527),
.B(n_1734),
.C(n_830),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1827),
.A2(n_1834),
.B1(n_1819),
.B2(n_1802),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1919),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1804),
.A2(n_835),
.B(n_839),
.C(n_827),
.Y(n_1984)
);

AO22x2_ASAP7_75t_L g1985 ( 
.A1(n_1829),
.A2(n_1698),
.B1(n_1775),
.B2(n_1732),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1919),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1791),
.B(n_1808),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1842),
.B(n_1698),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1789),
.B(n_1799),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1848),
.B(n_1892),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1864),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1810),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1807),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1904),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1906),
.A2(n_1717),
.B(n_1762),
.Y(n_1995)
);

OA21x2_ASAP7_75t_L g1996 ( 
.A1(n_1906),
.A2(n_1702),
.B(n_1731),
.Y(n_1996)
);

OA21x2_ASAP7_75t_L g1997 ( 
.A1(n_1926),
.A2(n_1741),
.B(n_1731),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1840),
.B(n_1698),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1873),
.A2(n_531),
.B1(n_536),
.B2(n_528),
.C(n_526),
.Y(n_1999)
);

OA21x2_ASAP7_75t_L g2000 ( 
.A1(n_1926),
.A2(n_1741),
.B(n_1769),
.Y(n_2000)
);

NAND2x1_ASAP7_75t_L g2001 ( 
.A(n_1866),
.B(n_1698),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1864),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1830),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_SL g2004 ( 
.A1(n_1895),
.A2(n_1775),
.B(n_1732),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1812),
.A2(n_721),
.B1(n_1748),
.B2(n_1346),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1928),
.A2(n_1762),
.B(n_1748),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1882),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_SL g2008 ( 
.A1(n_1800),
.A2(n_1732),
.B(n_1572),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1874),
.A2(n_1762),
.B1(n_585),
.B2(n_596),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1859),
.A2(n_841),
.B(n_840),
.C(n_599),
.Y(n_2010)
);

A2O1A1Ixp33_ASAP7_75t_L g2011 ( 
.A1(n_1876),
.A2(n_544),
.B(n_545),
.C(n_542),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1894),
.B(n_1748),
.Y(n_2012)
);

OA21x2_ASAP7_75t_L g2013 ( 
.A1(n_1928),
.A2(n_1769),
.B(n_1712),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1822),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1900),
.A2(n_1767),
.B(n_1716),
.Y(n_2015)
);

NAND3xp33_ASAP7_75t_L g2016 ( 
.A(n_1858),
.B(n_721),
.C(n_549),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1858),
.A2(n_1767),
.B(n_1716),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1828),
.A2(n_1748),
.B1(n_1346),
.B2(n_1517),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1861),
.A2(n_1763),
.B(n_1758),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1861),
.A2(n_1763),
.B(n_1758),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1930),
.A2(n_1837),
.B1(n_1856),
.B2(n_1887),
.Y(n_2021)
);

A2O1A1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1797),
.A2(n_550),
.B(n_551),
.C(n_548),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1865),
.A2(n_1755),
.B(n_1416),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1865),
.A2(n_1755),
.B(n_1202),
.Y(n_2024)
);

OAI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_1835),
.A2(n_558),
.B1(n_559),
.B2(n_554),
.C(n_553),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1822),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1867),
.A2(n_564),
.B(n_566),
.C(n_563),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_SL g2028 ( 
.A1(n_1921),
.A2(n_721),
.B1(n_588),
.B2(n_589),
.Y(n_2028)
);

AO21x2_ASAP7_75t_L g2029 ( 
.A1(n_1831),
.A2(n_1345),
.B(n_860),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1867),
.A2(n_1468),
.B(n_1465),
.Y(n_2030)
);

AO31x2_ASAP7_75t_L g2031 ( 
.A1(n_1901),
.A2(n_1489),
.A3(n_1492),
.B(n_1487),
.Y(n_2031)
);

OAI21x1_ASAP7_75t_L g2032 ( 
.A1(n_1900),
.A2(n_1575),
.B(n_1572),
.Y(n_2032)
);

NOR2xp67_ASAP7_75t_L g2033 ( 
.A(n_1911),
.B(n_3),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1914),
.A2(n_1468),
.B(n_1465),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1787),
.B(n_857),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1916),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1801),
.A2(n_593),
.B1(n_594),
.B2(n_578),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1875),
.Y(n_2038)
);

AO31x2_ASAP7_75t_L g2039 ( 
.A1(n_1901),
.A2(n_1489),
.A3(n_1492),
.B(n_1487),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1875),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1832),
.Y(n_2041)
);

OAI21x1_ASAP7_75t_L g2042 ( 
.A1(n_1910),
.A2(n_1227),
.B(n_1226),
.Y(n_2042)
);

AO21x1_ASAP7_75t_L g2043 ( 
.A1(n_1918),
.A2(n_860),
.B(n_857),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1850),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1871),
.Y(n_2045)
);

OA21x2_ASAP7_75t_L g2046 ( 
.A1(n_1902),
.A2(n_862),
.B(n_861),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1877),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1820),
.B(n_861),
.Y(n_2048)
);

BUFx12f_ASAP7_75t_L g2049 ( 
.A(n_1833),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1803),
.B(n_862),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1925),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1913),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1897),
.B(n_1509),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1814),
.B(n_1863),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1897),
.A2(n_1493),
.B(n_1299),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1842),
.B(n_1863),
.Y(n_2056)
);

OA21x2_ASAP7_75t_L g2057 ( 
.A1(n_1902),
.A2(n_866),
.B(n_863),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1897),
.A2(n_1493),
.B(n_1299),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1878),
.Y(n_2059)
);

OR2x6_ASAP7_75t_L g2060 ( 
.A(n_1921),
.B(n_1509),
.Y(n_2060)
);

OAI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1924),
.A2(n_1319),
.B(n_1316),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1920),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1886),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1908),
.A2(n_1287),
.B(n_1291),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1888),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1860),
.A2(n_1287),
.B(n_1291),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1883),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1913),
.Y(n_2068)
);

CKINVDCx11_ASAP7_75t_R g2069 ( 
.A(n_1909),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1911),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1844),
.B(n_1922),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_1883),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1912),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_SL g2074 ( 
.A1(n_1927),
.A2(n_1319),
.B1(n_1316),
.B2(n_1309),
.C(n_866),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1923),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_1913),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1847),
.B(n_863),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_1870),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_SL g2079 ( 
.A1(n_1870),
.A2(n_605),
.B1(n_613),
.B2(n_604),
.Y(n_2079)
);

OA21x2_ASAP7_75t_L g2080 ( 
.A1(n_1903),
.A2(n_616),
.B(n_615),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1866),
.A2(n_627),
.B1(n_634),
.B2(n_620),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1869),
.B(n_636),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1862),
.Y(n_2083)
);

OAI21x1_ASAP7_75t_L g2084 ( 
.A1(n_1783),
.A2(n_1238),
.B(n_1230),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1866),
.A2(n_640),
.B1(n_642),
.B2(n_638),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1885),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1881),
.A2(n_648),
.B1(n_649),
.B2(n_645),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1912),
.Y(n_2088)
);

OA21x2_ASAP7_75t_L g2089 ( 
.A1(n_1903),
.A2(n_652),
.B(n_650),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1872),
.A2(n_657),
.B(n_658),
.C(n_656),
.Y(n_2090)
);

AOI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_1957),
.A2(n_668),
.B1(n_672),
.B2(n_666),
.C(n_665),
.Y(n_2091)
);

BUFx12f_ASAP7_75t_L g2092 ( 
.A(n_1978),
.Y(n_2092)
);

A2O1A1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_1957),
.A2(n_2010),
.B(n_1965),
.C(n_2021),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1980),
.A2(n_1915),
.B1(n_1792),
.B2(n_1836),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2056),
.B(n_1885),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_1950),
.B(n_1891),
.Y(n_2096)
);

OAI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_2028),
.A2(n_686),
.B1(n_693),
.B2(n_685),
.C(n_673),
.Y(n_2097)
);

AOI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2037),
.A2(n_709),
.B1(n_710),
.B2(n_700),
.C(n_695),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_1954),
.A2(n_1786),
.B(n_1783),
.Y(n_2099)
);

OAI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2021),
.A2(n_1881),
.B1(n_1884),
.B2(n_1857),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_1980),
.A2(n_1792),
.B1(n_1836),
.B2(n_1817),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1938),
.B(n_1891),
.Y(n_2102)
);

OAI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1982),
.A2(n_1817),
.B1(n_1915),
.B2(n_1884),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1991),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1940),
.A2(n_1982),
.B(n_2016),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1990),
.B(n_1898),
.Y(n_2106)
);

OAI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2037),
.A2(n_1884),
.B1(n_1881),
.B2(n_1893),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1990),
.B(n_1898),
.Y(n_2108)
);

AOI21xp33_ASAP7_75t_L g2109 ( 
.A1(n_2081),
.A2(n_1931),
.B(n_1846),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1939),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1944),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2016),
.A2(n_1905),
.B(n_1793),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2009),
.A2(n_1879),
.B1(n_1868),
.B2(n_1823),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_1992),
.Y(n_2114)
);

OAI221xp5_ASAP7_75t_L g2115 ( 
.A1(n_2079),
.A2(n_719),
.B1(n_722),
.B2(n_717),
.C(n_712),
.Y(n_2115)
);

AOI222xp33_ASAP7_75t_L g2116 ( 
.A1(n_1937),
.A2(n_488),
.B1(n_479),
.B2(n_489),
.C1(n_487),
.C2(n_477),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1948),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1955),
.Y(n_2118)
);

HB1xp67_ASAP7_75t_L g2119 ( 
.A(n_2072),
.Y(n_2119)
);

BUFx4f_ASAP7_75t_SL g2120 ( 
.A(n_2049),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2054),
.B(n_1905),
.Y(n_2121)
);

OAI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2022),
.A2(n_1846),
.B1(n_1823),
.B2(n_1795),
.C(n_1815),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_2005),
.A2(n_1846),
.B1(n_1823),
.B2(n_1843),
.Y(n_2123)
);

NOR2x1p5_ASAP7_75t_L g2124 ( 
.A(n_1956),
.B(n_1823),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2009),
.A2(n_1846),
.B1(n_1795),
.B2(n_1815),
.C(n_1793),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2068),
.B(n_1973),
.Y(n_2126)
);

AOI221xp5_ASAP7_75t_L g2127 ( 
.A1(n_1943),
.A2(n_505),
.B1(n_507),
.B2(n_504),
.C(n_491),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_1998),
.B(n_1786),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2025),
.A2(n_516),
.B1(n_521),
.B2(n_514),
.C(n_508),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2071),
.B(n_1816),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_1942),
.A2(n_1862),
.B1(n_1308),
.B2(n_849),
.Y(n_2131)
);

AOI21xp33_ASAP7_75t_SL g2132 ( 
.A1(n_1989),
.A2(n_3),
.B(n_4),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_2015),
.A2(n_1961),
.B(n_1968),
.Y(n_2133)
);

NAND4xp25_ASAP7_75t_SL g2134 ( 
.A(n_2011),
.B(n_1826),
.C(n_6),
.D(n_4),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_SL g2135 ( 
.A1(n_2080),
.A2(n_1841),
.B1(n_1816),
.B2(n_1843),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2076),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1947),
.B(n_1849),
.Y(n_2137)
);

OAI211xp5_ASAP7_75t_SL g2138 ( 
.A1(n_1999),
.A2(n_1853),
.B(n_1849),
.C(n_751),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1947),
.B(n_1853),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1981),
.A2(n_1535),
.B1(n_1543),
.B2(n_1530),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1953),
.B(n_2007),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2002),
.Y(n_2142)
);

NAND2x1p5_ASAP7_75t_L g2143 ( 
.A(n_2001),
.B(n_1841),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1988),
.B(n_1509),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2071),
.B(n_1936),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_1975),
.A2(n_1308),
.B1(n_1241),
.B2(n_677),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2048),
.B(n_5),
.Y(n_2147)
);

INVx4_ASAP7_75t_L g2148 ( 
.A(n_1956),
.Y(n_2148)
);

INVx4_ASAP7_75t_L g2149 ( 
.A(n_1956),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2038),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_SL g2151 ( 
.A1(n_2080),
.A2(n_529),
.B1(n_535),
.B2(n_527),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2033),
.A2(n_1547),
.B1(n_1561),
.B2(n_1552),
.Y(n_2152)
);

OAI221xp5_ASAP7_75t_L g2153 ( 
.A1(n_2027),
.A2(n_560),
.B1(n_571),
.B2(n_557),
.C(n_538),
.Y(n_2153)
);

AOI22xp33_ASAP7_75t_SL g2154 ( 
.A1(n_2089),
.A2(n_574),
.B1(n_587),
.B2(n_572),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1935),
.A2(n_1561),
.B1(n_1564),
.B2(n_1552),
.Y(n_2155)
);

A2O1A1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_2033),
.A2(n_592),
.B(n_597),
.C(n_591),
.Y(n_2156)
);

OA21x2_ASAP7_75t_L g2157 ( 
.A1(n_2012),
.A2(n_751),
.B(n_749),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1953),
.B(n_5),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1960),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1987),
.A2(n_1308),
.B1(n_1163),
.B2(n_1159),
.Y(n_2160)
);

AOI21xp33_ASAP7_75t_L g2161 ( 
.A1(n_2081),
.A2(n_6),
.B(n_7),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2018),
.A2(n_1564),
.B1(n_1548),
.B2(n_1560),
.Y(n_2162)
);

OAI211xp5_ASAP7_75t_L g2163 ( 
.A1(n_1969),
.A2(n_609),
.B(n_614),
.C(n_603),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2018),
.A2(n_1560),
.B1(n_1563),
.B2(n_1513),
.Y(n_2164)
);

AOI222xp33_ASAP7_75t_L g2165 ( 
.A1(n_2061),
.A2(n_631),
.B1(n_621),
.B2(n_635),
.C1(n_628),
.C2(n_619),
.Y(n_2165)
);

OAI21xp33_ASAP7_75t_L g2166 ( 
.A1(n_1969),
.A2(n_644),
.B(n_637),
.Y(n_2166)
);

AOI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_2089),
.A2(n_1308),
.B1(n_1163),
.B2(n_1159),
.Y(n_2167)
);

AOI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_2062),
.A2(n_1308),
.B1(n_1186),
.B2(n_1192),
.Y(n_2168)
);

INVx4_ASAP7_75t_L g2169 ( 
.A(n_1992),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1988),
.B(n_1513),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_1992),
.A2(n_1186),
.B1(n_1192),
.B2(n_1182),
.Y(n_2171)
);

OAI221xp5_ASAP7_75t_SL g2172 ( 
.A1(n_1959),
.A2(n_1309),
.B1(n_9),
.B2(n_7),
.C(n_8),
.Y(n_2172)
);

OAI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_1995),
.A2(n_1560),
.B1(n_1563),
.B2(n_1513),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2078),
.A2(n_1962),
.B1(n_2087),
.B2(n_2085),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1976),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2006),
.A2(n_669),
.B(n_688),
.C(n_661),
.Y(n_2176)
);

A2O1A1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2090),
.A2(n_704),
.B(n_706),
.C(n_694),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1964),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1976),
.B(n_8),
.Y(n_2179)
);

OAI21x1_ASAP7_75t_L g2180 ( 
.A1(n_1968),
.A2(n_1516),
.B(n_1345),
.Y(n_2180)
);

AOI221xp5_ASAP7_75t_L g2181 ( 
.A1(n_2082),
.A2(n_715),
.B1(n_714),
.B2(n_753),
.C(n_749),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_SL g2182 ( 
.A1(n_1962),
.A2(n_1560),
.B1(n_1563),
.B2(n_1513),
.Y(n_2182)
);

OAI211xp5_ASAP7_75t_L g2183 ( 
.A1(n_1967),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_2183)
);

AOI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2085),
.A2(n_758),
.B1(n_756),
.B2(n_753),
.C(n_12),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_SL g2185 ( 
.A1(n_1994),
.A2(n_1570),
.B1(n_1563),
.B2(n_14),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1966),
.B(n_10),
.Y(n_2186)
);

OAI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2087),
.A2(n_758),
.B1(n_756),
.B2(n_1516),
.C(n_15),
.Y(n_2187)
);

OAI221xp5_ASAP7_75t_L g2188 ( 
.A1(n_1971),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.C(n_16),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2024),
.A2(n_1325),
.B(n_1302),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1974),
.B(n_17),
.Y(n_2190)
);

OAI211xp5_ASAP7_75t_L g2191 ( 
.A1(n_1967),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1979),
.B(n_19),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2061),
.A2(n_1186),
.B1(n_1192),
.B2(n_1182),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2077),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.C(n_23),
.Y(n_2194)
);

AOI221xp5_ASAP7_75t_L g2195 ( 
.A1(n_2035),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.C(n_29),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_1952),
.B(n_24),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2040),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2003),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_1941),
.A2(n_1186),
.B1(n_1192),
.B2(n_1182),
.Y(n_2199)
);

AOI221xp5_ASAP7_75t_L g2200 ( 
.A1(n_2050),
.A2(n_35),
.B1(n_30),
.B2(n_31),
.C(n_37),
.Y(n_2200)
);

CKINVDCx11_ASAP7_75t_R g2201 ( 
.A(n_2069),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2017),
.A2(n_1186),
.B(n_1182),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1970),
.A2(n_1265),
.B1(n_1192),
.B2(n_1570),
.Y(n_2203)
);

NAND4xp25_ASAP7_75t_L g2204 ( 
.A(n_1984),
.B(n_42),
.C(n_39),
.D(n_40),
.Y(n_2204)
);

OAI221xp5_ASAP7_75t_L g2205 ( 
.A1(n_1993),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.C(n_44),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2083),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2014),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_1949),
.A2(n_1265),
.B1(n_1570),
.B2(n_1262),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2074),
.A2(n_1570),
.B1(n_47),
.B2(n_43),
.Y(n_2209)
);

AOI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_1949),
.A2(n_1265),
.B1(n_1296),
.B2(n_1444),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_1949),
.A2(n_1265),
.B1(n_1502),
.B2(n_1494),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2075),
.Y(n_2212)
);

INVxp33_ASAP7_75t_L g2213 ( 
.A(n_2051),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2067),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_2070),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_SL g2216 ( 
.A1(n_2004),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_2216)
);

AOI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2017),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.C(n_53),
.Y(n_2217)
);

AOI21xp33_ASAP7_75t_L g2218 ( 
.A1(n_2008),
.A2(n_49),
.B(n_50),
.Y(n_2218)
);

OAI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_1977),
.A2(n_1504),
.B1(n_1214),
.B2(n_1229),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2026),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_SL g2221 ( 
.A1(n_1945),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2052),
.B(n_55),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2043),
.A2(n_1265),
.B1(n_1267),
.B2(n_1247),
.Y(n_2223)
);

OAI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_2060),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.Y(n_2224)
);

AOI222xp33_ASAP7_75t_L g2225 ( 
.A1(n_1945),
.A2(n_2045),
.B1(n_2041),
.B2(n_2059),
.C1(n_2047),
.C2(n_2044),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2063),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_SL g2227 ( 
.A1(n_1985),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_2073),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2065),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1934),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_1983),
.B(n_61),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2034),
.A2(n_1267),
.B1(n_1310),
.B2(n_1247),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_2086),
.Y(n_2233)
);

INVx5_ASAP7_75t_L g2234 ( 
.A(n_2060),
.Y(n_2234)
);

OAI221xp5_ASAP7_75t_SL g2235 ( 
.A1(n_2019),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.C(n_71),
.Y(n_2235)
);

OAI22xp33_ASAP7_75t_SL g2236 ( 
.A1(n_2012),
.A2(n_73),
.B1(n_65),
.B2(n_72),
.Y(n_2236)
);

BUFx3_ASAP7_75t_L g2237 ( 
.A(n_2060),
.Y(n_2237)
);

AOI22xp33_ASAP7_75t_L g2238 ( 
.A1(n_2023),
.A2(n_1494),
.B1(n_1502),
.B2(n_1310),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_1986),
.B(n_72),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2020),
.A2(n_1088),
.B1(n_1093),
.B2(n_1087),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_L g2241 ( 
.A1(n_2013),
.A2(n_1088),
.B1(n_1093),
.B2(n_1087),
.Y(n_2241)
);

AOI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2036),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.C(n_77),
.Y(n_2242)
);

OAI21x1_ASAP7_75t_SL g2243 ( 
.A1(n_2088),
.A2(n_77),
.B(n_78),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2030),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2244)
);

NAND3xp33_ASAP7_75t_L g2245 ( 
.A(n_2013),
.B(n_1229),
.C(n_1214),
.Y(n_2245)
);

OAI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_1997),
.A2(n_82),
.B(n_79),
.C(n_80),
.Y(n_2246)
);

OAI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_2053),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.Y(n_2247)
);

NOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2124),
.B(n_2046),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2121),
.B(n_1985),
.Y(n_2249)
);

OAI332xp33_ASAP7_75t_L g2250 ( 
.A1(n_2205),
.A2(n_83),
.A3(n_87),
.B1(n_90),
.B2(n_91),
.B3(n_92),
.C1(n_93),
.C2(n_94),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2215),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2207),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_2206),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_SL g2254 ( 
.A1(n_2105),
.A2(n_1997),
.B1(n_2000),
.B2(n_1996),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2126),
.B(n_1958),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2099),
.Y(n_2256)
);

NOR2x1_ASAP7_75t_SL g2257 ( 
.A(n_2234),
.B(n_1972),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2220),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2110),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2136),
.B(n_1958),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2141),
.B(n_1958),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2225),
.B(n_2000),
.Y(n_2262)
);

AO21x2_ASAP7_75t_L g2263 ( 
.A1(n_2133),
.A2(n_2032),
.B(n_1972),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2111),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2117),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2228),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2102),
.B(n_1963),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_2206),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2137),
.B(n_1963),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2119),
.B(n_2228),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2118),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2233),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2225),
.B(n_1996),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_2234),
.B(n_2144),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2139),
.B(n_1946),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2095),
.B(n_2175),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2175),
.B(n_1946),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2233),
.B(n_1951),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2145),
.B(n_2159),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2178),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2198),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2096),
.B(n_1951),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2226),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2229),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2130),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_2206),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2128),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2106),
.B(n_2031),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2104),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2108),
.B(n_2031),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2142),
.B(n_2031),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2150),
.B(n_2053),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2197),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2214),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_2201),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2196),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2231),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2143),
.B(n_2039),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2100),
.B(n_2039),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2239),
.Y(n_2300)
);

AND2x4_ASAP7_75t_SL g2301 ( 
.A(n_2148),
.B(n_2042),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2234),
.B(n_2084),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2186),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2190),
.Y(n_2304)
);

INVx2_ASAP7_75t_SL g2305 ( 
.A(n_2143),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2192),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_SL g2307 ( 
.A(n_2148),
.B(n_2055),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2179),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2157),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2234),
.B(n_2237),
.Y(n_2310)
);

OAI221xp5_ASAP7_75t_L g2311 ( 
.A1(n_2093),
.A2(n_2064),
.B1(n_2066),
.B2(n_2058),
.C(n_2057),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2112),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2144),
.B(n_2039),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_2092),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2170),
.B(n_2046),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2135),
.B(n_2174),
.Y(n_2316)
);

NOR2x1_ASAP7_75t_L g2317 ( 
.A(n_2149),
.B(n_2057),
.Y(n_2317)
);

AOI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2217),
.A2(n_2029),
.B1(n_95),
.B2(n_90),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2158),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2100),
.B(n_2029),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2114),
.Y(n_2321)
);

AOI21xp33_ASAP7_75t_L g2322 ( 
.A1(n_2165),
.A2(n_94),
.B(n_95),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2170),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2157),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2182),
.B(n_96),
.Y(n_2325)
);

INVxp67_ASAP7_75t_SL g2326 ( 
.A(n_2107),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2147),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2204),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_2328)
);

HB1xp67_ASAP7_75t_L g2329 ( 
.A(n_2173),
.Y(n_2329)
);

OR2x2_ASAP7_75t_L g2330 ( 
.A(n_2202),
.B(n_2125),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2222),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2169),
.B(n_98),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2180),
.B(n_99),
.Y(n_2333)
);

INVxp67_ASAP7_75t_L g2334 ( 
.A(n_2114),
.Y(n_2334)
);

OA21x2_ASAP7_75t_L g2335 ( 
.A1(n_2246),
.A2(n_1161),
.B(n_1249),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2202),
.B(n_100),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2169),
.B(n_101),
.Y(n_2337)
);

INVxp33_ASAP7_75t_SL g2338 ( 
.A(n_2212),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2103),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2114),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2094),
.B(n_101),
.Y(n_2341)
);

INVxp67_ASAP7_75t_L g2342 ( 
.A(n_2243),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2236),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2101),
.B(n_104),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2162),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2149),
.B(n_2230),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2213),
.B(n_105),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_2230),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2230),
.B(n_105),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2152),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2109),
.B(n_108),
.Y(n_2351)
);

INVx4_ASAP7_75t_L g2352 ( 
.A(n_2120),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2152),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2232),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2113),
.B(n_109),
.Y(n_2355)
);

NAND2x1_ASAP7_75t_L g2356 ( 
.A(n_2240),
.B(n_825),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2241),
.B(n_109),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_2204),
.A2(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2227),
.B(n_110),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2123),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2216),
.B(n_113),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2123),
.B(n_117),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2238),
.B(n_117),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2164),
.B(n_118),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2218),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2155),
.B(n_118),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2244),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2245),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2165),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2166),
.B(n_119),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_2244),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2183),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2221),
.B(n_121),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2211),
.B(n_122),
.Y(n_2374)
);

HB1xp67_ASAP7_75t_L g2375 ( 
.A(n_2270),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2312),
.B(n_2191),
.Y(n_2376)
);

AOI21x1_ASAP7_75t_L g2377 ( 
.A1(n_2346),
.A2(n_2163),
.B(n_2176),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2352),
.B(n_2132),
.Y(n_2378)
);

NAND4xp25_ASAP7_75t_L g2379 ( 
.A(n_2328),
.B(n_2200),
.C(n_2195),
.D(n_2194),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2250),
.A2(n_2235),
.B(n_2172),
.Y(n_2380)
);

OAI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2316),
.A2(n_2188),
.B1(n_2122),
.B2(n_2187),
.Y(n_2381)
);

CKINVDCx20_ASAP7_75t_R g2382 ( 
.A(n_2295),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2322),
.A2(n_2161),
.B(n_2209),
.Y(n_2383)
);

OAI21xp33_ASAP7_75t_L g2384 ( 
.A1(n_2262),
.A2(n_2273),
.B(n_2328),
.Y(n_2384)
);

OAI31xp33_ASAP7_75t_L g2385 ( 
.A1(n_2372),
.A2(n_2134),
.A3(n_2247),
.B(n_2224),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2311),
.A2(n_2209),
.B(n_2154),
.Y(n_2386)
);

OA21x2_ASAP7_75t_L g2387 ( 
.A1(n_2256),
.A2(n_2242),
.B(n_2167),
.Y(n_2387)
);

OAI211xp5_ASAP7_75t_L g2388 ( 
.A1(n_2371),
.A2(n_2185),
.B(n_2151),
.C(n_2098),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2259),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_2295),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_2296),
.B(n_2193),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2321),
.Y(n_2392)
);

OA21x2_ASAP7_75t_L g2393 ( 
.A1(n_2256),
.A2(n_2189),
.B(n_2156),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2264),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2321),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2358),
.A2(n_2343),
.B1(n_2318),
.B2(n_2367),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2265),
.Y(n_2397)
);

AOI22xp33_ASAP7_75t_L g2398 ( 
.A1(n_2365),
.A2(n_2184),
.B1(n_2153),
.B2(n_2129),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2253),
.B(n_2208),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2271),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2365),
.A2(n_2116),
.B1(n_2138),
.B2(n_2146),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2280),
.Y(n_2402)
);

AO21x2_ASAP7_75t_L g2403 ( 
.A1(n_2257),
.A2(n_2360),
.B(n_2277),
.Y(n_2403)
);

INVx4_ASAP7_75t_SL g2404 ( 
.A(n_2314),
.Y(n_2404)
);

AOI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2365),
.A2(n_2116),
.B(n_2097),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2286),
.B(n_2310),
.Y(n_2406)
);

BUFx3_ASAP7_75t_L g2407 ( 
.A(n_2314),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2352),
.B(n_2115),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_SL g2409 ( 
.A1(n_2368),
.A2(n_2219),
.B1(n_2140),
.B2(n_2091),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_SL g2410 ( 
.A1(n_2368),
.A2(n_2177),
.B1(n_2131),
.B2(n_2181),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2310),
.B(n_2210),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2368),
.B(n_2223),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2346),
.Y(n_2413)
);

AO31x2_ASAP7_75t_L g2414 ( 
.A1(n_2367),
.A2(n_124),
.A3(n_122),
.B(n_123),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2321),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2255),
.B(n_2168),
.Y(n_2416)
);

AOI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2370),
.A2(n_2160),
.B(n_2127),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_L g2418 ( 
.A(n_2352),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2281),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2283),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2358),
.A2(n_2203),
.B1(n_2199),
.B2(n_2171),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2338),
.B(n_125),
.Y(n_2422)
);

BUFx2_ASAP7_75t_L g2423 ( 
.A(n_2346),
.Y(n_2423)
);

OAI21xp33_ASAP7_75t_L g2424 ( 
.A1(n_2369),
.A2(n_125),
.B(n_126),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2321),
.Y(n_2425)
);

OAI221xp5_ASAP7_75t_L g2426 ( 
.A1(n_2369),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_2426)
);

OAI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_2326),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_2427)
);

INVxp67_ASAP7_75t_SL g2428 ( 
.A(n_2342),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2284),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2340),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2266),
.A2(n_2277),
.B(n_2339),
.Y(n_2431)
);

AO21x2_ASAP7_75t_L g2432 ( 
.A1(n_2266),
.A2(n_1325),
.B(n_1302),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2340),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2252),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2255),
.B(n_2261),
.Y(n_2435)
);

OAI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2254),
.A2(n_134),
.B(n_131),
.C(n_133),
.Y(n_2436)
);

A2O1A1Ixp33_ASAP7_75t_L g2437 ( 
.A1(n_2332),
.A2(n_137),
.B(n_134),
.C(n_136),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2258),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2318),
.A2(n_136),
.B(n_137),
.Y(n_2439)
);

OAI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2307),
.A2(n_145),
.B1(n_139),
.B2(n_142),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2340),
.Y(n_2441)
);

OAI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2373),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.C(n_149),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2340),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2368),
.B(n_146),
.Y(n_2444)
);

OAI211xp5_ASAP7_75t_SL g2445 ( 
.A1(n_2327),
.A2(n_152),
.B(n_147),
.C(n_151),
.Y(n_2445)
);

OAI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2330),
.A2(n_2362),
.B1(n_2344),
.B2(n_2268),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2296),
.Y(n_2447)
);

AO31x2_ASAP7_75t_L g2448 ( 
.A1(n_2309),
.A2(n_2324),
.A3(n_2332),
.B(n_2364),
.Y(n_2448)
);

OAI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2359),
.A2(n_2361),
.B(n_2355),
.Y(n_2449)
);

AND4x1_ASAP7_75t_L g2450 ( 
.A(n_2359),
.B(n_157),
.C(n_153),
.D(n_155),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2279),
.Y(n_2451)
);

AO21x2_ASAP7_75t_L g2452 ( 
.A1(n_2278),
.A2(n_1340),
.B(n_1338),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2268),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2366),
.A2(n_158),
.B(n_159),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2348),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2330),
.B(n_932),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2348),
.B(n_159),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2336),
.A2(n_160),
.B(n_162),
.Y(n_2458)
);

NAND3xp33_ASAP7_75t_L g2459 ( 
.A(n_2336),
.B(n_163),
.C(n_164),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2348),
.Y(n_2460)
);

A2O1A1Ixp33_ASAP7_75t_L g2461 ( 
.A1(n_2361),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2338),
.B(n_167),
.Y(n_2462)
);

AOI21xp33_ASAP7_75t_L g2463 ( 
.A1(n_2341),
.A2(n_168),
.B(n_169),
.Y(n_2463)
);

INVx4_ASAP7_75t_L g2464 ( 
.A(n_2349),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2329),
.B(n_170),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2251),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2260),
.Y(n_2467)
);

NAND2x1_ASAP7_75t_L g2468 ( 
.A(n_2274),
.B(n_170),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2261),
.B(n_171),
.Y(n_2469)
);

INVx5_ASAP7_75t_L g2470 ( 
.A(n_2337),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2292),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_2337),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2297),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2270),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2292),
.Y(n_2475)
);

AO21x2_ASAP7_75t_L g2476 ( 
.A1(n_2278),
.A2(n_1340),
.B(n_1338),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2345),
.B(n_172),
.C(n_173),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2289),
.Y(n_2478)
);

INVxp67_ASAP7_75t_L g2479 ( 
.A(n_2351),
.Y(n_2479)
);

INVx4_ASAP7_75t_L g2480 ( 
.A(n_2349),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_SL g2481 ( 
.A1(n_2355),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2260),
.Y(n_2482)
);

BUFx2_ASAP7_75t_L g2483 ( 
.A(n_2334),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2276),
.B(n_175),
.Y(n_2484)
);

HB1xp67_ASAP7_75t_L g2485 ( 
.A(n_2353),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2276),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2317),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2389),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2382),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2406),
.B(n_2274),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2394),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_2413),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2423),
.Y(n_2493)
);

BUFx3_ASAP7_75t_L g2494 ( 
.A(n_2390),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2470),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2397),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2390),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2470),
.Y(n_2498)
);

INVx5_ASAP7_75t_L g2499 ( 
.A(n_2418),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2400),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2402),
.Y(n_2501)
);

NAND4xp25_ASAP7_75t_L g2502 ( 
.A(n_2384),
.B(n_2341),
.C(n_2303),
.D(n_2306),
.Y(n_2502)
);

NAND4xp25_ASAP7_75t_L g2503 ( 
.A(n_2380),
.B(n_2304),
.C(n_2347),
.D(n_2354),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2419),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2390),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2470),
.B(n_2274),
.Y(n_2506)
);

OAI31xp33_ASAP7_75t_L g2507 ( 
.A1(n_2388),
.A2(n_2351),
.A3(n_2325),
.B(n_2305),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2472),
.B(n_2300),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2420),
.Y(n_2509)
);

AO21x2_ASAP7_75t_L g2510 ( 
.A1(n_2403),
.A2(n_2263),
.B(n_2325),
.Y(n_2510)
);

AND2x4_ASAP7_75t_L g2511 ( 
.A(n_2470),
.B(n_2263),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_L g2512 ( 
.A(n_2409),
.B(n_2354),
.C(n_2320),
.Y(n_2512)
);

BUFx2_ASAP7_75t_L g2513 ( 
.A(n_2404),
.Y(n_2513)
);

NAND4xp25_ASAP7_75t_SL g2514 ( 
.A(n_2380),
.B(n_2249),
.C(n_2347),
.D(n_2299),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2446),
.B(n_2376),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2428),
.B(n_2305),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2464),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2404),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2375),
.B(n_2290),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2435),
.B(n_2285),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2443),
.B(n_2285),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_2483),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2429),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2434),
.Y(n_2524)
);

BUFx2_ASAP7_75t_L g2525 ( 
.A(n_2404),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2438),
.Y(n_2526)
);

BUFx2_ASAP7_75t_L g2527 ( 
.A(n_2487),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2447),
.Y(n_2528)
);

OAI322xp33_ASAP7_75t_L g2529 ( 
.A1(n_2396),
.A2(n_2350),
.A3(n_2288),
.B1(n_2353),
.B2(n_2291),
.C1(n_2331),
.C2(n_2282),
.Y(n_2529)
);

OR2x6_ASAP7_75t_L g2530 ( 
.A(n_2468),
.B(n_2439),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2464),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2443),
.B(n_2323),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2480),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2478),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2480),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2418),
.B(n_2319),
.Y(n_2536)
);

INVxp67_ASAP7_75t_L g2537 ( 
.A(n_2378),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2418),
.B(n_2333),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2392),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2395),
.B(n_2313),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2473),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2415),
.B(n_2313),
.Y(n_2542)
);

CKINVDCx20_ASAP7_75t_R g2543 ( 
.A(n_2407),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2425),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2485),
.Y(n_2545)
);

INVx1_ASAP7_75t_SL g2546 ( 
.A(n_2457),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2430),
.Y(n_2547)
);

INVx1_ASAP7_75t_SL g2548 ( 
.A(n_2457),
.Y(n_2548)
);

OR2x2_ASAP7_75t_L g2549 ( 
.A(n_2474),
.B(n_2287),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2433),
.B(n_2275),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2441),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2484),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_2403),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2405),
.A2(n_2301),
.B(n_2333),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2379),
.A2(n_2333),
.B1(n_2300),
.B2(n_2335),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2455),
.B(n_2275),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2465),
.A2(n_2263),
.B(n_2309),
.Y(n_2557)
);

INVx5_ASAP7_75t_SL g2558 ( 
.A(n_2432),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2460),
.B(n_2287),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2431),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2453),
.B(n_2269),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2479),
.B(n_2448),
.Y(n_2562)
);

OA21x2_ASAP7_75t_L g2563 ( 
.A1(n_2376),
.A2(n_2324),
.B(n_2298),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2466),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_2486),
.B(n_2301),
.Y(n_2565)
);

OAI21xp33_ASAP7_75t_L g2566 ( 
.A1(n_2379),
.A2(n_2398),
.B(n_2386),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2414),
.Y(n_2567)
);

AOI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2396),
.A2(n_2308),
.B1(n_2374),
.B2(n_2248),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2431),
.Y(n_2569)
);

INVx5_ASAP7_75t_SL g2570 ( 
.A(n_2432),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2471),
.B(n_2269),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2475),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2482),
.B(n_2272),
.Y(n_2573)
);

AOI211xp5_ASAP7_75t_L g2574 ( 
.A1(n_2405),
.A2(n_2374),
.B(n_2363),
.C(n_2298),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2467),
.B(n_2272),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2492),
.Y(n_2576)
);

INVx3_ASAP7_75t_SL g2577 ( 
.A(n_2499),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2506),
.B(n_2448),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2492),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2490),
.B(n_2448),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2545),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2522),
.B(n_2465),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2507),
.B(n_2385),
.Y(n_2583)
);

OR2x2_ASAP7_75t_L g2584 ( 
.A(n_2493),
.B(n_2451),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2490),
.B(n_2467),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2506),
.B(n_2411),
.Y(n_2586)
);

NOR2x1_ASAP7_75t_SL g2587 ( 
.A(n_2530),
.B(n_2436),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2574),
.B(n_2381),
.Y(n_2588)
);

HB1xp67_ASAP7_75t_L g2589 ( 
.A(n_2493),
.Y(n_2589)
);

NAND2x1_ASAP7_75t_L g2590 ( 
.A(n_2511),
.B(n_2469),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2516),
.B(n_2399),
.Y(n_2591)
);

OR2x2_ASAP7_75t_L g2592 ( 
.A(n_2502),
.B(n_2391),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2546),
.B(n_2412),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2488),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2488),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2516),
.B(n_2416),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2508),
.B(n_2412),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2535),
.B(n_2393),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2535),
.B(n_2393),
.Y(n_2599)
);

NOR4xp25_ASAP7_75t_SL g2600 ( 
.A(n_2527),
.B(n_2456),
.C(n_2442),
.D(n_2463),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2548),
.B(n_2444),
.Y(n_2601)
);

CKINVDCx20_ASAP7_75t_R g2602 ( 
.A(n_2543),
.Y(n_2602)
);

NOR4xp25_ASAP7_75t_SL g2603 ( 
.A(n_2527),
.B(n_2442),
.C(n_2463),
.D(n_2426),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2495),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2517),
.B(n_2387),
.Y(n_2605)
);

NAND2x1p5_ASAP7_75t_L g2606 ( 
.A(n_2499),
.B(n_2450),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2517),
.B(n_2387),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2495),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2498),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2498),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2513),
.B(n_2459),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2491),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2519),
.B(n_2444),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2491),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2503),
.B(n_2449),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2496),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2496),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2500),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_2499),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2531),
.B(n_2449),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2566),
.B(n_2408),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2519),
.B(n_2414),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2549),
.B(n_2414),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2513),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2514),
.A2(n_2386),
.B1(n_2383),
.B2(n_2385),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2531),
.B(n_2267),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2533),
.B(n_2267),
.Y(n_2627)
);

INVx1_ASAP7_75t_SL g2628 ( 
.A(n_2489),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2500),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2552),
.B(n_2497),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2501),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2512),
.A2(n_2383),
.B1(n_2424),
.B2(n_2439),
.Y(n_2632)
);

BUFx3_ASAP7_75t_L g2633 ( 
.A(n_2489),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2501),
.Y(n_2634)
);

AO21x2_ASAP7_75t_L g2635 ( 
.A1(n_2560),
.A2(n_2454),
.B(n_2427),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2533),
.B(n_2308),
.Y(n_2636)
);

NOR2xp67_ASAP7_75t_L g2637 ( 
.A(n_2499),
.B(n_2422),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2552),
.B(n_2454),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2521),
.B(n_2315),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2552),
.B(n_2458),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2504),
.Y(n_2641)
);

INVxp67_ASAP7_75t_L g2642 ( 
.A(n_2518),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2521),
.B(n_2315),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2532),
.B(n_2540),
.Y(n_2644)
);

OR2x6_ASAP7_75t_L g2645 ( 
.A(n_2518),
.B(n_2477),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2560),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2494),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2549),
.B(n_2293),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2532),
.B(n_2294),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2568),
.B(n_2417),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2515),
.B(n_2461),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2569),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2572),
.B(n_2437),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2504),
.Y(n_2654)
);

NAND2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2525),
.B(n_2401),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2494),
.Y(n_2656)
);

BUFx3_ASAP7_75t_L g2657 ( 
.A(n_2525),
.Y(n_2657)
);

XOR2x2_ASAP7_75t_L g2658 ( 
.A(n_2583),
.B(n_2621),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2657),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2589),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2633),
.B(n_2505),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_2602),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2628),
.B(n_2537),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2633),
.B(n_2505),
.Y(n_2664)
);

XOR2xp5_ASAP7_75t_L g2665 ( 
.A(n_2602),
.B(n_2421),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2657),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2586),
.B(n_2499),
.Y(n_2667)
);

XOR2x2_ASAP7_75t_L g2668 ( 
.A(n_2583),
.B(n_2462),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2624),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2577),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2655),
.A2(n_2530),
.B1(n_2536),
.B2(n_2538),
.Y(n_2671)
);

XOR2xp5_ASAP7_75t_L g2672 ( 
.A(n_2615),
.B(n_2421),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2586),
.B(n_2530),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2646),
.Y(n_2674)
);

NAND3xp33_ASAP7_75t_L g2675 ( 
.A(n_2603),
.B(n_2530),
.C(n_2562),
.Y(n_2675)
);

XOR2x2_ASAP7_75t_L g2676 ( 
.A(n_2621),
.B(n_2426),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2576),
.Y(n_2677)
);

NAND4xp75_ASAP7_75t_L g2678 ( 
.A(n_2637),
.B(n_2588),
.C(n_2650),
.D(n_2599),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2576),
.Y(n_2679)
);

INVx2_ASAP7_75t_SL g2680 ( 
.A(n_2577),
.Y(n_2680)
);

NAND4xp75_ASAP7_75t_L g2681 ( 
.A(n_2598),
.B(n_2563),
.C(n_2554),
.D(n_2569),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2611),
.B(n_2539),
.Y(n_2682)
);

AOI22xp5_ASAP7_75t_L g2683 ( 
.A1(n_2655),
.A2(n_2410),
.B1(n_2510),
.B2(n_2555),
.Y(n_2683)
);

NAND4xp75_ASAP7_75t_L g2684 ( 
.A(n_2598),
.B(n_2563),
.C(n_2539),
.D(n_2547),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2591),
.B(n_2499),
.Y(n_2685)
);

NOR4xp25_ASAP7_75t_L g2686 ( 
.A(n_2625),
.B(n_2529),
.C(n_2562),
.D(n_2445),
.Y(n_2686)
);

NAND4xp75_ASAP7_75t_SL g2687 ( 
.A(n_2591),
.B(n_2563),
.C(n_2377),
.D(n_2542),
.Y(n_2687)
);

XOR2xp5_ASAP7_75t_L g2688 ( 
.A(n_2606),
.B(n_2481),
.Y(n_2688)
);

INVx4_ASAP7_75t_L g2689 ( 
.A(n_2619),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2652),
.Y(n_2690)
);

NAND2xp33_ASAP7_75t_R g2691 ( 
.A(n_2600),
.B(n_2553),
.Y(n_2691)
);

NAND4xp75_ASAP7_75t_L g2692 ( 
.A(n_2599),
.B(n_2563),
.C(n_2544),
.D(n_2551),
.Y(n_2692)
);

XNOR2xp5_ASAP7_75t_L g2693 ( 
.A(n_2606),
.B(n_2440),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2596),
.B(n_2520),
.Y(n_2694)
);

NAND3xp33_ASAP7_75t_SL g2695 ( 
.A(n_2632),
.B(n_2553),
.C(n_2567),
.Y(n_2695)
);

NOR3xp33_ASAP7_75t_L g2696 ( 
.A(n_2630),
.B(n_2547),
.C(n_2544),
.Y(n_2696)
);

XNOR2xp5_ASAP7_75t_L g2697 ( 
.A(n_2596),
.B(n_2363),
.Y(n_2697)
);

AOI211xp5_ASAP7_75t_SL g2698 ( 
.A1(n_2642),
.A2(n_2511),
.B(n_2567),
.C(n_2551),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2578),
.Y(n_2699)
);

XOR2x2_ASAP7_75t_L g2700 ( 
.A(n_2587),
.B(n_2510),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2579),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2579),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2619),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2611),
.B(n_2564),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2644),
.B(n_2520),
.Y(n_2705)
);

INVxp33_ASAP7_75t_SL g2706 ( 
.A(n_2582),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2604),
.Y(n_2707)
);

NAND4xp75_ASAP7_75t_SL g2708 ( 
.A(n_2605),
.B(n_2542),
.C(n_2540),
.D(n_2550),
.Y(n_2708)
);

NOR3xp33_ASAP7_75t_SL g2709 ( 
.A(n_2638),
.B(n_2564),
.C(n_2541),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_SL g2710 ( 
.A(n_2611),
.B(n_2647),
.Y(n_2710)
);

NAND4xp75_ASAP7_75t_SL g2711 ( 
.A(n_2605),
.B(n_2550),
.C(n_2575),
.D(n_2561),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2585),
.B(n_2559),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2647),
.B(n_2541),
.Y(n_2713)
);

XOR2xp5_ASAP7_75t_L g2714 ( 
.A(n_2592),
.B(n_2528),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2578),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2578),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2644),
.B(n_2559),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2604),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2656),
.B(n_2509),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2677),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2677),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2679),
.Y(n_2722)
);

AOI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2658),
.A2(n_2635),
.B1(n_2645),
.B2(n_2651),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2662),
.B(n_2585),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2669),
.B(n_2656),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2667),
.B(n_2620),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2669),
.B(n_2620),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2679),
.Y(n_2728)
);

NOR2xp67_ASAP7_75t_L g2729 ( 
.A(n_2689),
.B(n_2584),
.Y(n_2729)
);

INVxp67_ASAP7_75t_L g2730 ( 
.A(n_2710),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2667),
.B(n_2580),
.Y(n_2731)
);

INVx1_ASAP7_75t_SL g2732 ( 
.A(n_2685),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2659),
.B(n_2581),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2659),
.B(n_2635),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2701),
.B(n_2584),
.Y(n_2735)
);

INVxp67_ASAP7_75t_SL g2736 ( 
.A(n_2691),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2699),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2685),
.B(n_2580),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2702),
.Y(n_2739)
);

INVxp67_ASAP7_75t_L g2740 ( 
.A(n_2673),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2666),
.B(n_2635),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2704),
.B(n_2660),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2699),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2699),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2674),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2707),
.Y(n_2746)
);

INVxp67_ASAP7_75t_SL g2747 ( 
.A(n_2691),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2716),
.Y(n_2748)
);

NAND2x1p5_ASAP7_75t_L g2749 ( 
.A(n_2680),
.B(n_2590),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2666),
.B(n_2593),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2686),
.B(n_2658),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2718),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2690),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2716),
.Y(n_2754)
);

NOR2x1p5_ASAP7_75t_L g2755 ( 
.A(n_2678),
.B(n_2663),
.Y(n_2755)
);

INVx1_ASAP7_75t_SL g2756 ( 
.A(n_2661),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2705),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2706),
.B(n_2601),
.Y(n_2758)
);

INVxp67_ASAP7_75t_L g2759 ( 
.A(n_2664),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2705),
.B(n_2607),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2668),
.B(n_2640),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2668),
.B(n_2645),
.Y(n_2762)
);

INVx2_ASAP7_75t_SL g2763 ( 
.A(n_2716),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2682),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2683),
.B(n_2653),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2717),
.Y(n_2766)
);

OAI31xp33_ASAP7_75t_L g2767 ( 
.A1(n_2751),
.A2(n_2675),
.A3(n_2688),
.B(n_2693),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2728),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2736),
.B(n_2697),
.Y(n_2769)
);

OAI22xp33_ASAP7_75t_SL g2770 ( 
.A1(n_2747),
.A2(n_2706),
.B1(n_2671),
.B2(n_2645),
.Y(n_2770)
);

BUFx2_ASAP7_75t_L g2771 ( 
.A(n_2749),
.Y(n_2771)
);

OAI21xp33_ASAP7_75t_L g2772 ( 
.A1(n_2762),
.A2(n_2676),
.B(n_2695),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2723),
.A2(n_2676),
.B1(n_2700),
.B2(n_2645),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2744),
.Y(n_2774)
);

AOI21xp33_ASAP7_75t_L g2775 ( 
.A1(n_2730),
.A2(n_2680),
.B(n_2714),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2754),
.Y(n_2776)
);

OAI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_2765),
.A2(n_2700),
.B1(n_2709),
.B2(n_2761),
.C(n_2672),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2749),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2749),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2724),
.B(n_2665),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2720),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2724),
.B(n_2694),
.Y(n_2782)
);

O2A1O1Ixp33_ASAP7_75t_L g2783 ( 
.A1(n_2765),
.A2(n_2709),
.B(n_2698),
.C(n_2670),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2720),
.Y(n_2784)
);

OAI21xp33_ASAP7_75t_L g2785 ( 
.A1(n_2758),
.A2(n_2712),
.B(n_2717),
.Y(n_2785)
);

INVx2_ASAP7_75t_SL g2786 ( 
.A(n_2735),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2735),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2721),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2760),
.Y(n_2789)
);

AOI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2755),
.A2(n_2681),
.B1(n_2692),
.B2(n_2684),
.Y(n_2790)
);

OR2x2_ASAP7_75t_L g2791 ( 
.A(n_2727),
.B(n_2613),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2763),
.Y(n_2792)
);

OAI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2756),
.A2(n_2597),
.B1(n_2613),
.B2(n_2670),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2729),
.A2(n_2696),
.B1(n_2510),
.B2(n_2607),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2722),
.A2(n_2689),
.B1(n_2703),
.B2(n_2594),
.Y(n_2795)
);

OAI22xp33_ASAP7_75t_L g2796 ( 
.A1(n_2734),
.A2(n_2622),
.B1(n_2623),
.B2(n_2687),
.Y(n_2796)
);

AOI211xp5_ASAP7_75t_L g2797 ( 
.A1(n_2732),
.A2(n_2713),
.B(n_2719),
.C(n_2703),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2763),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2737),
.Y(n_2799)
);

INVxp67_ASAP7_75t_L g2800 ( 
.A(n_2760),
.Y(n_2800)
);

AOI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2759),
.A2(n_2636),
.B1(n_2689),
.B2(n_2609),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2740),
.A2(n_2622),
.B1(n_2623),
.B2(n_2609),
.Y(n_2802)
);

XNOR2xp5_ASAP7_75t_L g2803 ( 
.A(n_2757),
.B(n_2711),
.Y(n_2803)
);

INVx2_ASAP7_75t_SL g2804 ( 
.A(n_2737),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2786),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2787),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2789),
.B(n_2766),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2782),
.B(n_2726),
.Y(n_2808)
);

OAI322xp33_ASAP7_75t_L g2809 ( 
.A1(n_2790),
.A2(n_2742),
.A3(n_2741),
.B1(n_2725),
.B2(n_2753),
.C1(n_2745),
.C2(n_2766),
.Y(n_2809)
);

OR2x6_ASAP7_75t_L g2810 ( 
.A(n_2771),
.B(n_2750),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2804),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2792),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2798),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2772),
.A2(n_2726),
.B1(n_2764),
.B2(n_2557),
.Y(n_2814)
);

OAI32xp33_ASAP7_75t_L g2815 ( 
.A1(n_2777),
.A2(n_2742),
.A3(n_2733),
.B1(n_2745),
.B2(n_2731),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2790),
.A2(n_2731),
.B1(n_2738),
.B2(n_2636),
.Y(n_2816)
);

INVxp67_ASAP7_75t_SL g2817 ( 
.A(n_2778),
.Y(n_2817)
);

NOR2x1_ASAP7_75t_L g2818 ( 
.A(n_2779),
.B(n_2743),
.Y(n_2818)
);

NAND2xp33_ASAP7_75t_SL g2819 ( 
.A(n_2780),
.B(n_2738),
.Y(n_2819)
);

XNOR2x1_ASAP7_75t_L g2820 ( 
.A(n_2803),
.B(n_2773),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2799),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2800),
.B(n_2743),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2774),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2776),
.B(n_2748),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2768),
.Y(n_2825)
);

AOI211x1_ASAP7_75t_SL g2826 ( 
.A1(n_2775),
.A2(n_2748),
.B(n_2715),
.C(n_2610),
.Y(n_2826)
);

INVxp67_ASAP7_75t_L g2827 ( 
.A(n_2769),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2791),
.B(n_2608),
.Y(n_2828)
);

OAI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2773),
.A2(n_2715),
.B1(n_2610),
.B2(n_2608),
.Y(n_2829)
);

OAI21xp33_ASAP7_75t_SL g2830 ( 
.A1(n_2794),
.A2(n_2708),
.B(n_2739),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2781),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2785),
.B(n_2746),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2801),
.B(n_2752),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2784),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2795),
.Y(n_2835)
);

INVx1_ASAP7_75t_SL g2836 ( 
.A(n_2793),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2808),
.Y(n_2837)
);

INVx1_ASAP7_75t_SL g2838 ( 
.A(n_2807),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2805),
.B(n_2797),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2816),
.B(n_2767),
.Y(n_2840)
);

OAI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2830),
.A2(n_2783),
.B(n_2796),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2818),
.Y(n_2842)
);

OAI21xp33_ASAP7_75t_L g2843 ( 
.A1(n_2820),
.A2(n_2836),
.B(n_2770),
.Y(n_2843)
);

OAI32xp33_ASAP7_75t_L g2844 ( 
.A1(n_2830),
.A2(n_2802),
.A3(n_2788),
.B1(n_2595),
.B2(n_2634),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2817),
.B(n_2795),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2810),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2810),
.B(n_2794),
.Y(n_2847)
);

OAI21xp5_ASAP7_75t_SL g2848 ( 
.A1(n_2826),
.A2(n_2614),
.B(n_2612),
.Y(n_2848)
);

O2A1O1Ixp33_ASAP7_75t_SL g2849 ( 
.A1(n_2835),
.A2(n_2617),
.B(n_2618),
.C(n_2616),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2828),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2811),
.B(n_2806),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2822),
.Y(n_2852)
);

INVx1_ASAP7_75t_SL g2853 ( 
.A(n_2810),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2834),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2824),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2809),
.B(n_2629),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2829),
.B(n_2834),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2812),
.B(n_2631),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2832),
.Y(n_2859)
);

OAI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2814),
.A2(n_2827),
.B1(n_2813),
.B2(n_2833),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2823),
.Y(n_2861)
);

INVx1_ASAP7_75t_SL g2862 ( 
.A(n_2853),
.Y(n_2862)
);

NOR3x1_ASAP7_75t_L g2863 ( 
.A(n_2841),
.B(n_2825),
.C(n_2821),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2859),
.B(n_2831),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2843),
.B(n_2815),
.Y(n_2865)
);

NOR3x1_ASAP7_75t_L g2866 ( 
.A(n_2840),
.B(n_2819),
.C(n_2654),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2845),
.Y(n_2867)
);

OAI211xp5_ASAP7_75t_L g2868 ( 
.A1(n_2856),
.A2(n_2641),
.B(n_2523),
.C(n_2524),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2846),
.B(n_2649),
.Y(n_2869)
);

NOR3x1_ASAP7_75t_L g2870 ( 
.A(n_2848),
.B(n_2523),
.C(n_2509),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2842),
.B(n_2524),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2838),
.B(n_2649),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_2857),
.Y(n_2873)
);

NOR2x1_ASAP7_75t_L g2874 ( 
.A(n_2847),
.B(n_2857),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2859),
.B(n_2526),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2854),
.B(n_2850),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2856),
.B(n_2626),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2839),
.B(n_2639),
.Y(n_2878)
);

NOR3xp33_ASAP7_75t_L g2879 ( 
.A(n_2860),
.B(n_2627),
.C(n_2626),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2837),
.B(n_2526),
.Y(n_2880)
);

OAI21xp5_ASAP7_75t_SL g2881 ( 
.A1(n_2873),
.A2(n_2852),
.B(n_2851),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2877),
.A2(n_2862),
.B1(n_2874),
.B2(n_2872),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2878),
.B(n_2861),
.Y(n_2883)
);

NOR4xp25_ASAP7_75t_L g2884 ( 
.A(n_2876),
.B(n_2849),
.C(n_2855),
.D(n_2858),
.Y(n_2884)
);

O2A1O1Ixp33_ASAP7_75t_L g2885 ( 
.A1(n_2865),
.A2(n_2844),
.B(n_2849),
.C(n_2511),
.Y(n_2885)
);

AO22x2_ASAP7_75t_L g2886 ( 
.A1(n_2868),
.A2(n_2534),
.B1(n_2528),
.B2(n_2511),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2879),
.A2(n_2627),
.B1(n_2534),
.B2(n_2557),
.Y(n_2887)
);

A2O1A1Ixp33_ASAP7_75t_L g2888 ( 
.A1(n_2875),
.A2(n_2572),
.B(n_2565),
.C(n_2648),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2864),
.B(n_2639),
.Y(n_2889)
);

AND3x1_ASAP7_75t_L g2890 ( 
.A(n_2869),
.B(n_2643),
.C(n_2575),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2871),
.A2(n_2557),
.B(n_2643),
.Y(n_2891)
);

OAI211xp5_ASAP7_75t_SL g2892 ( 
.A1(n_2867),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2892)
);

OAI21xp33_ASAP7_75t_SL g2893 ( 
.A1(n_2871),
.A2(n_2880),
.B(n_2870),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2884),
.B(n_2863),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2886),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2890),
.A2(n_2565),
.B1(n_2573),
.B2(n_2561),
.Y(n_2896)
);

OAI221xp5_ASAP7_75t_L g2897 ( 
.A1(n_2881),
.A2(n_2866),
.B1(n_2573),
.B2(n_2556),
.C(n_2571),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2889),
.Y(n_2898)
);

AOI22xp33_ASAP7_75t_L g2899 ( 
.A1(n_2882),
.A2(n_2558),
.B1(n_2570),
.B2(n_2565),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2883),
.A2(n_2565),
.B1(n_2556),
.B2(n_2571),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2893),
.Y(n_2901)
);

OAI22x1_ASAP7_75t_L g2902 ( 
.A1(n_2887),
.A2(n_2357),
.B1(n_2302),
.B2(n_2335),
.Y(n_2902)
);

O2A1O1Ixp33_ASAP7_75t_SL g2903 ( 
.A1(n_2885),
.A2(n_2558),
.B(n_2570),
.C(n_2356),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2892),
.Y(n_2904)
);

AOI22x1_ASAP7_75t_L g2905 ( 
.A1(n_2891),
.A2(n_2888),
.B1(n_2357),
.B2(n_2570),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2886),
.Y(n_2906)
);

AOI221xp5_ASAP7_75t_L g2907 ( 
.A1(n_2894),
.A2(n_2570),
.B1(n_2558),
.B2(n_2302),
.C(n_2452),
.Y(n_2907)
);

AOI221xp5_ASAP7_75t_L g2908 ( 
.A1(n_2903),
.A2(n_2558),
.B1(n_2302),
.B2(n_2452),
.C(n_2476),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2901),
.B(n_2476),
.Y(n_2909)
);

AOI211xp5_ASAP7_75t_L g2910 ( 
.A1(n_2901),
.A2(n_181),
.B(n_177),
.C(n_180),
.Y(n_2910)
);

AOI221xp5_ASAP7_75t_L g2911 ( 
.A1(n_2897),
.A2(n_2899),
.B1(n_2895),
.B2(n_2906),
.C(n_2904),
.Y(n_2911)
);

NOR4xp75_ASAP7_75t_L g2912 ( 
.A(n_2900),
.B(n_183),
.C(n_180),
.D(n_181),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2905),
.Y(n_2913)
);

NOR4xp25_ASAP7_75t_L g2914 ( 
.A(n_2898),
.B(n_2896),
.C(n_2902),
.D(n_186),
.Y(n_2914)
);

NAND4xp25_ASAP7_75t_SL g2915 ( 
.A(n_2894),
.B(n_184),
.C(n_185),
.D(n_187),
.Y(n_2915)
);

O2A1O1Ixp5_ASAP7_75t_L g2916 ( 
.A1(n_2895),
.A2(n_185),
.B(n_187),
.C(n_188),
.Y(n_2916)
);

AOI221xp5_ASAP7_75t_L g2917 ( 
.A1(n_2894),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.C(n_192),
.Y(n_2917)
);

NAND3xp33_ASAP7_75t_L g2918 ( 
.A(n_2901),
.B(n_191),
.C(n_192),
.Y(n_2918)
);

AOI21xp33_ASAP7_75t_L g2919 ( 
.A1(n_2901),
.A2(n_193),
.B(n_194),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2894),
.A2(n_193),
.B(n_194),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_R g2921 ( 
.A(n_2894),
.B(n_195),
.Y(n_2921)
);

OAI211xp5_ASAP7_75t_SL g2922 ( 
.A1(n_2894),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_2922)
);

NOR3xp33_ASAP7_75t_L g2923 ( 
.A(n_2894),
.B(n_196),
.C(n_197),
.Y(n_2923)
);

AOI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2914),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.C(n_204),
.Y(n_2924)
);

NOR2x1p5_ASAP7_75t_L g2925 ( 
.A(n_2918),
.B(n_201),
.Y(n_2925)
);

NAND3xp33_ASAP7_75t_L g2926 ( 
.A(n_2911),
.B(n_204),
.C(n_205),
.Y(n_2926)
);

OAI221xp5_ASAP7_75t_SL g2927 ( 
.A1(n_2913),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.C(n_209),
.Y(n_2927)
);

AOI211xp5_ASAP7_75t_SL g2928 ( 
.A1(n_2920),
.A2(n_207),
.B(n_209),
.C(n_210),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2923),
.A2(n_2335),
.B1(n_211),
.B2(n_213),
.Y(n_2929)
);

NOR5xp2_ASAP7_75t_L g2930 ( 
.A(n_2922),
.B(n_210),
.C(n_213),
.D(n_214),
.E(n_215),
.Y(n_2930)
);

O2A1O1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2916),
.A2(n_215),
.B(n_216),
.C(n_217),
.Y(n_2931)
);

AOI211xp5_ASAP7_75t_L g2932 ( 
.A1(n_2915),
.A2(n_218),
.B(n_219),
.C(n_221),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2909),
.Y(n_2933)
);

AOI211x1_ASAP7_75t_L g2934 ( 
.A1(n_2919),
.A2(n_218),
.B(n_219),
.C(n_221),
.Y(n_2934)
);

AOI221xp5_ASAP7_75t_L g2935 ( 
.A1(n_2921),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.C(n_226),
.Y(n_2935)
);

NOR3xp33_ASAP7_75t_SL g2936 ( 
.A(n_2917),
.B(n_2912),
.C(n_2910),
.Y(n_2936)
);

AOI221xp5_ASAP7_75t_L g2937 ( 
.A1(n_2907),
.A2(n_223),
.B1(n_227),
.B2(n_1306),
.C(n_1301),
.Y(n_2937)
);

AOI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2908),
.A2(n_227),
.B1(n_1301),
.B2(n_932),
.C(n_1328),
.Y(n_2938)
);

NAND3xp33_ASAP7_75t_L g2939 ( 
.A(n_2928),
.B(n_1328),
.C(n_1304),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2931),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2924),
.B(n_1328),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2926),
.A2(n_2927),
.B1(n_2932),
.B2(n_2934),
.Y(n_2942)
);

NAND3x1_ASAP7_75t_L g2943 ( 
.A(n_2935),
.B(n_228),
.C(n_229),
.Y(n_2943)
);

NAND4xp25_ASAP7_75t_L g2944 ( 
.A(n_2938),
.B(n_2930),
.C(n_2937),
.D(n_2933),
.Y(n_2944)
);

AOI22x1_ASAP7_75t_L g2945 ( 
.A1(n_2925),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2933),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2936),
.A2(n_1005),
.B1(n_894),
.B2(n_1161),
.Y(n_2947)
);

NOR2x1_ASAP7_75t_L g2948 ( 
.A(n_2929),
.B(n_1180),
.Y(n_2948)
);

NAND3x1_ASAP7_75t_SL g2949 ( 
.A(n_2924),
.B(n_239),
.C(n_240),
.Y(n_2949)
);

NAND3xp33_ASAP7_75t_SL g2950 ( 
.A(n_2924),
.B(n_243),
.C(n_245),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2940),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2949),
.Y(n_2952)
);

NAND5xp2_ASAP7_75t_L g2953 ( 
.A(n_2942),
.B(n_251),
.C(n_252),
.D(n_253),
.E(n_255),
.Y(n_2953)
);

INVx3_ASAP7_75t_SL g2954 ( 
.A(n_2946),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2945),
.Y(n_2955)
);

NAND3xp33_ASAP7_75t_L g2956 ( 
.A(n_2939),
.B(n_1347),
.C(n_1304),
.Y(n_2956)
);

NAND4xp75_ASAP7_75t_L g2957 ( 
.A(n_2948),
.B(n_259),
.C(n_260),
.D(n_261),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2943),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2950),
.A2(n_2944),
.B1(n_2941),
.B2(n_2947),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2940),
.B(n_265),
.Y(n_2960)
);

NOR3xp33_ASAP7_75t_L g2961 ( 
.A(n_2940),
.B(n_900),
.C(n_876),
.Y(n_2961)
);

INVxp33_ASAP7_75t_SL g2962 ( 
.A(n_2960),
.Y(n_2962)
);

NOR3xp33_ASAP7_75t_L g2963 ( 
.A(n_2951),
.B(n_2958),
.C(n_2952),
.Y(n_2963)
);

OAI221xp5_ASAP7_75t_L g2964 ( 
.A1(n_2954),
.A2(n_1249),
.B1(n_269),
.B2(n_277),
.C(n_278),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2955),
.B(n_266),
.Y(n_2965)
);

OAI311xp33_ASAP7_75t_L g2966 ( 
.A1(n_2959),
.A2(n_2956),
.A3(n_2961),
.B1(n_2957),
.C1(n_2953),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2954),
.B(n_279),
.Y(n_2967)
);

NOR2x1p5_ASAP7_75t_L g2968 ( 
.A(n_2957),
.B(n_281),
.Y(n_2968)
);

OAI211xp5_ASAP7_75t_L g2969 ( 
.A1(n_2951),
.A2(n_285),
.B(n_286),
.C(n_289),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2957),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2960),
.Y(n_2971)
);

NOR4xp25_ASAP7_75t_L g2972 ( 
.A(n_2951),
.B(n_291),
.C(n_292),
.D(n_295),
.Y(n_2972)
);

OAI211xp5_ASAP7_75t_L g2973 ( 
.A1(n_2951),
.A2(n_297),
.B(n_300),
.C(n_307),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2960),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2968),
.Y(n_2975)
);

AOI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2963),
.A2(n_1005),
.B1(n_894),
.B2(n_932),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2965),
.Y(n_2977)
);

XNOR2xp5_ASAP7_75t_L g2978 ( 
.A(n_2962),
.B(n_2970),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_L g2979 ( 
.A1(n_2971),
.A2(n_932),
.B1(n_1005),
.B2(n_957),
.Y(n_2979)
);

XOR2xp5_ASAP7_75t_L g2980 ( 
.A(n_2967),
.B(n_308),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2974),
.Y(n_2981)
);

NAND4xp75_ASAP7_75t_L g2982 ( 
.A(n_2966),
.B(n_310),
.C(n_311),
.D(n_313),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2964),
.Y(n_2983)
);

OAI22x1_ASAP7_75t_L g2984 ( 
.A1(n_2980),
.A2(n_2972),
.B1(n_2973),
.B2(n_2969),
.Y(n_2984)
);

AOI22xp5_ASAP7_75t_L g2985 ( 
.A1(n_2982),
.A2(n_1005),
.B1(n_894),
.B2(n_932),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2981),
.A2(n_1087),
.B1(n_1093),
.B2(n_1097),
.Y(n_2986)
);

OAI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2975),
.A2(n_1097),
.B1(n_1027),
.B2(n_1029),
.Y(n_2987)
);

OAI221xp5_ASAP7_75t_L g2988 ( 
.A1(n_2978),
.A2(n_2977),
.B1(n_2983),
.B2(n_2979),
.C(n_2976),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2982),
.Y(n_2989)
);

OAI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2982),
.A2(n_1097),
.B1(n_1029),
.B2(n_1039),
.Y(n_2990)
);

AOI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2982),
.A2(n_1005),
.B1(n_894),
.B2(n_947),
.Y(n_2991)
);

OAI22x1_ASAP7_75t_L g2992 ( 
.A1(n_2980),
.A2(n_317),
.B1(n_323),
.B2(n_325),
.Y(n_2992)
);

HB1xp67_ASAP7_75t_L g2993 ( 
.A(n_2982),
.Y(n_2993)
);

OAI22x1_ASAP7_75t_L g2994 ( 
.A1(n_2980),
.A2(n_328),
.B1(n_335),
.B2(n_336),
.Y(n_2994)
);

HB1xp67_ASAP7_75t_L g2995 ( 
.A(n_2982),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2982),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2977),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_SL g2998 ( 
.A1(n_2977),
.A2(n_894),
.B1(n_1170),
.B2(n_947),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2982),
.A2(n_894),
.B1(n_963),
.B2(n_958),
.Y(n_2999)
);

OAI22x1_ASAP7_75t_L g3000 ( 
.A1(n_2980),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2982),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2977),
.Y(n_3002)
);

BUFx2_ASAP7_75t_L g3003 ( 
.A(n_2977),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2977),
.Y(n_3004)
);

OAI31xp33_ASAP7_75t_L g3005 ( 
.A1(n_3003),
.A2(n_340),
.A3(n_343),
.B(n_346),
.Y(n_3005)
);

BUFx2_ASAP7_75t_L g3006 ( 
.A(n_2993),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_2997),
.B(n_350),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2995),
.Y(n_3008)
);

OAI31xp33_ASAP7_75t_L g3009 ( 
.A1(n_3002),
.A2(n_352),
.A3(n_354),
.B(n_362),
.Y(n_3009)
);

AOI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_3004),
.A2(n_2989),
.B1(n_2996),
.B2(n_3001),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2984),
.Y(n_3011)
);

AOI22xp33_ASAP7_75t_SL g3012 ( 
.A1(n_2988),
.A2(n_894),
.B1(n_957),
.B2(n_947),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2991),
.A2(n_957),
.B1(n_958),
.B2(n_963),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2985),
.A2(n_957),
.B1(n_958),
.B2(n_963),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_2999),
.A2(n_947),
.B1(n_957),
.B2(n_958),
.Y(n_3015)
);

AOI31xp33_ASAP7_75t_L g3016 ( 
.A1(n_2990),
.A2(n_367),
.A3(n_371),
.B(n_376),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2992),
.Y(n_3017)
);

OAI31xp33_ASAP7_75t_SL g3018 ( 
.A1(n_2998),
.A2(n_379),
.A3(n_380),
.B(n_381),
.Y(n_3018)
);

AOI22xp5_ASAP7_75t_L g3019 ( 
.A1(n_2994),
.A2(n_947),
.B1(n_963),
.B2(n_958),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_3000),
.A2(n_963),
.B1(n_1059),
.B2(n_1070),
.Y(n_3020)
);

AOI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_2986),
.A2(n_918),
.B1(n_870),
.B2(n_1341),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2987),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_3003),
.B(n_382),
.Y(n_3023)
);

A2O1A1Ixp33_ASAP7_75t_SL g3024 ( 
.A1(n_2997),
.A2(n_918),
.B(n_870),
.C(n_1067),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_3003),
.B(n_383),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2997),
.A2(n_1351),
.B1(n_1347),
.B2(n_1304),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2992),
.Y(n_3027)
);

BUFx2_ASAP7_75t_L g3028 ( 
.A(n_3003),
.Y(n_3028)
);

OAI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2997),
.A2(n_1351),
.B1(n_1347),
.B2(n_1070),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_3003),
.A2(n_1059),
.B1(n_1074),
.B2(n_1071),
.Y(n_3030)
);

OAI31xp33_ASAP7_75t_L g3031 ( 
.A1(n_3003),
.A2(n_385),
.A3(n_386),
.B(n_391),
.Y(n_3031)
);

OAI31xp33_ASAP7_75t_L g3032 ( 
.A1(n_3003),
.A2(n_392),
.A3(n_393),
.B(n_394),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_3003),
.B(n_396),
.Y(n_3033)
);

NAND5xp2_ASAP7_75t_L g3034 ( 
.A(n_3010),
.B(n_398),
.C(n_400),
.D(n_403),
.E(n_406),
.Y(n_3034)
);

NAND4xp25_ASAP7_75t_SL g3035 ( 
.A(n_3023),
.B(n_412),
.C(n_414),
.D(n_415),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_3028),
.A2(n_1351),
.B1(n_918),
.B2(n_870),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_3006),
.A2(n_1050),
.B1(n_1043),
.B2(n_1046),
.Y(n_3037)
);

NAND4xp25_ASAP7_75t_L g3038 ( 
.A(n_3011),
.B(n_3008),
.C(n_3033),
.D(n_3025),
.Y(n_3038)
);

AOI322xp5_ASAP7_75t_L g3039 ( 
.A1(n_3017),
.A2(n_416),
.A3(n_418),
.B1(n_419),
.B2(n_1210),
.C1(n_1237),
.C2(n_1208),
.Y(n_3039)
);

NAND4xp25_ASAP7_75t_L g3040 ( 
.A(n_3027),
.B(n_876),
.C(n_900),
.D(n_1067),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_3019),
.A2(n_3013),
.B1(n_3014),
.B2(n_3016),
.Y(n_3041)
);

OAI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_3012),
.A2(n_1074),
.B(n_1071),
.Y(n_3042)
);

AOI221xp5_ASAP7_75t_L g3043 ( 
.A1(n_3026),
.A2(n_928),
.B1(n_1341),
.B2(n_1180),
.C(n_1295),
.Y(n_3043)
);

AOI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_3022),
.A2(n_1043),
.B1(n_1050),
.B2(n_1039),
.Y(n_3044)
);

O2A1O1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_3024),
.A2(n_1067),
.B(n_1084),
.C(n_1101),
.Y(n_3045)
);

NAND4xp25_ASAP7_75t_L g3046 ( 
.A(n_3018),
.B(n_876),
.C(n_900),
.D(n_1135),
.Y(n_3046)
);

A2O1A1Ixp33_ASAP7_75t_L g3047 ( 
.A1(n_3005),
.A2(n_1135),
.B(n_1101),
.C(n_1062),
.Y(n_3047)
);

NOR4xp25_ASAP7_75t_L g3048 ( 
.A(n_3015),
.B(n_1135),
.C(n_1084),
.D(n_1101),
.Y(n_3048)
);

NAND4xp25_ASAP7_75t_SL g3049 ( 
.A(n_3031),
.B(n_1046),
.C(n_1048),
.D(n_1019),
.Y(n_3049)
);

AOI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3007),
.A2(n_1278),
.B1(n_1295),
.B2(n_1196),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_3032),
.A2(n_1086),
.B1(n_1080),
.B2(n_1019),
.Y(n_3051)
);

AO22x2_ASAP7_75t_L g3052 ( 
.A1(n_3029),
.A2(n_3009),
.B1(n_3021),
.B2(n_3030),
.Y(n_3052)
);

AOI211xp5_ASAP7_75t_L g3053 ( 
.A1(n_3020),
.A2(n_1051),
.B(n_1015),
.C(n_1119),
.Y(n_3053)
);

NOR2x2_ASAP7_75t_L g3054 ( 
.A(n_3017),
.B(n_1080),
.Y(n_3054)
);

XOR2x2_ASAP7_75t_L g3055 ( 
.A(n_3010),
.B(n_1191),
.Y(n_3055)
);

XNOR2xp5_ASAP7_75t_L g3056 ( 
.A(n_3010),
.B(n_1048),
.Y(n_3056)
);

AOI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_3028),
.A2(n_1196),
.B1(n_1279),
.B2(n_1191),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_3038),
.A2(n_1211),
.B1(n_1271),
.B2(n_1279),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_3046),
.A2(n_1211),
.B1(n_1271),
.B2(n_1278),
.Y(n_3059)
);

AOI31xp33_ASAP7_75t_L g3060 ( 
.A1(n_3056),
.A2(n_1080),
.A3(n_1086),
.B(n_1019),
.Y(n_3060)
);

AOI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_3049),
.A2(n_1086),
.B1(n_1048),
.B2(n_1021),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_3055),
.A2(n_1021),
.B1(n_1015),
.B2(n_1134),
.Y(n_3062)
);

AOI22xp33_ASAP7_75t_L g3063 ( 
.A1(n_3034),
.A2(n_1021),
.B1(n_1015),
.B2(n_1134),
.Y(n_3063)
);

AOI31xp33_ASAP7_75t_L g3064 ( 
.A1(n_3041),
.A2(n_1237),
.A3(n_1210),
.B(n_1208),
.Y(n_3064)
);

AOI31xp33_ASAP7_75t_L g3065 ( 
.A1(n_3053),
.A2(n_1205),
.A3(n_1190),
.B(n_1184),
.Y(n_3065)
);

AOI31xp33_ASAP7_75t_L g3066 ( 
.A1(n_3047),
.A2(n_1205),
.A3(n_1190),
.B(n_1184),
.Y(n_3066)
);

AOI31xp33_ASAP7_75t_L g3067 ( 
.A1(n_3037),
.A2(n_1351),
.A3(n_1101),
.B(n_1135),
.Y(n_3067)
);

AOI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_3052),
.A2(n_1081),
.B1(n_1015),
.B2(n_1024),
.Y(n_3068)
);

AOI31xp33_ASAP7_75t_L g3069 ( 
.A1(n_3054),
.A2(n_1084),
.A3(n_1066),
.B(n_1040),
.Y(n_3069)
);

AOI31xp33_ASAP7_75t_L g3070 ( 
.A1(n_3036),
.A2(n_1084),
.A3(n_1066),
.B(n_1040),
.Y(n_3070)
);

AOI22xp33_ASAP7_75t_L g3071 ( 
.A1(n_3052),
.A2(n_1081),
.B1(n_1024),
.B2(n_1040),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_3040),
.A2(n_3050),
.B1(n_3043),
.B2(n_3035),
.Y(n_3072)
);

XNOR2xp5_ASAP7_75t_L g3073 ( 
.A(n_3072),
.B(n_3048),
.Y(n_3073)
);

AOI21x1_ASAP7_75t_L g3074 ( 
.A1(n_3069),
.A2(n_3042),
.B(n_3044),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_3062),
.Y(n_3075)
);

OAI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_3063),
.A2(n_3045),
.B(n_3057),
.Y(n_3076)
);

OAI22x1_ASAP7_75t_L g3077 ( 
.A1(n_3060),
.A2(n_3039),
.B1(n_3051),
.B2(n_1066),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_3070),
.A2(n_1119),
.B(n_1024),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_3068),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_3067),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_3065),
.Y(n_3081)
);

OAI21x1_ASAP7_75t_SL g3082 ( 
.A1(n_3071),
.A2(n_1119),
.B(n_1024),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_3066),
.A2(n_1119),
.B(n_1024),
.Y(n_3083)
);

CKINVDCx20_ASAP7_75t_R g3084 ( 
.A(n_3058),
.Y(n_3084)
);

INVx4_ASAP7_75t_L g3085 ( 
.A(n_3081),
.Y(n_3085)
);

AND2x4_ASAP7_75t_L g3086 ( 
.A(n_3076),
.B(n_3061),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_3073),
.A2(n_3064),
.B(n_3059),
.Y(n_3087)
);

NOR2xp67_ASAP7_75t_L g3088 ( 
.A(n_3077),
.B(n_1119),
.Y(n_3088)
);

OA21x2_ASAP7_75t_L g3089 ( 
.A1(n_3080),
.A2(n_3078),
.B(n_3079),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_3075),
.B(n_1119),
.Y(n_3090)
);

OAI21x1_ASAP7_75t_L g3091 ( 
.A1(n_3074),
.A2(n_1239),
.B(n_1024),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_3082),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_3087),
.A2(n_3083),
.B(n_3084),
.Y(n_3093)
);

NAND2xp33_ASAP7_75t_SL g3094 ( 
.A(n_3085),
.B(n_3090),
.Y(n_3094)
);

AO221x1_ASAP7_75t_L g3095 ( 
.A1(n_3092),
.A2(n_1134),
.B1(n_1040),
.B2(n_1045),
.C(n_1047),
.Y(n_3095)
);

OAI21x1_ASAP7_75t_SL g3096 ( 
.A1(n_3089),
.A2(n_1134),
.B(n_1040),
.Y(n_3096)
);

AOI21xp33_ASAP7_75t_SL g3097 ( 
.A1(n_3086),
.A2(n_1134),
.B(n_1040),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_3088),
.A2(n_3091),
.B(n_1045),
.Y(n_3098)
);

BUFx2_ASAP7_75t_L g3099 ( 
.A(n_3094),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3096),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_3099),
.A2(n_3093),
.B(n_3098),
.Y(n_3101)
);

AOI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_3101),
.A2(n_3100),
.B(n_3097),
.Y(n_3102)
);

AOI211xp5_ASAP7_75t_L g3103 ( 
.A1(n_3102),
.A2(n_3095),
.B(n_1045),
.C(n_1047),
.Y(n_3103)
);


endmodule