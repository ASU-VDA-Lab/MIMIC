module fake_jpeg_9012_n_92 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_2),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_3),
.C(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_13),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

XNOR2x1_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_20),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_15),
.C(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_11),
.C(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_24),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_24),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_15),
.B1(n_17),
.B2(n_13),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_51),
.B(n_54),
.Y(n_72)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_24),
.C(n_27),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_46),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_64),
.B1(n_51),
.B2(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_78),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_65),
.C(n_63),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_76),
.C(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_59),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_18),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_82),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_5),
.C(n_6),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_6),
.B(n_7),
.Y(n_88)
);

NOR2x1p5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_7),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_9),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_87),
.Y(n_92)
);


endmodule