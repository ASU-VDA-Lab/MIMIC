module real_jpeg_6784_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g89 ( 
.A(n_0),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_0),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_0),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_0),
.B(n_128),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_1),
.Y(n_293)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_2),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_2),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_2),
.B(n_258),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_2),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_3),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_3),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_4),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_4),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_4),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_4),
.B(n_443),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_7),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_7),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_8),
.Y(n_231)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_8),
.Y(n_245)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_8),
.Y(n_331)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_12),
.B(n_134),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_12),
.B(n_139),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_12),
.B(n_244),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_12),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_12),
.B(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_12),
.B(n_99),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_12),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_12),
.B(n_172),
.Y(n_483)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_14),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_14),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_14),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_14),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_15),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_15),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_15),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_15),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_15),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_15),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_225),
.Y(n_386)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_17),
.B(n_125),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_17),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_17),
.B(n_42),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_17),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_17),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_17),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_18),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_18),
.B(n_106),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_18),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_18),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_19),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_19),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_19),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_19),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_19),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_19),
.B(n_244),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_19),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_19),
.B(n_459),
.Y(n_458)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_117),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_116),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_75),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_75),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_58),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.C(n_41),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_41),
.B1(n_57),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_36),
.A2(n_62),
.B1(n_71),
.B2(n_107),
.Y(n_111)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_38),
.Y(n_258)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_40),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_44),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_44),
.Y(n_437)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_60),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_66),
.C(n_71),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_65),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_67),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_71),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_178)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_73),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_73),
.Y(n_347)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_74),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_112),
.C(n_113),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_76),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_101),
.C(n_108),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_77),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_93),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_97),
.C(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.C(n_88),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_88),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_89),
.B(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_101),
.A2(n_108),
.B1(n_109),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_105),
.B1(n_151),
.B2(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_104),
.B(n_147),
.C(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_112),
.B(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_186),
.B(n_525),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_184),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_119),
.B(n_184),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_176),
.C(n_181),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_120),
.B(n_511),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_156),
.C(n_158),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_121),
.B(n_514),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_137),
.C(n_146),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_122),
.B(n_137),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_131),
.C(n_136),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_125),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_129),
.Y(n_240)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_143),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_138),
.B(n_143),
.Y(n_474)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_142),
.B(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_146),
.B(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_161),
.C(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_151),
.A2(n_155),
.B1(n_161),
.B2(n_162),
.Y(n_470)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_154),
.Y(n_305)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_154),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_156),
.Y(n_515)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.C(n_173),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_160),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_161),
.A2(n_162),
.B1(n_454),
.B2(n_456),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_161),
.B(n_454),
.C(n_457),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_164),
.B(n_470),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_501)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_173),
.A2(n_174),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_174),
.B(n_484),
.C(n_499),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_176),
.B(n_181),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_180),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_177),
.B(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_179),
.B(n_180),
.Y(n_517)
);

AO21x1_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_506),
.B(n_522),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_489),
.B(n_505),
.Y(n_187)
);

AOI21x1_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_463),
.B(n_488),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_420),
.B(n_462),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_379),
.B(n_419),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_298),
.B(n_378),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_283),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_193),
.B(n_283),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_234),
.B2(n_282),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_194),
.B(n_235),
.C(n_266),
.Y(n_418)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_211),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_196),
.B(n_212),
.C(n_233),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.C(n_210),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_197),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_288)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_207),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_208),
.B(n_210),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_221),
.B1(n_232),
.B2(n_233),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_216),
.B(n_220),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_216),
.Y(n_220)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_220),
.B(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_220),
.B(n_384),
.C(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_222),
.B(n_227),
.C(n_230),
.Y(n_417)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_266),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_247),
.C(n_259),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_241),
.C(n_246),
.Y(n_281)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_245),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_248),
.B1(n_259),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.C(n_256),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_249),
.A2(n_250),
.B1(n_256),
.B2(n_257),
.Y(n_371)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_251),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_254),
.Y(n_406)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_264),
.Y(n_280)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

BUFx8_ASAP7_75t_L g455 ( 
.A(n_263),
.Y(n_455)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

XOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_279),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_267),
.B(n_280),
.C(n_281),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_268),
.B(n_273),
.C(n_277),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_273),
.B1(n_277),
.B2(n_278),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_272),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_273),
.Y(n_278)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_276),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.C(n_296),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_284),
.B(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_287),
.B(n_296),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_289),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_294),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_373),
.B(n_377),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_358),
.B(n_372),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_338),
.B(n_357),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_325),
.B(n_337),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_309),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_319),
.B2(n_320),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_316),
.C(n_319),
.Y(n_356)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_315),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_324),
.Y(n_342)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_332),
.B(n_336),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_328),
.Y(n_336)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_356),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_342),
.C(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_353),
.C(n_355),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx11_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_349),
.Y(n_355)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_361),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_368),
.C(n_369),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_375),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_418),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_418),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_399),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_383),
.C(n_399),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_396),
.B2(n_398),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_389),
.C(n_391),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_391),
.B2(n_392),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_396),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_402),
.C(n_412),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_412),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_408),
.C(n_409),
.Y(n_450)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_417),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_416),
.C(n_417),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_422),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_440),
.C(n_460),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_440),
.B1(n_460),
.B2(n_461),
.Y(n_424)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_428),
.B2(n_439),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_429),
.C(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_438),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_435),
.C(n_438),
.Y(n_480)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx6_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_449),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_450),
.C(n_451),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_441),
.Y(n_528)
);

FAx1_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_445),
.CI(n_448),
.CON(n_441),
.SN(n_441)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_442),
.B(n_445),
.C(n_448),
.Y(n_485)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_457),
.B2(n_458),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_454),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_487),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_487),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_467),
.C(n_476),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_476),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_475),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_472),
.C(n_473),
.Y(n_495)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_471),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_478),
.B1(n_479),
.B2(n_486),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_480),
.C(n_481),
.Y(n_491)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_479),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.Y(n_481)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_483),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_504),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_504),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_493),
.C(n_502),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_502),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_498),
.C(n_500),
.Y(n_518)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_519),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_509),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_512),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_512),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.C(n_518),
.Y(n_512)
);

FAx1_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_516),
.CI(n_518),
.CON(n_520),
.SN(n_520)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_521),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_520),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);


endmodule