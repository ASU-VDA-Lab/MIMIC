module real_jpeg_26553_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_37),
.B1(n_38),
.B2(n_60),
.Y(n_91)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_19),
.B1(n_44),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_19),
.B1(n_37),
.B2(n_38),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_25),
.B(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_135),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_6),
.B(n_38),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_58),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_5),
.A2(n_8),
.B(n_28),
.C(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_10),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_99),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_97),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_79),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_79),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_14),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_61),
.CI(n_66),
.CON(n_14),
.SN(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_16),
.A2(n_17),
.B1(n_69),
.B2(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_16),
.A2(n_17),
.B1(n_64),
.B2(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_16),
.A2(n_17),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_17),
.A2(n_67),
.B(n_78),
.Y(n_66)
);

AOI211xp5_ASAP7_75t_L g106 ( 
.A1(n_17),
.A2(n_94),
.B(n_96),
.C(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_19),
.A2(n_20),
.B(n_26),
.C(n_121),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_19),
.A2(n_40),
.B(n_45),
.C(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_19),
.B(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_19),
.B(n_157),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_19),
.A2(n_44),
.B(n_56),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_27),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_28),
.A2(n_29),
.B1(n_54),
.B2(n_56),
.Y(n_57)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_46),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_35),
.B(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_41),
.B1(n_46),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_41),
.B1(n_63),
.B2(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_37),
.B(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_72),
.Y(n_73)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_45),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_62),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_64),
.A2(n_88),
.B1(n_94),
.B2(n_108),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_122),
.C(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_64),
.A2(n_88),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_69),
.A2(n_75),
.B1(n_78),
.B2(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_73),
.B1(n_91),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_74),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_75),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_84),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_80),
.B(n_83),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_84),
.A2(n_85),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B(n_95),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_86),
.A2(n_95),
.B(n_197),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_87),
.A2(n_96),
.B(n_124),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_108),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_88),
.A2(n_108),
.B(n_169),
.C(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_89),
.A2(n_116),
.B1(n_117),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_89),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_90),
.A2(n_94),
.B1(n_108),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_90),
.Y(n_200)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_108),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_108),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_94),
.A2(n_108),
.B1(n_143),
.B2(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_122),
.C(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_94),
.A2(n_108),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_94),
.B(n_175),
.C(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_94),
.B(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_215),
.B(n_220),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_205),
.B(n_214),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_136),
.B(n_192),
.C(n_204),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_125),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_103),
.B(n_125),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_105),
.B(n_110),
.C(n_115),
.Y(n_193)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_111),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_124),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_116),
.A2(n_117),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_123),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_123),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_123),
.B1(n_133),
.B2(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.C(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_126),
.A2(n_127),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_129),
.B1(n_165),
.B2(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_191),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_184),
.B(n_190),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_171),
.B(n_183),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_162),
.B(n_170),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_150),
.B(n_161),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_174),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_194),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_197),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.C(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);


endmodule