module fake_jpeg_22247_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_29)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx12_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_12),
.B1(n_10),
.B2(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_23),
.B1(n_25),
.B2(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_31),
.B1(n_34),
.B2(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_38),
.B1(n_35),
.B2(n_43),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_36),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_11),
.C(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_23),
.B1(n_25),
.B2(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_56),
.B1(n_42),
.B2(n_38),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_23),
.B1(n_12),
.B2(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_66),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_60),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_62),
.B(n_65),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_35),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_45),
.B(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_43),
.C(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_52),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_76),
.C(n_64),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_54),
.B(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_81),
.C(n_13),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_58),
.C(n_65),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_84),
.C(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_63),
.C(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_73),
.B1(n_76),
.B2(n_57),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_90),
.C(n_21),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_67),
.B1(n_56),
.B2(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_21),
.C(n_19),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.C(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_94),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_97),
.B(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_35),
.B1(n_11),
.B2(n_9),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_4),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_4),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_103),
.B(n_6),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_100),
.C2(n_58),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_5),
.B(n_6),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_7),
.Y(n_108)
);


endmodule