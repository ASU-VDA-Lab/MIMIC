module fake_jpeg_26555_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_17),
.B1(n_23),
.B2(n_16),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_60),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_20),
.B1(n_27),
.B2(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_69),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_96),
.B1(n_98),
.B2(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_35),
.B1(n_43),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_84),
.B1(n_40),
.B2(n_27),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_37),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_26),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_36),
.B1(n_39),
.B2(n_34),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_95),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_93),
.B1(n_29),
.B2(n_19),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_41),
.C(n_43),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_41),
.C(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_21),
.B1(n_29),
.B2(n_18),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_102),
.B1(n_19),
.B2(n_33),
.Y(n_123)
);

AOI22x1_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_127),
.B1(n_129),
.B2(n_69),
.Y(n_139)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_107),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_36),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_116),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_70),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_41),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_110),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_126),
.B1(n_91),
.B2(n_103),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_41),
.C(n_34),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_88),
.C(n_98),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_77),
.C(n_85),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_71),
.A2(n_40),
.B1(n_26),
.B2(n_41),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_41),
.B1(n_34),
.B2(n_36),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_136),
.B(n_146),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_102),
.B(n_80),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_161),
.B1(n_164),
.B2(n_39),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_156),
.B1(n_158),
.B2(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_150),
.C(n_162),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_120),
.B(n_127),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_115),
.B(n_31),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_157),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_128),
.B(n_116),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_154),
.A3(n_160),
.B1(n_132),
.B2(n_28),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_95),
.C(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_67),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_109),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_68),
.B1(n_105),
.B2(n_75),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_106),
.A2(n_85),
.B(n_84),
.C(n_28),
.D(n_97),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_87),
.B1(n_99),
.B2(n_101),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_101),
.C(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_85),
.B1(n_96),
.B2(n_94),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_73),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_25),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_135),
.B1(n_115),
.B2(n_27),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_36),
.C(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_187),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_132),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_186),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_182),
.B(n_188),
.Y(n_213)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_32),
.A3(n_31),
.B1(n_19),
.B2(n_117),
.Y(n_176)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_184),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_138),
.B(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_134),
.B1(n_111),
.B2(n_66),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_144),
.B1(n_150),
.B2(n_143),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_189),
.C(n_3),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_111),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_1),
.B(n_2),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_34),
.C(n_39),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_200),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_25),
.B1(n_22),
.B2(n_15),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_215),
.B(n_198),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_211),
.B1(n_220),
.B2(n_222),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_141),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_210),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_167),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_25),
.B1(n_22),
.B2(n_15),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_25),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_173),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_190),
.B1(n_195),
.B2(n_172),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_22),
.B1(n_12),
.B2(n_11),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_182),
.A2(n_3),
.B(n_4),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_223),
.A2(n_228),
.B(n_176),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_3),
.C(n_5),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_181),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_174),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_3),
.B(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_178),
.B(n_198),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_233),
.B(n_238),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_244),
.B(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_246),
.B1(n_218),
.B2(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_173),
.B1(n_191),
.B2(n_185),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_192),
.B1(n_171),
.B2(n_197),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_247),
.A2(n_204),
.B1(n_224),
.B2(n_201),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_8),
.B(n_11),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_8),
.C(n_11),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_206),
.B(n_8),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_204),
.B1(n_203),
.B2(n_221),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_262),
.B1(n_270),
.B2(n_239),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_203),
.B(n_205),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_246),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_247),
.B1(n_239),
.B2(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_232),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_219),
.B1(n_207),
.B2(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_236),
.C(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_285),
.C(n_261),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_240),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_240),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_210),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_250),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_229),
.B1(n_207),
.B2(n_244),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_286),
.B(n_223),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_233),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_212),
.C(n_251),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_208),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_297),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_256),
.C(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_263),
.C(n_229),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_283),
.Y(n_295)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_235),
.CI(n_285),
.CON(n_298),
.SN(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_293),
.B(n_287),
.C(n_297),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_261),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_276),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_282),
.B1(n_278),
.B2(n_254),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_292),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_253),
.C(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_308),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_298),
.B1(n_302),
.B2(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_273),
.C(n_248),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_314),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_281),
.B1(n_269),
.B2(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_313),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_315),
.C(n_318),
.Y(n_321)
);

AO221x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_319),
.B1(n_310),
.B2(n_307),
.C(n_298),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_228),
.B(n_292),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_215),
.B(n_10),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_10),
.C(n_12),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_5),
.Y(n_326)
);


endmodule