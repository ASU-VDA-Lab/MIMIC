module fake_aes_11130_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
NAND2xp33_ASAP7_75t_L g15 ( .A(n_5), .B(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_4), .B(n_1), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
AOI22xp5_ASAP7_75t_SL g18 ( .A1(n_11), .A2(n_17), .B1(n_13), .B2(n_14), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_14), .B(n_2), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_15), .B(n_12), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI221xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_18), .B1(n_20), .B2(n_19), .C(n_6), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_20), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_27), .B(n_20), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_26), .B(n_24), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_29), .B(n_20), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g31 ( .A(n_28), .B(n_26), .Y(n_31) );
OAI22xp5_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_19), .B1(n_8), .B2(n_9), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OR3x2_ASAP7_75t_L g35 ( .A(n_34), .B(n_33), .C(n_19), .Y(n_35) );
endmodule