module fake_netlist_5_1663_n_3794 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_785, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_802, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_753, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_788, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_755, n_6, n_509, n_568, n_39, n_147, n_373, n_757, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_375, n_301, n_779, n_576, n_68, n_804, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_741, n_548, n_543, n_260, n_812, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_752, n_331, n_10, n_24, n_406, n_519, n_470, n_782, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_760, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_798, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_813, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_144, n_114, n_96, n_772, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_236, n_388, n_761, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_770, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_745, n_627, n_767, n_172, n_206, n_217, n_440, n_726, n_478, n_793, n_545, n_441, n_450, n_648, n_312, n_476, n_818, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_805, n_117, n_326, n_794, n_768, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_815, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_159, n_334, n_599, n_766, n_811, n_541, n_807, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_803, n_238, n_639, n_799, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_817, n_360, n_36, n_594, n_764, n_200, n_162, n_64, n_759, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_324, n_810, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_747, n_52, n_278, n_784, n_110, n_3794);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_755;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_757;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_375;
input n_301;
input n_779;
input n_576;
input n_68;
input n_804;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_782;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_813;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_144;
input n_114;
input n_96;
input n_772;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_761;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_805;
input n_117;
input n_326;
input n_794;
input n_768;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_238;
input n_639;
input n_799;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_817;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_162;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3794;

wire n_924;
wire n_1263;
wire n_3304;
wire n_2253;
wire n_2417;
wire n_1378;
wire n_977;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_2380;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_2899;
wire n_2955;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_880;
wire n_3086;
wire n_3297;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_2347;
wire n_1292;
wire n_2520;
wire n_2821;
wire n_1370;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_3641;
wire n_956;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_2487;
wire n_1695;
wire n_1466;
wire n_3766;
wire n_1353;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_854;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1462;
wire n_3621;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_1107;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_2963;
wire n_1098;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_2888;
wire n_1483;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1633;
wire n_1236;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_3631;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_976;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_3490;
wire n_3656;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_2099;
wire n_2408;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1749;
wire n_1036;
wire n_1097;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_897;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3702;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_2439;
wire n_1931;
wire n_1218;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_3744;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_2615;
wire n_1556;
wire n_1384;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1986;
wire n_1471;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3716;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_2713;
wire n_3544;
wire n_2700;
wire n_2644;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_3096;
wire n_2251;
wire n_1447;
wire n_1377;
wire n_2370;
wire n_3496;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_2248;
wire n_2356;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_2622;
wire n_1278;
wire n_2062;
wire n_2668;
wire n_3714;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_1058;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_3781;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_884;
wire n_3328;
wire n_944;
wire n_1754;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_3433;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_832;
wire n_857;
wire n_2305;
wire n_3430;
wire n_3392;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_2837;
wire n_847;
wire n_2319;
wire n_1393;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_3655;
wire n_2808;
wire n_3009;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_3640;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1847;
wire n_1199;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_1711;
wire n_931;
wire n_870;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_3790;
wire n_3491;
wire n_935;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_3643;
wire n_2222;
wire n_1892;
wire n_3510;
wire n_3745;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_2690;
wire n_1189;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1925;
wire n_1194;
wire n_3660;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_3775;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_2629;
wire n_1415;
wire n_2592;
wire n_3416;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_3770;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_3469;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_946;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_3113;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_3760;
wire n_1760;
wire n_2875;
wire n_936;
wire n_2960;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_3030;
wire n_1068;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_906;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_3031;
wire n_3396;
wire n_3701;
wire n_940;
wire n_1445;
wire n_3516;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_2507;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2320;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2093;
wire n_2473;
wire n_1079;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3741;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_2536;
wire n_1592;
wire n_1065;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_974;
wire n_1159;
wire n_957;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_2897;
wire n_2077;
wire n_1416;
wire n_3614;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_3411;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2879;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_860;
wire n_3229;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_3788;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_3421;
wire n_2240;
wire n_2696;
wire n_1351;
wire n_1205;
wire n_2436;
wire n_1044;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_1684;
wire n_996;
wire n_921;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_1840;
wire n_1082;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_2969;
wire n_2191;
wire n_2864;
wire n_1311;
wire n_3195;
wire n_1519;
wire n_950;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_912;
wire n_968;
wire n_3548;
wire n_2440;
wire n_1699;
wire n_1386;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_841;
wire n_1050;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1644;
wire n_1283;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_1203;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_2993;
wire n_1719;
wire n_1048;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_2499;
wire n_1200;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1668;
wire n_1363;
wire n_3737;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_828;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3572;
wire n_992;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_842;
wire n_3734;
wire n_984;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_3400;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_918;
wire n_3529;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1977;
wire n_1557;
wire n_2153;
wire n_1147;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_3196;
wire n_1422;
wire n_3078;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1511;
wire n_1470;
wire n_2094;
wire n_1096;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2393;
wire n_833;
wire n_2318;
wire n_3689;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_988;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_2751;
wire n_2707;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_2311;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_2285;
wire n_1446;
wire n_3147;
wire n_2758;
wire n_2471;
wire n_1472;
wire n_2298;
wire n_1176;
wire n_1458;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3708;
wire n_1204;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_3636;
wire n_2588;
wire n_2962;
wire n_1188;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_849;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3380;
wire n_3177;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_3393;
wire n_1603;
wire n_1232;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_3520;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_3192;
wire n_2608;
wire n_3764;
wire n_2657;
wire n_2995;
wire n_2494;
wire n_1375;
wire n_3547;
wire n_2649;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1929;
wire n_1392;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_2409;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_1253;
wire n_3408;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1514;
wire n_1777;
wire n_1335;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_2605;
wire n_1310;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_3308;
wire n_2665;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_3757;
wire n_3438;
wire n_872;
wire n_2012;
wire n_3792;
wire n_1291;
wire n_3381;
wire n_3503;
wire n_1753;
wire n_1297;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_2184;
wire n_1184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_827;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_2926;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_1137;
wire n_3046;
wire n_2213;
wire n_1170;
wire n_2023;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_823;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1817;
wire n_1944;
wire n_909;
wire n_1683;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3070;
wire n_3284;
wire n_1326;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_825;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_3700;
wire n_3609;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_1867;
wire n_1330;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2774;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_3391;
wire n_1567;
wire n_2567;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_839;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_2173;
wire n_1250;
wire n_3722;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_928;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_2030;
wire n_1348;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_2797;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_1028;
wire n_3336;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3114;
wire n_2594;
wire n_3125;
wire n_3234;
wire n_2394;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3591;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_3247;
wire n_1604;
wire n_2525;
wire n_2513;
wire n_1275;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_2225;
wire n_3613;
wire n_3567;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_1558;
wire n_1340;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_835;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_927;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_1004;
wire n_1186;
wire n_2614;
wire n_1032;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_2599;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_2524;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_3159;
wire n_2728;
wire n_2268;
wire n_3778;

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_524),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_559),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_464),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_594),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_554),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_701),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_12),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_481),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_496),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_529),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_784),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_390),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_14),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_507),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_138),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_475),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_485),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_375),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_71),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_271),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_718),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_181),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_229),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_493),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_581),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_609),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_742),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_105),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_334),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_708),
.Y(n_849)
);

CKINVDCx16_ASAP7_75t_R g850 ( 
.A(n_651),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_598),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_530),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_547),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_26),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_356),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_457),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_124),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_555),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_23),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_686),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_53),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_515),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_612),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_474),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_534),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_589),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_370),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_233),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_679),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_660),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_355),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_676),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_811),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_501),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_783),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_476),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_37),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_618),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_556),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_173),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_641),
.Y(n_882)
);

BUFx5_ASAP7_75t_L g883 ( 
.A(n_702),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_219),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_758),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_118),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_804),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_693),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_170),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_623),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_665),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_730),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_188),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_95),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_418),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_436),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_155),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_763),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_535),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_194),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_569),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_436),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_371),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_69),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_513),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_640),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_320),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_694),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_724),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_30),
.Y(n_910)
);

BUFx5_ASAP7_75t_L g911 ( 
.A(n_361),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_661),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_675),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_486),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_487),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_495),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_353),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_585),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_463),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_301),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_613),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_517),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_786),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_635),
.Y(n_924)
);

BUFx2_ASAP7_75t_SL g925 ( 
.A(n_326),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_169),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_403),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_780),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_165),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_256),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_684),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_752),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_750),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_697),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_740),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_721),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_582),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_733),
.Y(n_938)
);

BUFx10_ASAP7_75t_L g939 ( 
.A(n_372),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_816),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_801),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_389),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_765),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_89),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_197),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_266),
.Y(n_946)
);

CKINVDCx16_ASAP7_75t_R g947 ( 
.A(n_269),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_653),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_217),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_272),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_545),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_448),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_734),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_513),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_17),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_507),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_219),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_192),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_712),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_131),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_122),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_813),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_130),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_435),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_746),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_792),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_467),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_789),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_638),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_61),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_103),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_142),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_257),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_261),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_546),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_283),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_254),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_349),
.Y(n_978)
);

CKINVDCx16_ASAP7_75t_R g979 ( 
.A(n_456),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_551),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_53),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_245),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_500),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_604),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_518),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_417),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_288),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_146),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_154),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_814),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_189),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_768),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_295),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_626),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_326),
.Y(n_995)
);

INVxp67_ASAP7_75t_SL g996 ( 
.A(n_722),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_386),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_46),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_649),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_297),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_258),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_755),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_504),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_809),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_206),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_126),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_471),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_771),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_647),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_682),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_406),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_472),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_180),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_692),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_776),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_600),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_244),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_528),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_720),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_790),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_802),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_338),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_362),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_732),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_691),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_68),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_193),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_248),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_671),
.Y(n_1029)
);

BUFx8_ASAP7_75t_SL g1030 ( 
.A(n_634),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_631),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_302),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_621),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_406),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_529),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_544),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_685),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_605),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_185),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_118),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_411),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_312),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_266),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_140),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_51),
.Y(n_1045)
);

CKINVDCx16_ASAP7_75t_R g1046 ( 
.A(n_711),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_230),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_142),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_360),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_505),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_85),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_492),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_344),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_240),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_249),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_132),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_796),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_179),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_482),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_442),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_40),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_8),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_580),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_710),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_293),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_11),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_429),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_350),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_462),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_532),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_473),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_300),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_762),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_666),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_390),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_428),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_40),
.Y(n_1077)
);

BUFx10_ASAP7_75t_L g1078 ( 
.A(n_125),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_189),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_549),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_32),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_119),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_99),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_362),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_591),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_431),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_367),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_566),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_497),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_565),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_808),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_514),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_175),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_775),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_429),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_739),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_163),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_214),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_560),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_663),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_484),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_491),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_778),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_664),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_508),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_331),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_134),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_375),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_644),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_267),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_599),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_650),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_633),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_494),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_736),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_59),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_648),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_403),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_163),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_143),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_550),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_476),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_200),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_539),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_688),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_616),
.Y(n_1126)
);

BUFx5_ASAP7_75t_L g1127 ( 
.A(n_656),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_532),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_639),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_807),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_596),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_731),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_158),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_98),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_818),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_286),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_90),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_495),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_231),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_333),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_58),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_254),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_646),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_144),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_696),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_788),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_198),
.Y(n_1147)
);

BUFx10_ASAP7_75t_L g1148 ( 
.A(n_608),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_218),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_446),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_748),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_322),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_11),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_363),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_719),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_713),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_799),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_430),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_628),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_133),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_29),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_329),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_237),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_537),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_310),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_667),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_277),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_497),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_23),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_615),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_817),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_173),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_506),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_251),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_204),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_330),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_700),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_361),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_678),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_203),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_520),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_695),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_738),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_153),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_680),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_548),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_745),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_510),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_271),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_761),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_220),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_759),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_256),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_527),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_417),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_259),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_224),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_145),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_709),
.Y(n_1199)
);

BUFx5_ASAP7_75t_L g1200 ( 
.A(n_593),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_66),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_157),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_194),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_726),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_629),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_418),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_463),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_531),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_757),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_442),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_488),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_772),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_381),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_652),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_22),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_774),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_520),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_499),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_595),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_112),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_543),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_462),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_578),
.Y(n_1223)
);

BUFx5_ASAP7_75t_L g1224 ( 
.A(n_766),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_503),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_617),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_320),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_249),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_183),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_563),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_528),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_293),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_376),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_373),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_575),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_502),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_433),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_448),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_735),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_769),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_669),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_672),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_819),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_553),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_627),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_466),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_662),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_681),
.Y(n_1248)
);

BUFx10_ASAP7_75t_L g1249 ( 
.A(n_716),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_114),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_453),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_557),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_453),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_420),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_150),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_199),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_80),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_198),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_568),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_630),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_572),
.Y(n_1261)
);

CKINVDCx12_ASAP7_75t_R g1262 ( 
.A(n_98),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_798),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_527),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_525),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_276),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_642),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_655),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_279),
.Y(n_1269)
);

INVxp33_ASAP7_75t_L g1270 ( 
.A(n_96),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_521),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_445),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_574),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_365),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_597),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_365),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_756),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_728),
.Y(n_1278)
);

BUFx10_ASAP7_75t_L g1279 ( 
.A(n_420),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_135),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_455),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_319),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_744),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_413),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_499),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_491),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_425),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_60),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_637),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_619),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_767),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_760),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_221),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_39),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_622),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_360),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_567),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_538),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_571),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_717),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_795),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_246),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_704),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_6),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_232),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_213),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_606),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_741),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_533),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_358),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_441),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_312),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_601),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_247),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_625),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_677),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_570),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_690),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_564),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_501),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_614),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_673),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_274),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_522),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_200),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_725),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_446),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_534),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_175),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_437),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_3),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_208),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_577),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_586),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_715),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_643),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_803),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_636),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_815),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_607),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_787),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_192),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_689),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_558),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_52),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_810),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_97),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_348),
.Y(n_1349)
);

CKINVDCx14_ASAP7_75t_R g1350 ( 
.A(n_498),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_723),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_227),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_9),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_141),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_505),
.Y(n_1355)
);

CKINVDCx14_ASAP7_75t_R g1356 ( 
.A(n_151),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_542),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_285),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_632),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_533),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_473),
.Y(n_1361)
);

CKINVDCx14_ASAP7_75t_R g1362 ( 
.A(n_182),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_157),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_674),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_79),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_93),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_373),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_523),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_773),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_516),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_645),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_228),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_84),
.Y(n_1373)
);

BUFx5_ASAP7_75t_L g1374 ( 
.A(n_791),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_525),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_521),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_576),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_93),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_358),
.Y(n_1379)
);

CKINVDCx14_ASAP7_75t_R g1380 ( 
.A(n_61),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_754),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_785),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_714),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_751),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_253),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_812),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_592),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_610),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_602),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_354),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_654),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_583),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_137),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_35),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_327),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_279),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_526),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_82),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_541),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_223),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_176),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_518),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_437),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_806),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_319),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_166),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_603),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_380),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_611),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_377),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_454),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_579),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_698),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_260),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_737),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_770),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_506),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_330),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_729),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_540),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_588),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_805),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_657),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_100),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_269),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_183),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_19),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_398),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_280),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_286),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_341),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_561),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_519),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_797),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_743),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_624),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_699),
.Y(n_1437)
);

CKINVDCx16_ASAP7_75t_R g1438 ( 
.A(n_388),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_466),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_706),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_703),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_125),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_327),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_388),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_323),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_573),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_781),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_24),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_509),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_687),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_504),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_291),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_227),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_707),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_584),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_338),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_324),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_590),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_150),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_512),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_562),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_705),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_237),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_794),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_210),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_469),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_317),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_511),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_782),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_793),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_409),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_196),
.Y(n_1472)
);

BUFx10_ASAP7_75t_L g1473 ( 
.A(n_668),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_407),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_683),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_620),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_434),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_281),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_727),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_777),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_275),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_222),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_478),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_658),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_96),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_470),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_779),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_308),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_490),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_483),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_158),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_587),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_489),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_276),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_749),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_281),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_4),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_670),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_477),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_88),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_247),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_800),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_764),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_224),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_469),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_480),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_202),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_753),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_425),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_39),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_479),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_747),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_552),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_866),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1030),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_926),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_866),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_866),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_866),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_866),
.Y(n_1520)
);

INVxp33_ASAP7_75t_SL g1521 ( 
.A(n_926),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_845),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_866),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_911),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1148),
.Y(n_1525)
);

CKINVDCx16_ASAP7_75t_R g1526 ( 
.A(n_826),
.Y(n_1526)
);

BUFx5_ASAP7_75t_L g1527 ( 
.A(n_823),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_911),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1503),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_911),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_911),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_821),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1428),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_859),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_911),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1428),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_986),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1262),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1145),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_828),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_941),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_986),
.Y(n_1542)
);

INVxp67_ASAP7_75t_SL g1543 ( 
.A(n_1145),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1011),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_820),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_830),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1431),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1391),
.B(n_1),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1011),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1391),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1013),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1013),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_840),
.Y(n_1553)
);

CKINVDCx16_ASAP7_75t_R g1554 ( 
.A(n_947),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1075),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1105),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1105),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_844),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1140),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_846),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1140),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1141),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1141),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1258),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1258),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1264),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_849),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_820),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1264),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1333),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_820),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1349),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_960),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1349),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1398),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1398),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1408),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1453),
.Y(n_1578)
);

INVxp33_ASAP7_75t_L g1579 ( 
.A(n_963),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_853),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1453),
.Y(n_1581)
);

INVxp33_ASAP7_75t_SL g1582 ( 
.A(n_1213),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1504),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1504),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_894),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_864),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1414),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1414),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_867),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_894),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_894),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_903),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_874),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_903),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_903),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_871),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_913),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_919),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_919),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_873),
.Y(n_1600)
);

INVxp33_ASAP7_75t_L g1601 ( 
.A(n_1321),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_979),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1026),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1438),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1026),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1355),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1026),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1089),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1089),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1089),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_876),
.Y(n_1611)
);

INVxp33_ASAP7_75t_L g1612 ( 
.A(n_1390),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1089),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_913),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_932),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1172),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1172),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1172),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1172),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_879),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1180),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1180),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1180),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1457),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1457),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1457),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_932),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1457),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_882),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_888),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1505),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1507),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_822),
.Y(n_1633)
);

BUFx10_ASAP7_75t_L g1634 ( 
.A(n_827),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1270),
.Y(n_1635)
);

CKINVDCx16_ASAP7_75t_R g1636 ( 
.A(n_1488),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_829),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_891),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_833),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_892),
.Y(n_1640)
);

INVxp33_ASAP7_75t_SL g1641 ( 
.A(n_831),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_836),
.Y(n_1642)
);

CKINVDCx16_ASAP7_75t_R g1643 ( 
.A(n_850),
.Y(n_1643)
);

CKINVDCx16_ASAP7_75t_R g1644 ( 
.A(n_1046),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1499),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_835),
.Y(n_1646)
);

INVxp33_ASAP7_75t_SL g1647 ( 
.A(n_832),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_899),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_883),
.Y(n_1649)
);

BUFx2_ASAP7_75t_SL g1650 ( 
.A(n_923),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_839),
.Y(n_1651)
);

INVxp33_ASAP7_75t_SL g1652 ( 
.A(n_834),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_852),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_883),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_965),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_857),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_865),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_933),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_856),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_856),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_897),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_883),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_902),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_883),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_939),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_920),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1024),
.B(n_0),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_956),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_957),
.Y(n_1669)
);

INVxp33_ASAP7_75t_SL g1670 ( 
.A(n_841),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_961),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1509),
.Y(n_1672)
);

CKINVDCx16_ASAP7_75t_R g1673 ( 
.A(n_1299),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_981),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_991),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_883),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_949),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1148),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_995),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_909),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_997),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_998),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1545),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1568),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1571),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1525),
.B(n_1678),
.Y(n_1686)
);

INVx5_ASAP7_75t_L g1687 ( 
.A(n_1646),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1568),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1585),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1602),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1622),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1624),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1626),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1628),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1590),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1546),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1591),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1604),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1592),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1553),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1539),
.B(n_933),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1558),
.B(n_1029),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1521),
.A2(n_1356),
.B1(n_1362),
.B2(n_1350),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1594),
.Y(n_1704)
);

AND2x2_ASAP7_75t_SL g1705 ( 
.A(n_1643),
.B(n_1364),
.Y(n_1705)
);

BUFx8_ASAP7_75t_L g1706 ( 
.A(n_1516),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1595),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1667),
.B(n_1024),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1537),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1543),
.B(n_1025),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1541),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1598),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1599),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1582),
.A2(n_838),
.B1(n_945),
.B2(n_942),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1603),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1541),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1526),
.A2(n_967),
.B1(n_993),
.B2(n_958),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1560),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1605),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1607),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1608),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1541),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1550),
.B(n_1025),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1567),
.B(n_1104),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1609),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1540),
.A2(n_1573),
.B1(n_1673),
.B2(n_1644),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1610),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1613),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1554),
.A2(n_1636),
.B1(n_1548),
.B2(n_1606),
.Y(n_1729)
);

BUFx12f_ASAP7_75t_L g1730 ( 
.A(n_1515),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1616),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1617),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1618),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1672),
.Y(n_1734)
);

AND2x6_ASAP7_75t_L g1735 ( 
.A(n_1542),
.B(n_1063),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1659),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1634),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1580),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1619),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1597),
.B(n_1063),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1621),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1623),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1625),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1517),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1518),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1544),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1549),
.Y(n_1747)
);

CKINVDCx11_ASAP7_75t_R g1748 ( 
.A(n_1522),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1551),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1570),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1528),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1514),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1586),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1589),
.Y(n_1754)
);

OA21x2_ASAP7_75t_L g1755 ( 
.A1(n_1519),
.A2(n_931),
.B(n_825),
.Y(n_1755)
);

OA21x2_ASAP7_75t_L g1756 ( 
.A1(n_1520),
.A2(n_851),
.B(n_824),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1631),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1587),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1523),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1614),
.B(n_1261),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1615),
.B(n_1268),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1588),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1660),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1579),
.A2(n_1022),
.B1(n_1061),
.B2(n_1043),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1632),
.Y(n_1765)
);

AOI22x1_ASAP7_75t_SL g1766 ( 
.A1(n_1529),
.A2(n_1067),
.B1(n_1069),
.B2(n_1066),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1633),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1538),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1637),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1639),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1524),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1627),
.B(n_1268),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1534),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1601),
.A2(n_1356),
.B1(n_1380),
.B2(n_1362),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1530),
.Y(n_1775)
);

INVx6_ASAP7_75t_L g1776 ( 
.A(n_1527),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1531),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1642),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1535),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1645),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1527),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1527),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1596),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1651),
.Y(n_1784)
);

CKINVDCx8_ASAP7_75t_R g1785 ( 
.A(n_1650),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1653),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1656),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1657),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1658),
.B(n_1261),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1661),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1533),
.B(n_1536),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1612),
.A2(n_1380),
.B1(n_1652),
.B2(n_1647),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1600),
.B(n_1611),
.Y(n_1793)
);

AND2x2_ASAP7_75t_SL g1794 ( 
.A(n_1547),
.B(n_1190),
.Y(n_1794)
);

AND2x2_ASAP7_75t_SL g1795 ( 
.A(n_1552),
.B(n_1190),
.Y(n_1795)
);

OA21x2_ASAP7_75t_L g1796 ( 
.A1(n_1649),
.A2(n_861),
.B(n_854),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1663),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1620),
.B(n_1273),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1629),
.B(n_1296),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1666),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1593),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1630),
.B(n_1334),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1668),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1555),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1669),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1671),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1674),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1640),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1556),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1557),
.Y(n_1810)
);

BUFx12f_ASAP7_75t_L g1811 ( 
.A(n_1648),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1680),
.B(n_1273),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1559),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1670),
.B(n_1292),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1675),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1679),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1561),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1527),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1681),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1638),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1682),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1562),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1563),
.B(n_1290),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1665),
.Y(n_1824)
);

AOI22x1_ASAP7_75t_SL g1825 ( 
.A1(n_1655),
.A2(n_1102),
.B1(n_1133),
.B2(n_1076),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1654),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1564),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1662),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1677),
.A2(n_1292),
.B1(n_1289),
.B2(n_1232),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1565),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1664),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1676),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1566),
.B(n_1290),
.Y(n_1833)
);

AOI22x1_ASAP7_75t_SL g1834 ( 
.A1(n_1569),
.A2(n_1217),
.B1(n_1237),
.B2(n_1202),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1572),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1574),
.B(n_1249),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1575),
.A2(n_1331),
.B1(n_1346),
.B2(n_1294),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1576),
.Y(n_1838)
);

CKINVDCx8_ASAP7_75t_R g1839 ( 
.A(n_1577),
.Y(n_1839)
);

CKINVDCx14_ASAP7_75t_R g1840 ( 
.A(n_1578),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1584),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1581),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1583),
.Y(n_1843)
);

INVx6_ASAP7_75t_L g1844 ( 
.A(n_1634),
.Y(n_1844)
);

NOR2x1_ASAP7_75t_L g1845 ( 
.A(n_1667),
.B(n_1419),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1545),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1545),
.Y(n_1847)
);

AOI22x1_ASAP7_75t_SL g1848 ( 
.A1(n_1522),
.A2(n_1373),
.B1(n_1385),
.B2(n_1361),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1525),
.B(n_1484),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1545),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1545),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1537),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1602),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1545),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1545),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1641),
.B(n_962),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1635),
.B(n_1484),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1602),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1545),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1545),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1545),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1602),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1545),
.Y(n_1863)
);

NAND2xp33_ASAP7_75t_L g1864 ( 
.A(n_1672),
.B(n_1501),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1545),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1517),
.A2(n_928),
.B(n_908),
.Y(n_1866)
);

AND2x6_ASAP7_75t_L g1867 ( 
.A(n_1548),
.B(n_1018),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1545),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1545),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1532),
.Y(n_1870)
);

CKINVDCx11_ASAP7_75t_R g1871 ( 
.A(n_1634),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1525),
.B(n_984),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1545),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1568),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1568),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1545),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1532),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1545),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1545),
.Y(n_1879)
);

OA22x2_ASAP7_75t_SL g1880 ( 
.A1(n_1539),
.A2(n_1472),
.B1(n_855),
.B2(n_944),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1545),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1545),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1545),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1545),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1545),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1525),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1568),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1545),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1521),
.A2(n_1468),
.B1(n_842),
.B2(n_847),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1541),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1545),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1537),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1532),
.B(n_943),
.Y(n_1893)
);

INVx6_ASAP7_75t_L g1894 ( 
.A(n_1634),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1545),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1545),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1568),
.Y(n_1897)
);

INVx5_ASAP7_75t_L g1898 ( 
.A(n_1646),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1537),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1582),
.A2(n_1090),
.B1(n_1121),
.B2(n_1074),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1545),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1541),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1568),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1545),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1568),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1545),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1545),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1517),
.A2(n_1020),
.B(n_953),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1545),
.Y(n_1909)
);

CKINVDCx11_ASAP7_75t_R g1910 ( 
.A(n_1634),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1634),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1545),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1545),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1517),
.A2(n_1088),
.B(n_1021),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1532),
.B(n_1192),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1521),
.A2(n_843),
.B1(n_858),
.B2(n_848),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1545),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1643),
.B(n_1249),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1643),
.B(n_1277),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1545),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1545),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1641),
.B(n_1117),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1541),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1541),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1545),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1514),
.A2(n_880),
.B(n_870),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1541),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1545),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1532),
.B(n_1239),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1541),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1545),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1545),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1602),
.Y(n_1933)
);

OAI21x1_ASAP7_75t_L g1934 ( 
.A1(n_1517),
.A2(n_1248),
.B(n_1240),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1545),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1541),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1545),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1541),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1532),
.B(n_1252),
.Y(n_1939)
);

OAI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1517),
.A2(n_1345),
.B(n_1301),
.Y(n_1940)
);

INVxp67_ASAP7_75t_L g1941 ( 
.A(n_1602),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1545),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1532),
.B(n_1371),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1521),
.A2(n_860),
.B1(n_863),
.B2(n_862),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1532),
.Y(n_1945)
);

CKINVDCx16_ASAP7_75t_R g1946 ( 
.A(n_1526),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1545),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1582),
.A2(n_1204),
.B1(n_1205),
.B2(n_1159),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1545),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1545),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1545),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1545),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1521),
.A2(n_1402),
.B1(n_1433),
.B2(n_1394),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1545),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1525),
.B(n_1131),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1545),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1545),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1545),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1582),
.A2(n_1235),
.B1(n_1245),
.B2(n_1221),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1641),
.B(n_1164),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1545),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1545),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1545),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1545),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1545),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1532),
.Y(n_1966)
);

OA21x2_ASAP7_75t_L g1967 ( 
.A1(n_1514),
.A2(n_887),
.B(n_885),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1545),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1525),
.B(n_1309),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1568),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1700),
.Y(n_1971)
);

NOR2xp67_ASAP7_75t_L g1972 ( 
.A(n_1696),
.B(n_912),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1754),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1711),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1822),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1785),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1877),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1945),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1750),
.B(n_1259),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1966),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1748),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1830),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1835),
.Y(n_1983)
);

CKINVDCx20_ASAP7_75t_R g1984 ( 
.A(n_1773),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1820),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1711),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1863),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1842),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1857),
.B(n_949),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1751),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1709),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1893),
.B(n_1440),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1801),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1872),
.B(n_1277),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1869),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1780),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1811),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1730),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1784),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1718),
.Y(n_2000)
);

INVxp67_ASAP7_75t_SL g2001 ( 
.A(n_1751),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1786),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_1946),
.Y(n_2003)
);

CKINVDCx20_ASAP7_75t_R g2004 ( 
.A(n_1783),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_R g2005 ( 
.A(n_1840),
.B(n_1871),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1808),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1955),
.B(n_1078),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1910),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1738),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1788),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1753),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1878),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1870),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1879),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_1726),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1793),
.Y(n_2016)
);

BUFx2_ASAP7_75t_L g2017 ( 
.A(n_1706),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1737),
.Y(n_2018)
);

AO21x2_ASAP7_75t_L g2019 ( 
.A1(n_1915),
.A2(n_898),
.B(n_890),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1900),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1844),
.Y(n_2021)
);

BUFx6f_ASAP7_75t_L g2022 ( 
.A(n_1716),
.Y(n_2022)
);

BUFx10_ASAP7_75t_L g2023 ( 
.A(n_1894),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1886),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1856),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_1736),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1922),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1960),
.Y(n_2028)
);

CKINVDCx20_ASAP7_75t_R g2029 ( 
.A(n_1948),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1929),
.B(n_1454),
.Y(n_2030)
);

INVxp67_ASAP7_75t_L g2031 ( 
.A(n_1763),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1722),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1959),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1911),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1705),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1814),
.Y(n_2036)
);

INVxp33_ASAP7_75t_L g2037 ( 
.A(n_1853),
.Y(n_2037)
);

INVxp33_ASAP7_75t_L g2038 ( 
.A(n_1858),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1698),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1702),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_R g2041 ( 
.A(n_1864),
.B(n_1336),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1724),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1799),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1802),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1969),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1790),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1939),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1882),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_1933),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1943),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1798),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1812),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1686),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1690),
.Y(n_2054)
);

BUFx10_ASAP7_75t_L g2055 ( 
.A(n_1791),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1734),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1839),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1797),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1800),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1766),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1825),
.Y(n_2061)
);

NOR2xp67_ASAP7_75t_L g2062 ( 
.A(n_1862),
.B(n_918),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1848),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1761),
.B(n_924),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1824),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1883),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1717),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1792),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_R g2069 ( 
.A(n_1795),
.B(n_1342),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_1768),
.B(n_895),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1941),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_1729),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1714),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1805),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1953),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1807),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1916),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_1746),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1890),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1944),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1821),
.Y(n_2081)
);

NOR2xp67_ASAP7_75t_L g2082 ( 
.A(n_1747),
.B(n_935),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_R g2083 ( 
.A(n_1772),
.B(n_1399),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1867),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1884),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1867),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1794),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1803),
.Y(n_2088)
);

CKINVDCx16_ASAP7_75t_R g2089 ( 
.A(n_1774),
.Y(n_2089)
);

CKINVDCx20_ASAP7_75t_R g2090 ( 
.A(n_1764),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1703),
.Y(n_2091)
);

INVxp33_ASAP7_75t_L g2092 ( 
.A(n_1837),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1834),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1947),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1806),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1952),
.Y(n_2096)
);

INVxp33_ASAP7_75t_L g2097 ( 
.A(n_1889),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1829),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1849),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1817),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1852),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_SL g2102 ( 
.A(n_1701),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1892),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1899),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1740),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1760),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_R g2107 ( 
.A(n_1779),
.B(n_1404),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1890),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1789),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1710),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_1723),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1956),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_1918),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1957),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1919),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1735),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_1836),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1958),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1735),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1962),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_1823),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1841),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1815),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1841),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_1964),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1816),
.Y(n_2126)
);

CKINVDCx20_ASAP7_75t_R g2127 ( 
.A(n_1833),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1819),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1843),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1704),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1757),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1725),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_R g2133 ( 
.A(n_1755),
.B(n_868),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1765),
.Y(n_2134)
);

NOR2x1p5_ASAP7_75t_L g2135 ( 
.A(n_1749),
.B(n_869),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1725),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_R g2137 ( 
.A(n_1804),
.B(n_938),
.Y(n_2137)
);

BUFx10_ASAP7_75t_L g2138 ( 
.A(n_1758),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1752),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1767),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1769),
.Y(n_2141)
);

CKINVDCx20_ASAP7_75t_R g2142 ( 
.A(n_1769),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1770),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1684),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1902),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1759),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1778),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1778),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1771),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1787),
.Y(n_2150)
);

CKINVDCx6p67_ASAP7_75t_R g2151 ( 
.A(n_1687),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_1845),
.Y(n_2152)
);

BUFx10_ASAP7_75t_L g2153 ( 
.A(n_1762),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1787),
.Y(n_2154)
);

CKINVDCx20_ASAP7_75t_R g2155 ( 
.A(n_1756),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_1926),
.Y(n_2156)
);

CKINVDCx16_ASAP7_75t_R g2157 ( 
.A(n_1708),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_1688),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1775),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_1874),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1902),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1728),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1739),
.Y(n_2163)
);

AOI21x1_ASAP7_75t_L g2164 ( 
.A1(n_1777),
.A2(n_906),
.B(n_901),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1739),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_1923),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1687),
.B(n_1409),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_1875),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1744),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1967),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1743),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_1809),
.B(n_940),
.Y(n_2172)
);

CKINVDCx20_ASAP7_75t_R g2173 ( 
.A(n_1880),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1810),
.Y(n_2174)
);

NOR2xp67_ASAP7_75t_L g2175 ( 
.A(n_1813),
.B(n_1827),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1838),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1745),
.Y(n_2177)
);

XNOR2xp5_ASAP7_75t_L g2178 ( 
.A(n_1796),
.B(n_1442),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1826),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1828),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1887),
.Y(n_2181)
);

CKINVDCx20_ASAP7_75t_R g2182 ( 
.A(n_1898),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1897),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1903),
.Y(n_2184)
);

CKINVDCx20_ASAP7_75t_R g2185 ( 
.A(n_1898),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_1905),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1831),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_1970),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1832),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_1924),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1697),
.Y(n_2191)
);

INVx6_ASAP7_75t_L g2192 ( 
.A(n_1924),
.Y(n_2192)
);

CKINVDCx20_ASAP7_75t_R g2193 ( 
.A(n_1713),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1719),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1927),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_R g2196 ( 
.A(n_1776),
.B(n_951),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1930),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1692),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1930),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1720),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_1936),
.Y(n_2201)
);

CKINVDCx16_ASAP7_75t_R g2202 ( 
.A(n_1936),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_1683),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1721),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1727),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_R g2206 ( 
.A(n_1866),
.B(n_872),
.Y(n_2206)
);

CKINVDCx5p33_ASAP7_75t_R g2207 ( 
.A(n_1938),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1731),
.Y(n_2208)
);

INVx4_ASAP7_75t_L g2209 ( 
.A(n_1938),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1693),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1732),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1694),
.Y(n_2212)
);

CKINVDCx20_ASAP7_75t_R g2213 ( 
.A(n_1733),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1846),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1742),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1851),
.B(n_1001),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1854),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_R g2218 ( 
.A(n_1685),
.B(n_959),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1855),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1859),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1873),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1888),
.Y(n_2222)
);

NOR2xp67_ASAP7_75t_L g2223 ( 
.A(n_1689),
.B(n_966),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_1891),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_2025),
.B(n_1092),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1992),
.B(n_1781),
.Y(n_2226)
);

CKINVDCx20_ASAP7_75t_R g2227 ( 
.A(n_1984),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1996),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_2039),
.Y(n_2229)
);

AND2x2_ASAP7_75t_SL g2230 ( 
.A(n_2089),
.B(n_855),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1999),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2030),
.B(n_1782),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_2047),
.B(n_968),
.Y(n_2233)
);

INVx4_ASAP7_75t_SL g2234 ( 
.A(n_1976),
.Y(n_2234)
);

INVx4_ASAP7_75t_SL g2235 ( 
.A(n_2102),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_L g2236 ( 
.A(n_2027),
.B(n_877),
.C(n_875),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2155),
.A2(n_996),
.B1(n_934),
.B2(n_936),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_1989),
.B(n_1162),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2156),
.A2(n_975),
.B1(n_980),
.B2(n_969),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_2142),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1991),
.B(n_1691),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2050),
.B(n_990),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_2126),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2198),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_2144),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1971),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2078),
.B(n_1847),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2002),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_2128),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_2135),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2055),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_2168),
.B(n_1850),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2170),
.A2(n_999),
.B1(n_1008),
.B2(n_992),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2217),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2040),
.B(n_1009),
.Y(n_2255)
);

INVx8_ASAP7_75t_L g2256 ( 
.A(n_1993),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2219),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1987),
.B(n_1860),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2169),
.Y(n_2259)
);

BUFx4f_ASAP7_75t_L g2260 ( 
.A(n_1979),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2028),
.B(n_2042),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2010),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2046),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2043),
.B(n_1010),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_2071),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2044),
.B(n_1818),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2064),
.B(n_1895),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2058),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2059),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1995),
.B(n_1861),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2074),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2076),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1974),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2081),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2019),
.B(n_1896),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1988),
.Y(n_2276)
);

INVx4_ASAP7_75t_L g2277 ( 
.A(n_2130),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2191),
.Y(n_2278)
);

BUFx4f_ASAP7_75t_L g2279 ( 
.A(n_1979),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_1974),
.Y(n_2280)
);

INVx1_ASAP7_75t_SL g2281 ( 
.A(n_2049),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_L g2282 ( 
.A(n_2087),
.B(n_881),
.C(n_878),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_2202),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2177),
.B(n_1906),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2194),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2200),
.Y(n_2286)
);

INVx5_ASAP7_75t_L g2287 ( 
.A(n_2023),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2204),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2205),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2179),
.Y(n_2290)
);

INVx4_ASAP7_75t_SL g2291 ( 
.A(n_2102),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_2192),
.Y(n_2292)
);

INVx3_ASAP7_75t_L g2293 ( 
.A(n_2192),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2208),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2180),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2007),
.B(n_1161),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2211),
.Y(n_2297)
);

OR2x6_ASAP7_75t_L g2298 ( 
.A(n_2017),
.B(n_2152),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2187),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2097),
.B(n_1208),
.Y(n_2300)
);

INVx4_ASAP7_75t_L g2301 ( 
.A(n_2131),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2083),
.B(n_1014),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2036),
.B(n_1236),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2215),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2189),
.Y(n_2305)
);

AOI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2092),
.A2(n_2146),
.B1(n_2149),
.B2(n_2139),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2216),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_L g2308 ( 
.A1(n_2159),
.A2(n_925),
.B1(n_1118),
.B2(n_1057),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1990),
.Y(n_2309)
);

NOR2x1p5_ASAP7_75t_L g2310 ( 
.A(n_2018),
.B(n_884),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_1974),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2012),
.B(n_2014),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2026),
.B(n_1282),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2134),
.B(n_1175),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_1986),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2216),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_2031),
.B(n_1295),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2158),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2160),
.Y(n_2319)
);

NAND2x1p5_ASAP7_75t_L g2320 ( 
.A(n_2188),
.B(n_1865),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2186),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2210),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2173),
.A2(n_937),
.B1(n_948),
.B2(n_921),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1990),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2001),
.B(n_1907),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2132),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2212),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2214),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2054),
.B(n_1312),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2220),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2136),
.Y(n_2331)
);

AO22x2_ASAP7_75t_L g2332 ( 
.A1(n_1994),
.A2(n_1324),
.B1(n_1486),
.B2(n_1401),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2221),
.Y(n_2333)
);

AND2x6_ASAP7_75t_L g2334 ( 
.A(n_2070),
.B(n_944),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2037),
.B(n_896),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2048),
.B(n_1868),
.Y(n_2336)
);

BUFx3_ASAP7_75t_L g2337 ( 
.A(n_2162),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2163),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_2022),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2222),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2022),
.Y(n_2341)
);

BUFx10_ASAP7_75t_L g2342 ( 
.A(n_2008),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1972),
.B(n_2224),
.Y(n_2343)
);

AND2x6_ASAP7_75t_L g2344 ( 
.A(n_2066),
.B(n_1493),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2045),
.Y(n_2345)
);

INVx2_ASAP7_75t_SL g2346 ( 
.A(n_2140),
.Y(n_2346)
);

AO21x2_ASAP7_75t_L g2347 ( 
.A1(n_2041),
.A2(n_1914),
.B(n_1908),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2038),
.B(n_886),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_2032),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2201),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2141),
.B(n_1197),
.Y(n_2351)
);

INVx5_ASAP7_75t_L g2352 ( 
.A(n_2032),
.Y(n_2352)
);

INVx3_ASAP7_75t_L g2353 ( 
.A(n_2032),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2057),
.B(n_889),
.Y(n_2354)
);

AND2x6_ASAP7_75t_L g2355 ( 
.A(n_2085),
.B(n_1493),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_1973),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2143),
.B(n_1016),
.Y(n_2357)
);

AND2x2_ASAP7_75t_SL g2358 ( 
.A(n_2157),
.B(n_837),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2203),
.Y(n_2359)
);

AO22x2_ASAP7_75t_L g2360 ( 
.A1(n_2073),
.A2(n_917),
.B1(n_1167),
.B2(n_1062),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2108),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2121),
.B(n_893),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2125),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2108),
.Y(n_2364)
);

BUFx10_ASAP7_75t_L g2365 ( 
.A(n_2021),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2165),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2082),
.B(n_1917),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2094),
.B(n_1876),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2079),
.Y(n_2369)
);

AND2x6_ASAP7_75t_L g2370 ( 
.A(n_2096),
.B(n_1003),
.Y(n_2370)
);

AND2x6_ASAP7_75t_L g2371 ( 
.A(n_2112),
.B(n_1006),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2079),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2166),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2166),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2199),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2174),
.B(n_1920),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2147),
.B(n_1019),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2065),
.B(n_1233),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2176),
.B(n_1921),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2127),
.B(n_900),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2088),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2095),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2024),
.B(n_1315),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2148),
.B(n_2150),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2108),
.Y(n_2385)
);

BUFx4f_ASAP7_75t_L g2386 ( 
.A(n_2151),
.Y(n_2386)
);

INVx3_ASAP7_75t_L g2387 ( 
.A(n_2145),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2145),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2077),
.B(n_904),
.Y(n_2389)
);

OR2x6_ASAP7_75t_L g2390 ( 
.A(n_2114),
.B(n_1489),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2161),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2080),
.B(n_905),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2129),
.B(n_907),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2161),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2223),
.B(n_1928),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2154),
.B(n_1279),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2118),
.B(n_1881),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2009),
.B(n_910),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2123),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2033),
.B(n_914),
.Y(n_2400)
);

AND2x6_ASAP7_75t_L g2401 ( 
.A(n_2120),
.B(n_1017),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2069),
.B(n_1036),
.Y(n_2402)
);

AND2x2_ASAP7_75t_SL g2403 ( 
.A(n_2067),
.B(n_915),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2062),
.B(n_1942),
.Y(n_2404)
);

BUFx10_ASAP7_75t_L g2405 ( 
.A(n_1981),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1975),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2196),
.B(n_1949),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_1982),
.B(n_1885),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2161),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2122),
.B(n_2124),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1983),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2164),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2011),
.B(n_1951),
.Y(n_2413)
);

INVx4_ASAP7_75t_L g2414 ( 
.A(n_2171),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2209),
.Y(n_2415)
);

INVxp67_ASAP7_75t_SL g2416 ( 
.A(n_2175),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2209),
.Y(n_2417)
);

INVx2_ASAP7_75t_SL g2418 ( 
.A(n_2138),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2013),
.B(n_1954),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2138),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2190),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2195),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2300),
.A2(n_2091),
.B1(n_2178),
.B2(n_2029),
.Y(n_2423)
);

AO22x2_ASAP7_75t_L g2424 ( 
.A1(n_2237),
.A2(n_1039),
.B1(n_1045),
.B2(n_1023),
.Y(n_2424)
);

INVxp67_ASAP7_75t_L g2425 ( 
.A(n_2238),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2273),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2228),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2231),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2229),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2248),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2265),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2225),
.B(n_2016),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2244),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2262),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2303),
.B(n_1977),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2263),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2268),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2269),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_SL g2439 ( 
.A1(n_2403),
.A2(n_2075),
.B1(n_2020),
.B2(n_2090),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2266),
.B(n_2107),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2273),
.Y(n_2441)
);

AO22x2_ASAP7_75t_L g2442 ( 
.A1(n_2400),
.A2(n_1059),
.B1(n_1060),
.B2(n_1056),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2271),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2254),
.Y(n_2444)
);

INVxp67_ASAP7_75t_SL g2445 ( 
.A(n_2280),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_2240),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2257),
.Y(n_2447)
);

AOI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2389),
.A2(n_2133),
.B1(n_2115),
.B2(n_2113),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2359),
.B(n_2000),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2246),
.Y(n_2450)
);

AO22x2_ASAP7_75t_L g2451 ( 
.A1(n_2281),
.A2(n_1071),
.B1(n_1072),
.B2(n_1070),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2261),
.B(n_2313),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2272),
.Y(n_2453)
);

NAND2x1p5_ASAP7_75t_L g2454 ( 
.A(n_2301),
.B(n_1961),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2274),
.Y(n_2455)
);

AOI22x1_ASAP7_75t_L g2456 ( 
.A1(n_2276),
.A2(n_2098),
.B1(n_2119),
.B2(n_2116),
.Y(n_2456)
);

AND2x4_ASAP7_75t_SL g2457 ( 
.A(n_2365),
.B(n_2004),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_2356),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2329),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2278),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2317),
.B(n_2006),
.Y(n_2461)
);

A2O1A1Ixp33_ASAP7_75t_L g2462 ( 
.A1(n_2226),
.A2(n_2068),
.B(n_2086),
.C(n_2084),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2392),
.A2(n_2206),
.B1(n_2035),
.B2(n_2072),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2232),
.B(n_2105),
.Y(n_2464)
);

INVxp67_ASAP7_75t_L g2465 ( 
.A(n_2296),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2285),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2286),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2283),
.B(n_2197),
.Y(n_2468)
);

NOR2xp67_ASAP7_75t_L g2469 ( 
.A(n_2287),
.B(n_1978),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2243),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2288),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2267),
.B(n_2106),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2289),
.Y(n_2473)
);

NAND2xp33_ASAP7_75t_L g2474 ( 
.A(n_2343),
.B(n_1980),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2294),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2297),
.Y(n_2476)
);

AO22x2_ASAP7_75t_L g2477 ( 
.A1(n_2323),
.A2(n_2236),
.B1(n_2378),
.B2(n_2327),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2304),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2259),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2284),
.Y(n_2480)
);

BUFx8_ASAP7_75t_L g2481 ( 
.A(n_2249),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2416),
.B(n_2109),
.Y(n_2482)
);

NOR2xp67_ASAP7_75t_L g2483 ( 
.A(n_2277),
.B(n_1985),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2234),
.B(n_2207),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2348),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2290),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2398),
.B(n_2100),
.Y(n_2487)
);

AND2x4_ASAP7_75t_L g2488 ( 
.A(n_2235),
.B(n_2003),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2239),
.A2(n_2111),
.B1(n_2110),
.B2(n_2117),
.Y(n_2489)
);

OAI21xp33_ASAP7_75t_L g2490 ( 
.A1(n_2393),
.A2(n_2354),
.B(n_2306),
.Y(n_2490)
);

AO22x2_ASAP7_75t_L g2491 ( 
.A1(n_2322),
.A2(n_1086),
.B1(n_1087),
.B2(n_1081),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2253),
.A2(n_2052),
.B1(n_2051),
.B2(n_2101),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2260),
.A2(n_2034),
.B1(n_2099),
.B2(n_2103),
.Y(n_2493)
);

AO22x2_ASAP7_75t_L g2494 ( 
.A1(n_2328),
.A2(n_2015),
.B1(n_1110),
.B2(n_1119),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2307),
.Y(n_2495)
);

AO22x2_ASAP7_75t_L g2496 ( 
.A1(n_2330),
.A2(n_1123),
.B1(n_1128),
.B2(n_1093),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2295),
.Y(n_2497)
);

OAI22xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2227),
.A2(n_2056),
.B1(n_2061),
.B2(n_2060),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2299),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2316),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2305),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2291),
.B(n_2053),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2334),
.A2(n_994),
.B1(n_1015),
.B2(n_1002),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2314),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2334),
.A2(n_1031),
.B1(n_1037),
.B2(n_1033),
.Y(n_2505)
);

NAND2x1p5_ASAP7_75t_L g2506 ( 
.A(n_2414),
.B(n_1901),
.Y(n_2506)
);

BUFx3_ASAP7_75t_L g2507 ( 
.A(n_2337),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2366),
.B(n_2104),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2376),
.B(n_2181),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2258),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2270),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2362),
.B(n_2183),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2336),
.Y(n_2513)
);

NAND2x1p5_ASAP7_75t_L g2514 ( 
.A(n_2422),
.B(n_1904),
.Y(n_2514)
);

NAND2x1p5_ASAP7_75t_L g2515 ( 
.A(n_2384),
.B(n_1909),
.Y(n_2515)
);

INVxp67_ASAP7_75t_SL g2516 ( 
.A(n_2280),
.Y(n_2516)
);

NAND2x1p5_ASAP7_75t_L g2517 ( 
.A(n_2346),
.B(n_1912),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2368),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2397),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2245),
.B(n_2193),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2379),
.B(n_2184),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2369),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2413),
.B(n_2137),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2326),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2241),
.B(n_2213),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2373),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2374),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2380),
.B(n_2153),
.Y(n_2528)
);

AO22x2_ASAP7_75t_L g2529 ( 
.A1(n_2333),
.A2(n_1136),
.B1(n_1138),
.B2(n_1134),
.Y(n_2529)
);

AO22x2_ASAP7_75t_L g2530 ( 
.A1(n_2340),
.A2(n_1142),
.B1(n_1147),
.B2(n_1139),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2331),
.Y(n_2531)
);

AND2x6_ASAP7_75t_L g2532 ( 
.A(n_2420),
.B(n_1064),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2419),
.B(n_2172),
.Y(n_2533)
);

NAND2x1_ASAP7_75t_L g2534 ( 
.A(n_2412),
.B(n_1913),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2338),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2309),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2324),
.Y(n_2537)
);

INVx6_ASAP7_75t_L g2538 ( 
.A(n_2256),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2408),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2391),
.Y(n_2540)
);

INVx4_ASAP7_75t_L g2541 ( 
.A(n_2352),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2404),
.B(n_2153),
.Y(n_2542)
);

INVx8_ASAP7_75t_L g2543 ( 
.A(n_2352),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2233),
.B(n_2242),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2409),
.Y(n_2545)
);

INVxp67_ASAP7_75t_SL g2546 ( 
.A(n_2311),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2275),
.B(n_2218),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_2350),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2358),
.B(n_2005),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2282),
.A2(n_2250),
.B1(n_2279),
.B2(n_2230),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2372),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2375),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2247),
.B(n_2182),
.Y(n_2553)
);

BUFx2_ASAP7_75t_L g2554 ( 
.A(n_2345),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_2418),
.B(n_1997),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2325),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2292),
.B(n_2185),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2308),
.A2(n_1085),
.B1(n_1111),
.B2(n_1091),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2381),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2293),
.B(n_1998),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2382),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2255),
.B(n_1113),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2399),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_2332),
.A2(n_1115),
.B1(n_1126),
.B2(n_1125),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2264),
.B(n_1130),
.Y(n_2565)
);

AO22x2_ASAP7_75t_L g2566 ( 
.A1(n_2383),
.A2(n_1158),
.B1(n_1168),
.B2(n_1152),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2415),
.B(n_1132),
.Y(n_2567)
);

OR2x2_ASAP7_75t_SL g2568 ( 
.A(n_2421),
.B(n_2335),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2417),
.B(n_1151),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2406),
.Y(n_2570)
);

OR2x2_ASAP7_75t_SL g2571 ( 
.A(n_2363),
.B(n_927),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2351),
.B(n_2167),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2318),
.Y(n_2573)
);

OR2x2_ASAP7_75t_SL g2574 ( 
.A(n_2319),
.B(n_982),
.Y(n_2574)
);

INVx2_ASAP7_75t_SL g2575 ( 
.A(n_2252),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2411),
.Y(n_2576)
);

INVx2_ASAP7_75t_SL g2577 ( 
.A(n_2396),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2321),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2315),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2367),
.A2(n_1170),
.B1(n_1179),
.B2(n_1166),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2347),
.A2(n_1185),
.B1(n_1186),
.B2(n_1183),
.Y(n_2581)
);

INVx4_ASAP7_75t_L g2582 ( 
.A(n_2311),
.Y(n_2582)
);

BUFx6f_ASAP7_75t_L g2583 ( 
.A(n_2426),
.Y(n_2583)
);

NOR3xp33_ASAP7_75t_L g2584 ( 
.A(n_2432),
.B(n_2410),
.C(n_2357),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2452),
.B(n_2480),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2453),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2460),
.Y(n_2587)
);

OAI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2547),
.A2(n_2395),
.B(n_2402),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2490),
.A2(n_2302),
.B1(n_2407),
.B2(n_2377),
.Y(n_2589)
);

AOI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2534),
.A2(n_1940),
.B(n_1934),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2426),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2544),
.A2(n_2556),
.B(n_2533),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2435),
.B(n_2251),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2523),
.A2(n_2320),
.B(n_2339),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2485),
.B(n_2339),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2440),
.B(n_2387),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_L g2597 ( 
.A(n_2543),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2509),
.A2(n_2349),
.B(n_2341),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2521),
.A2(n_2361),
.B(n_2353),
.Y(n_2599)
);

BUFx12f_ASAP7_75t_L g2600 ( 
.A(n_2481),
.Y(n_2600)
);

A2O1A1Ixp33_ASAP7_75t_L g2601 ( 
.A1(n_2528),
.A2(n_1212),
.B(n_1214),
.C(n_1187),
.Y(n_2601)
);

A2O1A1Ixp33_ASAP7_75t_L g2602 ( 
.A1(n_2448),
.A2(n_1219),
.B(n_1226),
.C(n_1216),
.Y(n_2602)
);

OAI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2581),
.A2(n_2312),
.B(n_1260),
.Y(n_2603)
);

OAI321xp33_ASAP7_75t_L g2604 ( 
.A1(n_2564),
.A2(n_2423),
.A3(n_2425),
.B1(n_2463),
.B2(n_2461),
.C(n_2503),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2427),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2464),
.B(n_2388),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2449),
.B(n_2360),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2487),
.B(n_2394),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2470),
.Y(n_2609)
);

OAI21xp33_ASAP7_75t_L g2610 ( 
.A1(n_2512),
.A2(n_1482),
.B(n_2298),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2542),
.A2(n_2385),
.B(n_2364),
.Y(n_2611)
);

AOI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2477),
.A2(n_2310),
.B1(n_2093),
.B2(n_1038),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2472),
.B(n_1695),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2431),
.B(n_2390),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2428),
.B(n_1699),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2459),
.B(n_2405),
.Y(n_2616)
);

AO21x2_ASAP7_75t_L g2617 ( 
.A1(n_2567),
.A2(n_1304),
.B(n_1263),
.Y(n_2617)
);

AOI221x1_ASAP7_75t_L g2618 ( 
.A1(n_2477),
.A2(n_1319),
.B1(n_1320),
.B2(n_1316),
.C(n_1308),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2473),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2569),
.A2(n_1004),
.B(n_941),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2430),
.B(n_1707),
.Y(n_2621)
);

A2O1A1Ixp33_ASAP7_75t_L g2622 ( 
.A1(n_2478),
.A2(n_1335),
.B(n_1338),
.C(n_1323),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2434),
.B(n_1712),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2436),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2437),
.Y(n_2625)
);

O2A1O1Ixp33_ASAP7_75t_L g2626 ( 
.A1(n_2462),
.A2(n_1359),
.B(n_1369),
.C(n_1347),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2438),
.Y(n_2627)
);

CKINVDCx8_ASAP7_75t_R g2628 ( 
.A(n_2450),
.Y(n_2628)
);

NAND2x1p5_ASAP7_75t_L g2629 ( 
.A(n_2507),
.B(n_2386),
.Y(n_2629)
);

INVx4_ASAP7_75t_L g2630 ( 
.A(n_2543),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2482),
.A2(n_1004),
.B(n_941),
.Y(n_2631)
);

A2O1A1Ixp33_ASAP7_75t_L g2632 ( 
.A1(n_2443),
.A2(n_1382),
.B(n_1383),
.C(n_1381),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2455),
.B(n_1715),
.Y(n_2633)
);

O2A1O1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2465),
.A2(n_1420),
.B(n_1432),
.C(n_1407),
.Y(n_2634)
);

AO21x2_ASAP7_75t_L g2635 ( 
.A1(n_2562),
.A2(n_1437),
.B(n_1435),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_L g2636 ( 
.A(n_2429),
.B(n_2342),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2433),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2466),
.B(n_1741),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2467),
.B(n_2344),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2471),
.B(n_2344),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2484),
.B(n_2355),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2504),
.B(n_2063),
.Y(n_2642)
);

OAI21xp33_ASAP7_75t_L g2643 ( 
.A1(n_2578),
.A2(n_922),
.B(n_916),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2444),
.A2(n_1004),
.B(n_941),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2483),
.B(n_1409),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2447),
.A2(n_1073),
.B(n_1004),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2479),
.A2(n_2497),
.B(n_2486),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2572),
.B(n_2355),
.Y(n_2648)
);

AOI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2499),
.A2(n_1124),
.B(n_1073),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2475),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2501),
.A2(n_1124),
.B(n_1073),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2476),
.A2(n_1461),
.B1(n_1462),
.B2(n_1450),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2565),
.A2(n_1242),
.B(n_1124),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2495),
.Y(n_2654)
);

BUFx2_ASAP7_75t_L g2655 ( 
.A(n_2525),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2576),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2500),
.B(n_1925),
.Y(n_2657)
);

OAI21xp33_ASAP7_75t_L g2658 ( 
.A1(n_2573),
.A2(n_2548),
.B(n_2577),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2559),
.B(n_1931),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2561),
.B(n_1932),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2474),
.A2(n_2552),
.B(n_2551),
.Y(n_2661)
);

AOI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2540),
.A2(n_1937),
.B(n_1935),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2458),
.B(n_1473),
.Y(n_2663)
);

O2A1O1Ixp33_ASAP7_75t_SL g2664 ( 
.A1(n_2522),
.A2(n_2527),
.B(n_2526),
.C(n_2545),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2524),
.A2(n_1291),
.B(n_1242),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2446),
.Y(n_2666)
);

OAI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2563),
.A2(n_1470),
.B1(n_1475),
.B2(n_1464),
.Y(n_2667)
);

AOI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2445),
.A2(n_1291),
.B(n_1242),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2570),
.Y(n_2669)
);

NOR3xp33_ASAP7_75t_L g2670 ( 
.A(n_2439),
.B(n_930),
.C(n_929),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2531),
.B(n_1950),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2575),
.B(n_2539),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2538),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2516),
.A2(n_1291),
.B(n_1242),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2546),
.A2(n_1337),
.B(n_1291),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2554),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2508),
.B(n_2370),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2456),
.A2(n_1487),
.B1(n_1492),
.B2(n_1476),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2535),
.B(n_1963),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2536),
.B(n_1965),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2550),
.A2(n_1502),
.B1(n_1508),
.B2(n_1495),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2537),
.B(n_1968),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2469),
.B(n_1473),
.Y(n_2683)
);

BUFx4f_ASAP7_75t_L g2684 ( 
.A(n_2488),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2510),
.A2(n_1384),
.B(n_1337),
.Y(n_2685)
);

O2A1O1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2493),
.A2(n_1174),
.B(n_1178),
.C(n_1173),
.Y(n_2686)
);

AOI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2511),
.A2(n_1384),
.B(n_1337),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2520),
.B(n_2370),
.Y(n_2688)
);

A2O1A1Ixp33_ASAP7_75t_L g2689 ( 
.A1(n_2580),
.A2(n_1203),
.B(n_1206),
.C(n_1196),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2579),
.Y(n_2690)
);

AOI21xp5_ASAP7_75t_L g2691 ( 
.A1(n_2513),
.A2(n_1384),
.B(n_1498),
.Y(n_2691)
);

AOI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2489),
.A2(n_1513),
.B1(n_1512),
.B2(n_1080),
.Y(n_2692)
);

AOI21x1_ASAP7_75t_L g2693 ( 
.A1(n_2518),
.A2(n_1210),
.B(n_1207),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2424),
.B(n_2558),
.Y(n_2694)
);

AOI21xp5_ASAP7_75t_L g2695 ( 
.A1(n_2519),
.A2(n_1096),
.B(n_1094),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2442),
.B(n_2371),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_2492),
.B(n_2549),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2505),
.A2(n_1100),
.B1(n_1103),
.B2(n_1099),
.Y(n_2698)
);

AOI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2515),
.A2(n_1112),
.B(n_1109),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2568),
.B(n_946),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2585),
.B(n_2457),
.Y(n_2701)
);

A2O1A1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2592),
.A2(n_2555),
.B(n_2441),
.C(n_2468),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2650),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2605),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2673),
.Y(n_2705)
);

AND2x4_ASAP7_75t_SL g2706 ( 
.A(n_2673),
.B(n_2502),
.Y(n_2706)
);

A2O1A1Ixp33_ASAP7_75t_L g2707 ( 
.A1(n_2604),
.A2(n_1250),
.B(n_1254),
.C(n_1228),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2593),
.B(n_2532),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2624),
.Y(n_2709)
);

BUFx8_ASAP7_75t_L g2710 ( 
.A(n_2600),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2697),
.A2(n_2498),
.B1(n_2553),
.B2(n_2557),
.Y(n_2711)
);

AOI21x1_ASAP7_75t_L g2712 ( 
.A1(n_2662),
.A2(n_2496),
.B(n_2491),
.Y(n_2712)
);

OAI21xp33_ASAP7_75t_SL g2713 ( 
.A1(n_2589),
.A2(n_2582),
.B(n_2541),
.Y(n_2713)
);

OAI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2625),
.A2(n_2574),
.B1(n_2571),
.B2(n_2506),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2666),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2588),
.A2(n_2514),
.B(n_2454),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2627),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2610),
.B(n_2517),
.Y(n_2718)
);

INVx4_ASAP7_75t_L g2719 ( 
.A(n_2666),
.Y(n_2719)
);

BUFx6f_ASAP7_75t_L g2720 ( 
.A(n_2583),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2608),
.A2(n_2442),
.B(n_2530),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2606),
.B(n_2532),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2584),
.B(n_2491),
.Y(n_2723)
);

BUFx2_ASAP7_75t_L g2724 ( 
.A(n_2676),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2596),
.B(n_2496),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2613),
.A2(n_2529),
.B(n_2566),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2628),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2648),
.B(n_2566),
.Y(n_2728)
);

NOR3xp33_ASAP7_75t_L g2729 ( 
.A(n_2663),
.B(n_2560),
.C(n_1465),
.Y(n_2729)
);

INVx1_ASAP7_75t_SL g2730 ( 
.A(n_2609),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2669),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2594),
.A2(n_2529),
.B(n_1135),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2654),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2586),
.Y(n_2734)
);

BUFx2_ASAP7_75t_SL g2735 ( 
.A(n_2630),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2661),
.A2(n_1143),
.B(n_1129),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2587),
.A2(n_2494),
.B1(n_2451),
.B2(n_1146),
.Y(n_2737)
);

INVxp67_ASAP7_75t_L g2738 ( 
.A(n_2636),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2619),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2656),
.B(n_2451),
.Y(n_2740)
);

O2A1O1Ixp33_ASAP7_75t_L g2741 ( 
.A1(n_2601),
.A2(n_1257),
.B(n_1266),
.C(n_1256),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2694),
.B(n_2401),
.Y(n_2742)
);

AO21x2_ASAP7_75t_L g2743 ( 
.A1(n_2631),
.A2(n_2599),
.B(n_2602),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2607),
.B(n_2401),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2658),
.B(n_1279),
.Y(n_2745)
);

AOI21x1_ASAP7_75t_L g2746 ( 
.A1(n_2590),
.A2(n_1287),
.B(n_1284),
.Y(n_2746)
);

BUFx2_ASAP7_75t_L g2747 ( 
.A(n_2591),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2616),
.B(n_1306),
.Y(n_2748)
);

AND2x2_ASAP7_75t_SL g2749 ( 
.A(n_2670),
.B(n_1297),
.Y(n_2749)
);

AOI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2603),
.A2(n_1156),
.B(n_1155),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2597),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2637),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2642),
.B(n_1306),
.Y(n_2753)
);

AND2x6_ASAP7_75t_L g2754 ( 
.A(n_2696),
.B(n_1310),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2690),
.Y(n_2755)
);

O2A1O1Ixp5_ASAP7_75t_L g2756 ( 
.A1(n_2681),
.A2(n_1358),
.B(n_1363),
.C(n_1354),
.Y(n_2756)
);

AND2x4_ASAP7_75t_L g2757 ( 
.A(n_2641),
.B(n_1365),
.Y(n_2757)
);

CKINVDCx20_ASAP7_75t_R g2758 ( 
.A(n_2655),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2700),
.B(n_950),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2614),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2598),
.A2(n_1177),
.B(n_1171),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2659),
.B(n_1157),
.Y(n_2762)
);

O2A1O1Ixp33_ASAP7_75t_L g2763 ( 
.A1(n_2686),
.A2(n_1378),
.B(n_1393),
.C(n_1372),
.Y(n_2763)
);

O2A1O1Ixp33_ASAP7_75t_L g2764 ( 
.A1(n_2645),
.A2(n_1405),
.B(n_1406),
.C(n_1400),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2641),
.Y(n_2765)
);

O2A1O1Ixp33_ASAP7_75t_L g2766 ( 
.A1(n_2678),
.A2(n_1417),
.B(n_1418),
.C(n_1410),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2647),
.A2(n_1209),
.B(n_1182),
.Y(n_2767)
);

OR2x6_ASAP7_75t_L g2768 ( 
.A(n_2629),
.B(n_1424),
.Y(n_2768)
);

O2A1O1Ixp33_ASAP7_75t_L g2769 ( 
.A1(n_2634),
.A2(n_1426),
.B(n_1427),
.C(n_1425),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2660),
.B(n_1199),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2672),
.B(n_1343),
.Y(n_2771)
);

INVx6_ASAP7_75t_L g2772 ( 
.A(n_2677),
.Y(n_2772)
);

O2A1O1Ixp33_ASAP7_75t_L g2773 ( 
.A1(n_2683),
.A2(n_1448),
.B(n_1451),
.C(n_1429),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_2684),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2664),
.A2(n_1230),
.B(n_1223),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2657),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2615),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2688),
.Y(n_2778)
);

BUFx12f_ASAP7_75t_L g2779 ( 
.A(n_2672),
.Y(n_2779)
);

O2A1O1Ixp33_ASAP7_75t_L g2780 ( 
.A1(n_2595),
.A2(n_2626),
.B(n_2689),
.C(n_2632),
.Y(n_2780)
);

O2A1O1Ixp33_ASAP7_75t_L g2781 ( 
.A1(n_2622),
.A2(n_1474),
.B(n_1481),
.C(n_1459),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2621),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2639),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2693),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2640),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2612),
.B(n_952),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2692),
.B(n_954),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2643),
.A2(n_1127),
.B1(n_1200),
.B2(n_883),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2698),
.A2(n_1200),
.B1(n_1224),
.B2(n_1127),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2623),
.Y(n_2790)
);

CKINVDCx20_ASAP7_75t_R g2791 ( 
.A(n_2680),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2633),
.B(n_1241),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2638),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2611),
.B(n_1243),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2671),
.B(n_1244),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_L g2796 ( 
.A(n_2679),
.B(n_955),
.Y(n_2796)
);

OR2x2_ASAP7_75t_L g2797 ( 
.A(n_2682),
.B(n_964),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2695),
.B(n_970),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2618),
.B(n_1247),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_SL g2800 ( 
.A1(n_2652),
.A2(n_972),
.B1(n_973),
.B2(n_971),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2699),
.B(n_1267),
.Y(n_2801)
);

NAND3xp33_ASAP7_75t_SL g2802 ( 
.A(n_2691),
.B(n_2667),
.C(n_976),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2635),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2620),
.A2(n_1278),
.B(n_1275),
.Y(n_2804)
);

AOI21x1_ASAP7_75t_L g2805 ( 
.A1(n_2668),
.A2(n_1485),
.B(n_1007),
.Y(n_2805)
);

A2O1A1Ixp33_ASAP7_75t_L g2806 ( 
.A1(n_2685),
.A2(n_1032),
.B(n_1041),
.C(n_989),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2617),
.Y(n_2807)
);

OAI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2687),
.A2(n_1293),
.B(n_1283),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2674),
.B(n_1298),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2675),
.B(n_1300),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2776),
.B(n_974),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2715),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2704),
.Y(n_2813)
);

INVx1_ASAP7_75t_SL g2814 ( 
.A(n_2724),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2777),
.B(n_977),
.Y(n_2815)
);

INVx4_ASAP7_75t_L g2816 ( 
.A(n_2720),
.Y(n_2816)
);

INVx8_ASAP7_75t_L g2817 ( 
.A(n_2720),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2727),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2782),
.B(n_978),
.Y(n_2819)
);

BUFx12f_ASAP7_75t_L g2820 ( 
.A(n_2710),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2747),
.Y(n_2821)
);

NAND2x1p5_ASAP7_75t_L g2822 ( 
.A(n_2719),
.B(n_2730),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2728),
.B(n_1302),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2790),
.B(n_983),
.Y(n_2824)
);

INVx4_ASAP7_75t_L g2825 ( 
.A(n_2774),
.Y(n_2825)
);

BUFx3_ASAP7_75t_L g2826 ( 
.A(n_2705),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2791),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2706),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2793),
.B(n_985),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2709),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2731),
.Y(n_2831)
);

BUFx12f_ASAP7_75t_L g2832 ( 
.A(n_2778),
.Y(n_2832)
);

INVx2_ASAP7_75t_SL g2833 ( 
.A(n_2772),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2765),
.Y(n_2834)
);

INVx6_ASAP7_75t_L g2835 ( 
.A(n_2779),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2717),
.Y(n_2836)
);

CKINVDCx8_ASAP7_75t_R g2837 ( 
.A(n_2735),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2733),
.Y(n_2838)
);

INVx4_ASAP7_75t_L g2839 ( 
.A(n_2751),
.Y(n_2839)
);

INVx5_ASAP7_75t_L g2840 ( 
.A(n_2768),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2703),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2701),
.B(n_1314),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2734),
.Y(n_2843)
);

INVx4_ASAP7_75t_L g2844 ( 
.A(n_2772),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_L g2845 ( 
.A(n_2785),
.Y(n_2845)
);

INVx4_ASAP7_75t_L g2846 ( 
.A(n_2785),
.Y(n_2846)
);

BUFx6f_ASAP7_75t_L g2847 ( 
.A(n_2757),
.Y(n_2847)
);

BUFx5_ASAP7_75t_L g2848 ( 
.A(n_2803),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2739),
.Y(n_2849)
);

INVx3_ASAP7_75t_L g2850 ( 
.A(n_2755),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2752),
.Y(n_2851)
);

BUFx8_ASAP7_75t_L g2852 ( 
.A(n_2744),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2768),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2758),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2740),
.Y(n_2855)
);

BUFx3_ASAP7_75t_L g2856 ( 
.A(n_2760),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2725),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2784),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2783),
.Y(n_2859)
);

INVx8_ASAP7_75t_L g2860 ( 
.A(n_2754),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2754),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2807),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2754),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2742),
.Y(n_2864)
);

BUFx6f_ASAP7_75t_L g2865 ( 
.A(n_2771),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2786),
.A2(n_1200),
.B1(n_1224),
.B2(n_1127),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2712),
.Y(n_2867)
);

BUFx6f_ASAP7_75t_L g2868 ( 
.A(n_2708),
.Y(n_2868)
);

INVx6_ASAP7_75t_SL g2869 ( 
.A(n_2738),
.Y(n_2869)
);

INVx3_ASAP7_75t_L g2870 ( 
.A(n_2797),
.Y(n_2870)
);

INVx4_ASAP7_75t_L g2871 ( 
.A(n_2749),
.Y(n_2871)
);

INVx4_ASAP7_75t_L g2872 ( 
.A(n_2787),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2722),
.Y(n_2873)
);

INVx5_ASAP7_75t_L g2874 ( 
.A(n_2729),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2805),
.Y(n_2875)
);

BUFx3_ASAP7_75t_L g2876 ( 
.A(n_2711),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2796),
.B(n_1317),
.Y(n_2877)
);

CKINVDCx11_ASAP7_75t_R g2878 ( 
.A(n_2737),
.Y(n_2878)
);

INVx2_ASAP7_75t_SL g2879 ( 
.A(n_2748),
.Y(n_2879)
);

BUFx12f_ASAP7_75t_L g2880 ( 
.A(n_2702),
.Y(n_2880)
);

BUFx12f_ASAP7_75t_L g2881 ( 
.A(n_2713),
.Y(n_2881)
);

INVx4_ASAP7_75t_L g2882 ( 
.A(n_2743),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2723),
.Y(n_2883)
);

INVx1_ASAP7_75t_SL g2884 ( 
.A(n_2745),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2756),
.Y(n_2885)
);

HB1xp67_ASAP7_75t_L g2886 ( 
.A(n_2714),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2746),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2792),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2759),
.Y(n_2889)
);

INVx4_ASAP7_75t_L g2890 ( 
.A(n_2718),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2781),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2741),
.Y(n_2892)
);

INVx8_ASAP7_75t_L g2893 ( 
.A(n_2806),
.Y(n_2893)
);

BUFx12f_ASAP7_75t_L g2894 ( 
.A(n_2753),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2726),
.B(n_987),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2707),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2766),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2794),
.Y(n_2898)
);

HB1xp67_ASAP7_75t_L g2899 ( 
.A(n_2721),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2762),
.Y(n_2900)
);

AO21x2_ASAP7_75t_L g2901 ( 
.A1(n_2887),
.A2(n_2716),
.B(n_2875),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2836),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2838),
.Y(n_2903)
);

HB1xp67_ASAP7_75t_L g2904 ( 
.A(n_2859),
.Y(n_2904)
);

OAI21x1_ASAP7_75t_SL g2905 ( 
.A1(n_2890),
.A2(n_2732),
.B(n_2780),
.Y(n_2905)
);

OAI21x1_ASAP7_75t_L g2906 ( 
.A1(n_2867),
.A2(n_2651),
.B(n_2653),
.Y(n_2906)
);

AO31x2_ASAP7_75t_L g2907 ( 
.A1(n_2882),
.A2(n_2799),
.A3(n_2775),
.B(n_2649),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2888),
.B(n_2770),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2856),
.Y(n_2909)
);

AO31x2_ASAP7_75t_L g2910 ( 
.A1(n_2885),
.A2(n_2750),
.A3(n_2646),
.B(n_2665),
.Y(n_2910)
);

CKINVDCx12_ASAP7_75t_R g2911 ( 
.A(n_2900),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2813),
.Y(n_2912)
);

NAND2x1p5_ASAP7_75t_L g2913 ( 
.A(n_2846),
.B(n_2801),
.Y(n_2913)
);

OAI21x1_ASAP7_75t_L g2914 ( 
.A1(n_2858),
.A2(n_2644),
.B(n_2809),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2837),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2812),
.Y(n_2916)
);

CKINVDCx6p67_ASAP7_75t_R g2917 ( 
.A(n_2820),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2849),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2850),
.Y(n_2919)
);

AOI22xp33_ASAP7_75t_L g2920 ( 
.A1(n_2876),
.A2(n_2798),
.B1(n_2802),
.B2(n_2800),
.Y(n_2920)
);

OAI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2889),
.A2(n_2795),
.B1(n_2789),
.B2(n_2788),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2864),
.B(n_2898),
.Y(n_2922)
);

HB1xp67_ASAP7_75t_L g2923 ( 
.A(n_2873),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2830),
.Y(n_2924)
);

AO31x2_ASAP7_75t_L g2925 ( 
.A1(n_2862),
.A2(n_2896),
.A3(n_2895),
.B(n_2892),
.Y(n_2925)
);

AO21x2_ASAP7_75t_L g2926 ( 
.A1(n_2899),
.A2(n_2808),
.B(n_2736),
.Y(n_2926)
);

CKINVDCx11_ASAP7_75t_R g2927 ( 
.A(n_2854),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2831),
.Y(n_2928)
);

OAI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2891),
.A2(n_2810),
.B(n_2767),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2866),
.A2(n_2761),
.B(n_2804),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2823),
.B(n_1127),
.Y(n_2931)
);

CKINVDCx5p33_ASAP7_75t_R g2932 ( 
.A(n_2818),
.Y(n_2932)
);

OAI21x1_ASAP7_75t_L g2933 ( 
.A1(n_2843),
.A2(n_2769),
.B(n_2764),
.Y(n_2933)
);

OAI21x1_ASAP7_75t_L g2934 ( 
.A1(n_2851),
.A2(n_2763),
.B(n_2773),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2857),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2855),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2841),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2868),
.B(n_1127),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2883),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2870),
.B(n_1496),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2880),
.A2(n_1322),
.B(n_1318),
.Y(n_2941)
);

OAI21x1_ASAP7_75t_L g2942 ( 
.A1(n_2897),
.A2(n_1065),
.B(n_1054),
.Y(n_2942)
);

AOI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2872),
.A2(n_2871),
.B1(n_2878),
.B2(n_2884),
.Y(n_2943)
);

OA21x2_ASAP7_75t_L g2944 ( 
.A1(n_2886),
.A2(n_1225),
.B(n_1160),
.Y(n_2944)
);

BUFx2_ASAP7_75t_L g2945 ( 
.A(n_2869),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2883),
.Y(n_2946)
);

AND2x2_ASAP7_75t_SL g2947 ( 
.A(n_2861),
.B(n_2863),
.Y(n_2947)
);

OA21x2_ASAP7_75t_L g2948 ( 
.A1(n_2829),
.A2(n_1395),
.B(n_1251),
.Y(n_2948)
);

AOI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2879),
.A2(n_1000),
.B1(n_1005),
.B2(n_988),
.Y(n_2949)
);

INVxp67_ASAP7_75t_SL g2950 ( 
.A(n_2848),
.Y(n_2950)
);

OAI21x1_ASAP7_75t_L g2951 ( 
.A1(n_2848),
.A2(n_2822),
.B(n_2819),
.Y(n_2951)
);

AO21x2_ASAP7_75t_L g2952 ( 
.A1(n_2815),
.A2(n_1169),
.B(n_1116),
.Y(n_2952)
);

BUFx2_ASAP7_75t_SL g2953 ( 
.A(n_2828),
.Y(n_2953)
);

OAI21x1_ASAP7_75t_L g2954 ( 
.A1(n_2848),
.A2(n_1265),
.B(n_1231),
.Y(n_2954)
);

INVx2_ASAP7_75t_SL g2955 ( 
.A(n_2817),
.Y(n_2955)
);

OAI21x1_ASAP7_75t_L g2956 ( 
.A1(n_2824),
.A2(n_1368),
.B(n_1269),
.Y(n_2956)
);

OAI21x1_ASAP7_75t_L g2957 ( 
.A1(n_2811),
.A2(n_1430),
.B(n_1379),
.Y(n_2957)
);

INVx6_ASAP7_75t_L g2958 ( 
.A(n_2852),
.Y(n_2958)
);

CKINVDCx6p67_ASAP7_75t_R g2959 ( 
.A(n_2840),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2881),
.Y(n_2960)
);

O2A1O1Ixp5_ASAP7_75t_L g2961 ( 
.A1(n_2842),
.A2(n_1483),
.B(n_1200),
.C(n_1224),
.Y(n_2961)
);

BUFx3_ASAP7_75t_L g2962 ( 
.A(n_2826),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2845),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2853),
.A2(n_1200),
.B(n_1127),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2874),
.A2(n_1374),
.B1(n_1224),
.B2(n_1027),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2814),
.B(n_1327),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2902),
.Y(n_2967)
);

CKINVDCx6p67_ASAP7_75t_R g2968 ( 
.A(n_2927),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2920),
.A2(n_2893),
.B1(n_2874),
.B2(n_2894),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2903),
.Y(n_2970)
);

BUFx3_ASAP7_75t_L g2971 ( 
.A(n_2962),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2935),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2924),
.Y(n_2973)
);

INVx2_ASAP7_75t_SL g2974 ( 
.A(n_2916),
.Y(n_2974)
);

INVx4_ASAP7_75t_L g2975 ( 
.A(n_2959),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2928),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2937),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2936),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2912),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2939),
.B(n_2827),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2958),
.Y(n_2981)
);

BUFx2_ASAP7_75t_L g2982 ( 
.A(n_2950),
.Y(n_2982)
);

AOI22xp33_ASAP7_75t_SL g2983 ( 
.A1(n_2905),
.A2(n_2860),
.B1(n_2877),
.B2(n_2840),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2946),
.B(n_2845),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2923),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2904),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2909),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2958),
.Y(n_2988)
);

NOR2x1_ASAP7_75t_SL g2989 ( 
.A(n_2901),
.B(n_2926),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2918),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2919),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2922),
.Y(n_2992)
);

INVx2_ASAP7_75t_SL g2993 ( 
.A(n_2963),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2925),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2925),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2915),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2951),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2953),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2938),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2947),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2911),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2964),
.Y(n_3002)
);

BUFx2_ASAP7_75t_SL g3003 ( 
.A(n_2960),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2908),
.Y(n_3004)
);

BUFx2_ASAP7_75t_L g3005 ( 
.A(n_2948),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_2932),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2931),
.B(n_2952),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2944),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2943),
.B(n_2821),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2942),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2929),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2906),
.Y(n_3012)
);

OAI21x1_ASAP7_75t_L g3013 ( 
.A1(n_2954),
.A2(n_1374),
.B(n_1224),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2956),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2914),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2957),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2921),
.A2(n_2865),
.B1(n_1374),
.B2(n_1224),
.Y(n_3017)
);

CKINVDCx16_ASAP7_75t_R g3018 ( 
.A(n_2971),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2967),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_R g3020 ( 
.A(n_2968),
.B(n_2917),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2985),
.B(n_2945),
.Y(n_3021)
);

AO21x2_ASAP7_75t_L g3022 ( 
.A1(n_2989),
.A2(n_2941),
.B(n_2930),
.Y(n_3022)
);

NAND2xp33_ASAP7_75t_R g3023 ( 
.A(n_2981),
.B(n_2940),
.Y(n_3023)
);

AOI21xp33_ASAP7_75t_L g3024 ( 
.A1(n_3007),
.A2(n_2961),
.B(n_2965),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2986),
.B(n_2955),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2982),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2999),
.A2(n_1374),
.B1(n_2934),
.B2(n_2933),
.Y(n_3027)
);

OR2x2_ASAP7_75t_L g3028 ( 
.A(n_2970),
.B(n_2966),
.Y(n_3028)
);

AND2x6_ASAP7_75t_L g3029 ( 
.A(n_3000),
.B(n_2847),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2987),
.B(n_2913),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_3001),
.B(n_2833),
.Y(n_3031)
);

CKINVDCx20_ASAP7_75t_R g3032 ( 
.A(n_3006),
.Y(n_3032)
);

INVx3_ASAP7_75t_L g3033 ( 
.A(n_2996),
.Y(n_3033)
);

NAND2xp33_ASAP7_75t_R g3034 ( 
.A(n_2988),
.B(n_3009),
.Y(n_3034)
);

CKINVDCx11_ASAP7_75t_R g3035 ( 
.A(n_2998),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2980),
.B(n_2825),
.Y(n_3036)
);

CKINVDCx16_ASAP7_75t_R g3037 ( 
.A(n_2975),
.Y(n_3037)
);

NAND2xp33_ASAP7_75t_R g3038 ( 
.A(n_2984),
.B(n_0),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2983),
.A2(n_2835),
.B1(n_2949),
.B2(n_2844),
.Y(n_3039)
);

CKINVDCx16_ASAP7_75t_R g3040 ( 
.A(n_2975),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_R g3041 ( 
.A(n_2974),
.B(n_2832),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2989),
.A2(n_2907),
.B(n_2839),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2972),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_3003),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2982),
.B(n_2816),
.Y(n_3045)
);

AO31x2_ASAP7_75t_L g3046 ( 
.A1(n_2995),
.A2(n_2907),
.A3(n_2910),
.B(n_1374),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_3004),
.B(n_1374),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2977),
.B(n_2834),
.Y(n_3048)
);

NAND2xp33_ASAP7_75t_R g3049 ( 
.A(n_2992),
.B(n_2),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2990),
.B(n_1012),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2973),
.B(n_1028),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2978),
.B(n_2910),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2993),
.Y(n_3053)
);

INVxp67_ASAP7_75t_L g3054 ( 
.A(n_2991),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2976),
.B(n_1034),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2979),
.Y(n_3056)
);

NAND2xp33_ASAP7_75t_R g3057 ( 
.A(n_3005),
.B(n_2997),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2994),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3005),
.Y(n_3059)
);

OR2x6_ASAP7_75t_L g3060 ( 
.A(n_3008),
.B(n_3014),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_3011),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_3012),
.B(n_2),
.Y(n_3062)
);

INVx4_ASAP7_75t_L g3063 ( 
.A(n_3016),
.Y(n_3063)
);

INVx2_ASAP7_75t_SL g3064 ( 
.A(n_3002),
.Y(n_3064)
);

NAND2xp33_ASAP7_75t_R g3065 ( 
.A(n_3010),
.B(n_3),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_3015),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_3019),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_3033),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_3032),
.Y(n_3069)
);

AND2x4_ASAP7_75t_L g3070 ( 
.A(n_3026),
.B(n_3013),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_3059),
.B(n_2969),
.Y(n_3071)
);

AO21x2_ASAP7_75t_L g3072 ( 
.A1(n_3042),
.A2(n_3017),
.B(n_4),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_3043),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_3056),
.Y(n_3074)
);

NOR2x1_ASAP7_75t_L g3075 ( 
.A(n_3047),
.B(n_5),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_3025),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_3054),
.B(n_1035),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_3058),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_3024),
.A2(n_1478),
.B1(n_1490),
.B2(n_1477),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_3018),
.B(n_5),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_3021),
.B(n_6),
.Y(n_3081)
);

OR2x2_ASAP7_75t_L g3082 ( 
.A(n_3052),
.B(n_7),
.Y(n_3082)
);

AND2x4_ASAP7_75t_L g3083 ( 
.A(n_3060),
.B(n_8),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_3030),
.B(n_9),
.Y(n_3084)
);

OR2x2_ASAP7_75t_L g3085 ( 
.A(n_3060),
.B(n_10),
.Y(n_3085)
);

NAND2x1p5_ASAP7_75t_L g3086 ( 
.A(n_3045),
.B(n_536),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_3063),
.B(n_3064),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_3061),
.Y(n_3088)
);

INVx2_ASAP7_75t_SL g3089 ( 
.A(n_3053),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_3066),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3037),
.B(n_12),
.Y(n_3091)
);

OR2x2_ASAP7_75t_L g3092 ( 
.A(n_3028),
.B(n_13),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3062),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_3040),
.B(n_13),
.Y(n_3094)
);

INVxp67_ASAP7_75t_SL g3095 ( 
.A(n_3057),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_3048),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_3069),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_3095),
.B(n_3044),
.Y(n_3098)
);

INVx3_ASAP7_75t_SL g3099 ( 
.A(n_3083),
.Y(n_3099)
);

OA21x2_ASAP7_75t_L g3100 ( 
.A1(n_3078),
.A2(n_3027),
.B(n_3051),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_3068),
.B(n_3036),
.Y(n_3101)
);

INVxp67_ASAP7_75t_SL g3102 ( 
.A(n_3085),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_3073),
.Y(n_3103)
);

OA21x2_ASAP7_75t_L g3104 ( 
.A1(n_3067),
.A2(n_3055),
.B(n_3031),
.Y(n_3104)
);

INVx2_ASAP7_75t_SL g3105 ( 
.A(n_3089),
.Y(n_3105)
);

OAI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_3079),
.A2(n_3050),
.B(n_3039),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_3074),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3093),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_3096),
.B(n_3035),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_3090),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_3082),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3088),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_3087),
.Y(n_3113)
);

AOI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_3072),
.A2(n_3022),
.B(n_3065),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3087),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_3070),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_3070),
.Y(n_3117)
);

OAI221xp5_ASAP7_75t_L g3118 ( 
.A1(n_3075),
.A2(n_3049),
.B1(n_3023),
.B2(n_3034),
.C(n_3038),
.Y(n_3118)
);

OAI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_3092),
.A2(n_3029),
.B1(n_3041),
.B2(n_3020),
.Y(n_3119)
);

OAI22xp33_ASAP7_75t_L g3120 ( 
.A1(n_3086),
.A2(n_3029),
.B1(n_1042),
.B2(n_1044),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_3071),
.B(n_3076),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3071),
.Y(n_3122)
);

INVx5_ASAP7_75t_L g3123 ( 
.A(n_3080),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_3091),
.A2(n_3029),
.B1(n_1047),
.B2(n_1048),
.Y(n_3124)
);

INVx5_ASAP7_75t_L g3125 ( 
.A(n_3094),
.Y(n_3125)
);

OAI221xp5_ASAP7_75t_L g3126 ( 
.A1(n_3118),
.A2(n_3077),
.B1(n_3084),
.B2(n_3081),
.C(n_1050),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3104),
.B(n_3083),
.Y(n_3127)
);

OAI21xp33_ASAP7_75t_L g3128 ( 
.A1(n_3114),
.A2(n_1049),
.B(n_1040),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3102),
.B(n_3046),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_3122),
.B(n_3113),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_3108),
.B(n_3046),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3110),
.Y(n_3132)
);

AOI222xp33_ASAP7_75t_L g3133 ( 
.A1(n_3106),
.A2(n_1055),
.B1(n_1052),
.B2(n_1058),
.C1(n_1053),
.C2(n_1051),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_3098),
.B(n_14),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3103),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3107),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_3115),
.B(n_15),
.Y(n_3137)
);

AND2x2_ASAP7_75t_L g3138 ( 
.A(n_3116),
.B(n_15),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_3117),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3111),
.Y(n_3140)
);

INVx3_ASAP7_75t_L g3141 ( 
.A(n_3123),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_3121),
.Y(n_3142)
);

INVxp67_ASAP7_75t_SL g3143 ( 
.A(n_3119),
.Y(n_3143)
);

INVxp67_ASAP7_75t_L g3144 ( 
.A(n_3112),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_3125),
.B(n_1068),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3125),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3123),
.B(n_16),
.Y(n_3147)
);

BUFx3_ASAP7_75t_L g3148 ( 
.A(n_3097),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3123),
.Y(n_3149)
);

OAI21xp5_ASAP7_75t_SL g3150 ( 
.A1(n_3124),
.A2(n_17),
.B(n_18),
.Y(n_3150)
);

NAND4xp25_ASAP7_75t_SL g3151 ( 
.A(n_3109),
.B(n_20),
.C(n_18),
.D(n_19),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_3100),
.A2(n_1079),
.B1(n_1082),
.B2(n_1077),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_3099),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3101),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_3105),
.B(n_1083),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_3153),
.B(n_20),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_3152),
.B(n_3120),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_3130),
.B(n_21),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_3141),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_3154),
.B(n_21),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_3149),
.B(n_22),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_3141),
.B(n_25),
.Y(n_3162)
);

OAI31xp33_ASAP7_75t_L g3163 ( 
.A1(n_3128),
.A2(n_27),
.A3(n_25),
.B(n_26),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3142),
.B(n_27),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_3140),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3132),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3146),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3135),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_3143),
.B(n_1084),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3136),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3139),
.B(n_28),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_3144),
.B(n_28),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_3148),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3127),
.B(n_3137),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3138),
.B(n_30),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_3134),
.B(n_31),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3147),
.B(n_31),
.Y(n_3177)
);

AND2x4_ASAP7_75t_L g3178 ( 
.A(n_3129),
.B(n_32),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3131),
.B(n_33),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3145),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3155),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_3126),
.Y(n_3182)
);

OR2x2_ASAP7_75t_L g3183 ( 
.A(n_3151),
.B(n_33),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3133),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_3150),
.B(n_34),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_3173),
.B(n_35),
.Y(n_3186)
);

INVxp67_ASAP7_75t_L g3187 ( 
.A(n_3159),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3168),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_3174),
.B(n_36),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3168),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3180),
.B(n_37),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3170),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_3181),
.B(n_38),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3178),
.B(n_3179),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_3178),
.B(n_38),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_3162),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3156),
.B(n_41),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_3167),
.B(n_3166),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3160),
.B(n_42),
.Y(n_3199)
);

INVxp67_ASAP7_75t_L g3200 ( 
.A(n_3169),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3184),
.B(n_1095),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3165),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3182),
.B(n_1097),
.Y(n_3203)
);

AND2x2_ASAP7_75t_L g3204 ( 
.A(n_3158),
.B(n_42),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3161),
.Y(n_3205)
);

INVxp67_ASAP7_75t_SL g3206 ( 
.A(n_3157),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_3164),
.Y(n_3207)
);

OR2x2_ASAP7_75t_L g3208 ( 
.A(n_3172),
.B(n_43),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3171),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3176),
.B(n_43),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3177),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3175),
.Y(n_3212)
);

INVxp67_ASAP7_75t_SL g3213 ( 
.A(n_3183),
.Y(n_3213)
);

INVx3_ASAP7_75t_R g3214 ( 
.A(n_3185),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3163),
.Y(n_3215)
);

AND2x4_ASAP7_75t_L g3216 ( 
.A(n_3159),
.B(n_44),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3173),
.B(n_44),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3178),
.B(n_1098),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3168),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3173),
.B(n_45),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_3159),
.B(n_46),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3188),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3190),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3192),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_3196),
.B(n_47),
.Y(n_3225)
);

HB1xp67_ASAP7_75t_L g3226 ( 
.A(n_3187),
.Y(n_3226)
);

INVx2_ASAP7_75t_SL g3227 ( 
.A(n_3221),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_3207),
.Y(n_3228)
);

INVx2_ASAP7_75t_SL g3229 ( 
.A(n_3221),
.Y(n_3229)
);

INVx5_ASAP7_75t_L g3230 ( 
.A(n_3186),
.Y(n_3230)
);

NAND4xp25_ASAP7_75t_L g3231 ( 
.A(n_3215),
.B(n_1106),
.C(n_1107),
.D(n_1101),
.Y(n_3231)
);

NAND2xp33_ASAP7_75t_R g3232 ( 
.A(n_3189),
.B(n_47),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3206),
.B(n_1108),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3205),
.B(n_1114),
.Y(n_3234)
);

HB1xp67_ASAP7_75t_L g3235 ( 
.A(n_3194),
.Y(n_3235)
);

AO21x2_ASAP7_75t_L g3236 ( 
.A1(n_3201),
.A2(n_48),
.B(n_49),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3212),
.B(n_1120),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3211),
.B(n_1122),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3219),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3198),
.Y(n_3240)
);

CKINVDCx16_ASAP7_75t_R g3241 ( 
.A(n_3197),
.Y(n_3241)
);

NOR2xp33_ASAP7_75t_L g3242 ( 
.A(n_3214),
.B(n_1137),
.Y(n_3242)
);

INVx1_ASAP7_75t_SL g3243 ( 
.A(n_3195),
.Y(n_3243)
);

AND2x4_ASAP7_75t_L g3244 ( 
.A(n_3209),
.B(n_49),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3202),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_3200),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3193),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3217),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3191),
.Y(n_3249)
);

NOR2xp67_ASAP7_75t_L g3250 ( 
.A(n_3208),
.B(n_50),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_3204),
.B(n_50),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_3220),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3210),
.Y(n_3253)
);

OR2x2_ASAP7_75t_L g3254 ( 
.A(n_3203),
.B(n_52),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3199),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3218),
.Y(n_3256)
);

INVx1_ASAP7_75t_SL g3257 ( 
.A(n_3195),
.Y(n_3257)
);

NOR2x1_ASAP7_75t_L g3258 ( 
.A(n_3216),
.B(n_54),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3213),
.B(n_1144),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3188),
.Y(n_3260)
);

AOI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_3206),
.A2(n_1150),
.B1(n_1153),
.B2(n_1149),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3216),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_3216),
.Y(n_3263)
);

AOI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_3215),
.A2(n_1471),
.B1(n_1491),
.B2(n_1467),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3216),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3213),
.B(n_1154),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3196),
.B(n_55),
.Y(n_3267)
);

OAI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3215),
.A2(n_1165),
.B1(n_1194),
.B2(n_1184),
.Y(n_3268)
);

INVx1_ASAP7_75t_SL g3269 ( 
.A(n_3195),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3188),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3241),
.B(n_1163),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3228),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3226),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3243),
.B(n_56),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3246),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_3255),
.A2(n_3252),
.B1(n_3253),
.B2(n_3248),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_3230),
.B(n_1176),
.Y(n_3277)
);

INVxp67_ASAP7_75t_L g3278 ( 
.A(n_3232),
.Y(n_3278)
);

OR2x2_ASAP7_75t_L g3279 ( 
.A(n_3257),
.B(n_56),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3227),
.B(n_1181),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3269),
.B(n_57),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3225),
.Y(n_3282)
);

HB1xp67_ASAP7_75t_L g3283 ( 
.A(n_3250),
.Y(n_3283)
);

INVx2_ASAP7_75t_SL g3284 ( 
.A(n_3263),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3263),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3229),
.B(n_1188),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3262),
.B(n_1189),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3267),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3265),
.B(n_1191),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3258),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3235),
.B(n_1193),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3247),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3249),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3242),
.B(n_1195),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3240),
.Y(n_3295)
);

HB1xp67_ASAP7_75t_L g3296 ( 
.A(n_3236),
.Y(n_3296)
);

INVx2_ASAP7_75t_SL g3297 ( 
.A(n_3244),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_R g3298 ( 
.A(n_3264),
.B(n_58),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3222),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3223),
.Y(n_3300)
);

HB1xp67_ASAP7_75t_L g3301 ( 
.A(n_3224),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3256),
.A2(n_3261),
.B1(n_3268),
.B2(n_3233),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3239),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3260),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_3231),
.B(n_1198),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3251),
.B(n_1201),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3270),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3254),
.B(n_1211),
.Y(n_3308)
);

OR2x2_ASAP7_75t_L g3309 ( 
.A(n_3259),
.B(n_59),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3234),
.B(n_3245),
.Y(n_3310)
);

NAND3xp33_ASAP7_75t_L g3311 ( 
.A(n_3266),
.B(n_1218),
.C(n_1215),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3237),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3238),
.Y(n_3313)
);

INVxp67_ASAP7_75t_L g3314 ( 
.A(n_3232),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3228),
.Y(n_3315)
);

INVx1_ASAP7_75t_SL g3316 ( 
.A(n_3230),
.Y(n_3316)
);

INVx1_ASAP7_75t_SL g3317 ( 
.A(n_3230),
.Y(n_3317)
);

HB1xp67_ASAP7_75t_L g3318 ( 
.A(n_3230),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3241),
.B(n_1220),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_3241),
.B(n_1222),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3241),
.B(n_1227),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_3241),
.B(n_60),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3228),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3228),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3263),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3263),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3241),
.B(n_1229),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3228),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3241),
.B(n_1234),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3241),
.B(n_1238),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3228),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_3227),
.B(n_62),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3228),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3228),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3318),
.Y(n_3335)
);

AOI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3314),
.A2(n_1253),
.B1(n_1255),
.B2(n_1246),
.Y(n_3336)
);

OR2x2_ASAP7_75t_L g3337 ( 
.A(n_3290),
.B(n_3283),
.Y(n_3337)
);

OAI22xp33_ASAP7_75t_SL g3338 ( 
.A1(n_3317),
.A2(n_1497),
.B1(n_1500),
.B2(n_1494),
.Y(n_3338)
);

OAI21xp33_ASAP7_75t_L g3339 ( 
.A1(n_3276),
.A2(n_1272),
.B(n_1271),
.Y(n_3339)
);

AOI221x1_ASAP7_75t_L g3340 ( 
.A1(n_3273),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3332),
.Y(n_3341)
);

AND2x4_ASAP7_75t_L g3342 ( 
.A(n_3284),
.B(n_63),
.Y(n_3342)
);

O2A1O1Ixp33_ASAP7_75t_L g3343 ( 
.A1(n_3275),
.A2(n_67),
.B(n_64),
.C(n_65),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_3272),
.B(n_1452),
.C(n_1449),
.Y(n_3344)
);

AOI32xp33_ASAP7_75t_L g3345 ( 
.A1(n_3285),
.A2(n_1280),
.A3(n_1281),
.B1(n_1276),
.B2(n_1274),
.Y(n_3345)
);

AOI211xp5_ASAP7_75t_L g3346 ( 
.A1(n_3315),
.A2(n_1286),
.B(n_1288),
.C(n_1285),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3332),
.Y(n_3347)
);

OR2x2_ASAP7_75t_L g3348 ( 
.A(n_3322),
.B(n_3328),
.Y(n_3348)
);

AOI221xp5_ASAP7_75t_L g3349 ( 
.A1(n_3323),
.A2(n_1307),
.B1(n_1311),
.B2(n_1305),
.C(n_1303),
.Y(n_3349)
);

OAI21xp33_ASAP7_75t_SL g3350 ( 
.A1(n_3324),
.A2(n_67),
.B(n_68),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3325),
.B(n_1313),
.Y(n_3351)
);

INVx2_ASAP7_75t_SL g3352 ( 
.A(n_3331),
.Y(n_3352)
);

O2A1O1Ixp33_ASAP7_75t_L g3353 ( 
.A1(n_3333),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3353)
);

INVxp67_ASAP7_75t_SL g3354 ( 
.A(n_3277),
.Y(n_3354)
);

OAI21xp33_ASAP7_75t_L g3355 ( 
.A1(n_3326),
.A2(n_1326),
.B(n_1325),
.Y(n_3355)
);

XOR2x2_ASAP7_75t_L g3356 ( 
.A(n_3297),
.B(n_70),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3334),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3274),
.Y(n_3358)
);

OR2x2_ASAP7_75t_L g3359 ( 
.A(n_3282),
.B(n_72),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3288),
.B(n_1328),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3271),
.B(n_1329),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3279),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3319),
.B(n_1330),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3281),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_SL g3365 ( 
.A1(n_3302),
.A2(n_73),
.B(n_74),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3320),
.B(n_1332),
.Y(n_3366)
);

HB1xp67_ASAP7_75t_L g3367 ( 
.A(n_3301),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3321),
.B(n_1348),
.Y(n_3368)
);

OR2x2_ASAP7_75t_L g3369 ( 
.A(n_3327),
.B(n_75),
.Y(n_3369)
);

AOI221x1_ASAP7_75t_L g3370 ( 
.A1(n_3329),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_3330),
.B(n_3309),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3313),
.A2(n_3312),
.B1(n_3293),
.B2(n_3292),
.Y(n_3372)
);

OAI21xp33_ASAP7_75t_L g3373 ( 
.A1(n_3295),
.A2(n_1353),
.B(n_1352),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_3287),
.B(n_76),
.Y(n_3374)
);

OAI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3280),
.A2(n_3286),
.B1(n_3307),
.B2(n_3311),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3306),
.B(n_1360),
.Y(n_3376)
);

OAI31xp33_ASAP7_75t_L g3377 ( 
.A1(n_3291),
.A2(n_80),
.A3(n_77),
.B(n_78),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3289),
.A2(n_1367),
.B1(n_1370),
.B2(n_1366),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3308),
.B(n_1375),
.Y(n_3379)
);

OAI21xp5_ASAP7_75t_SL g3380 ( 
.A1(n_3310),
.A2(n_81),
.B(n_82),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3299),
.Y(n_3381)
);

INVxp67_ASAP7_75t_L g3382 ( 
.A(n_3305),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_3294),
.B(n_1376),
.Y(n_3383)
);

NAND3xp33_ASAP7_75t_L g3384 ( 
.A(n_3300),
.B(n_1460),
.C(n_1456),
.Y(n_3384)
);

OR2x2_ASAP7_75t_L g3385 ( 
.A(n_3303),
.B(n_81),
.Y(n_3385)
);

XNOR2x1_ASAP7_75t_L g3386 ( 
.A(n_3304),
.B(n_83),
.Y(n_3386)
);

AOI21xp33_ASAP7_75t_L g3387 ( 
.A1(n_3298),
.A2(n_1397),
.B(n_1396),
.Y(n_3387)
);

INVx3_ASAP7_75t_L g3388 ( 
.A(n_3332),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3278),
.B(n_1403),
.Y(n_3389)
);

AND2x4_ASAP7_75t_L g3390 ( 
.A(n_3318),
.B(n_84),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3318),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_L g3392 ( 
.A(n_3278),
.B(n_1411),
.Y(n_3392)
);

OAI21xp5_ASAP7_75t_SL g3393 ( 
.A1(n_3278),
.A2(n_86),
.B(n_87),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3318),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3318),
.Y(n_3395)
);

OAI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3278),
.A2(n_1443),
.B(n_1439),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3318),
.Y(n_3397)
);

OAI21xp33_ASAP7_75t_L g3398 ( 
.A1(n_3278),
.A2(n_1445),
.B(n_1444),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3318),
.Y(n_3399)
);

NAND2x1p5_ASAP7_75t_L g3400 ( 
.A(n_3316),
.B(n_89),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3278),
.A2(n_1466),
.B(n_1463),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3318),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3278),
.B(n_1506),
.Y(n_3403)
);

AOI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_3278),
.A2(n_1510),
.B1(n_1511),
.B2(n_1447),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3318),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3278),
.B(n_90),
.Y(n_3406)
);

NAND2x1p5_ASAP7_75t_L g3407 ( 
.A(n_3316),
.B(n_91),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3278),
.B(n_91),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_3322),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3318),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3318),
.Y(n_3411)
);

OR2x2_ASAP7_75t_L g3412 ( 
.A(n_3278),
.B(n_92),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3278),
.B(n_94),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_SL g3414 ( 
.A(n_3278),
.B(n_1339),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3318),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3278),
.A2(n_1458),
.B1(n_1421),
.B2(n_1341),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3278),
.B(n_94),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3278),
.B(n_97),
.Y(n_3418)
);

OAI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3296),
.A2(n_1344),
.B1(n_1351),
.B2(n_1340),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3318),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3278),
.A2(n_1377),
.B1(n_1386),
.B2(n_1357),
.Y(n_3421)
);

NOR2xp67_ASAP7_75t_L g3422 ( 
.A(n_3318),
.B(n_100),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3318),
.Y(n_3423)
);

OR2x2_ASAP7_75t_L g3424 ( 
.A(n_3278),
.B(n_99),
.Y(n_3424)
);

NOR4xp25_ASAP7_75t_L g3425 ( 
.A(n_3316),
.B(n_103),
.C(n_101),
.D(n_102),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_3278),
.B(n_102),
.Y(n_3426)
);

AOI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3278),
.A2(n_1455),
.B1(n_1415),
.B2(n_1388),
.Y(n_3427)
);

OAI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3278),
.A2(n_1389),
.B1(n_1392),
.B2(n_1387),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_3278),
.A2(n_1413),
.B(n_1412),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3278),
.B(n_104),
.Y(n_3430)
);

AOI221xp5_ASAP7_75t_L g3431 ( 
.A1(n_3278),
.A2(n_1479),
.B1(n_1480),
.B2(n_1469),
.C(n_1446),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3278),
.B(n_104),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3278),
.A2(n_1422),
.B1(n_1423),
.B2(n_1416),
.Y(n_3433)
);

OAI21xp33_ASAP7_75t_L g3434 ( 
.A1(n_3278),
.A2(n_1436),
.B(n_1434),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3318),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3318),
.Y(n_3436)
);

OAI322xp33_ASAP7_75t_L g3437 ( 
.A1(n_3278),
.A2(n_111),
.A3(n_110),
.B1(n_108),
.B2(n_106),
.C1(n_107),
.C2(n_109),
.Y(n_3437)
);

NOR3xp33_ASAP7_75t_L g3438 ( 
.A(n_3278),
.B(n_1441),
.C(n_106),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3318),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3318),
.Y(n_3440)
);

OAI21xp33_ASAP7_75t_SL g3441 ( 
.A1(n_3296),
.A2(n_109),
.B(n_110),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3318),
.Y(n_3442)
);

OAI21xp33_ASAP7_75t_SL g3443 ( 
.A1(n_3296),
.A2(n_112),
.B(n_113),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3388),
.B(n_113),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3341),
.B(n_115),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3422),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3425),
.B(n_115),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3400),
.Y(n_3448)
);

NOR2x1_ASAP7_75t_L g3449 ( 
.A(n_3337),
.B(n_116),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3347),
.B(n_116),
.Y(n_3450)
);

OR2x2_ASAP7_75t_L g3451 ( 
.A(n_3409),
.B(n_117),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3407),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3367),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3335),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3348),
.B(n_120),
.Y(n_3455)
);

INVxp67_ASAP7_75t_L g3456 ( 
.A(n_3426),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3342),
.B(n_121),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3411),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_SL g3459 ( 
.A1(n_3340),
.A2(n_123),
.B(n_124),
.Y(n_3459)
);

OR2x2_ASAP7_75t_L g3460 ( 
.A(n_3440),
.B(n_123),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3342),
.B(n_126),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3391),
.B(n_127),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3358),
.B(n_3362),
.Y(n_3463)
);

INVx1_ASAP7_75t_SL g3464 ( 
.A(n_3356),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3394),
.Y(n_3465)
);

INVxp67_ASAP7_75t_L g3466 ( 
.A(n_3395),
.Y(n_3466)
);

OR2x2_ASAP7_75t_L g3467 ( 
.A(n_3412),
.B(n_128),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3397),
.B(n_3399),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3402),
.Y(n_3469)
);

INVxp67_ASAP7_75t_L g3470 ( 
.A(n_3405),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3410),
.B(n_128),
.Y(n_3471)
);

AOI211xp5_ASAP7_75t_L g3472 ( 
.A1(n_3441),
.A2(n_139),
.B(n_149),
.C(n_129),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3350),
.B(n_129),
.Y(n_3473)
);

OR2x2_ASAP7_75t_L g3474 ( 
.A(n_3424),
.B(n_130),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3415),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_3364),
.B(n_131),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3420),
.B(n_134),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3354),
.B(n_135),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3352),
.B(n_136),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3423),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3435),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3436),
.Y(n_3482)
);

O2A1O1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_3443),
.A2(n_143),
.B(n_139),
.C(n_140),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3439),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3338),
.B(n_145),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3442),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3390),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3406),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3408),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3413),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3361),
.B(n_147),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3417),
.Y(n_3492)
);

INVxp67_ASAP7_75t_L g3493 ( 
.A(n_3418),
.Y(n_3493)
);

INVxp67_ASAP7_75t_L g3494 ( 
.A(n_3430),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3357),
.B(n_148),
.Y(n_3495)
);

OA21x2_ASAP7_75t_SL g3496 ( 
.A1(n_3414),
.A2(n_148),
.B(n_152),
.Y(n_3496)
);

NOR2x1_ASAP7_75t_L g3497 ( 
.A(n_3393),
.B(n_152),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3432),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_3386),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3382),
.B(n_156),
.Y(n_3500)
);

INVx1_ASAP7_75t_SL g3501 ( 
.A(n_3359),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3380),
.B(n_156),
.Y(n_3502)
);

OR2x2_ASAP7_75t_L g3503 ( 
.A(n_3365),
.B(n_159),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3385),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3371),
.B(n_159),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3369),
.Y(n_3506)
);

XNOR2x2_ASAP7_75t_L g3507 ( 
.A(n_3344),
.B(n_3368),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3351),
.B(n_160),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3374),
.Y(n_3509)
);

OAI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3353),
.A2(n_164),
.B(n_162),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3360),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3381),
.Y(n_3512)
);

OAI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3370),
.A2(n_165),
.B1(n_161),
.B2(n_162),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3389),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3372),
.B(n_166),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3377),
.B(n_167),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3392),
.B(n_167),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3403),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3383),
.B(n_168),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3375),
.B(n_168),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3379),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3438),
.B(n_169),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3345),
.B(n_170),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3376),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3343),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3363),
.Y(n_3526)
);

INVxp67_ASAP7_75t_L g3527 ( 
.A(n_3366),
.Y(n_3527)
);

OAI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3336),
.A2(n_174),
.B(n_172),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3437),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3384),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3446),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3487),
.B(n_3398),
.Y(n_3532)
);

AOI32xp33_ASAP7_75t_L g3533 ( 
.A1(n_3529),
.A2(n_3419),
.A3(n_3346),
.B1(n_3339),
.B2(n_3349),
.Y(n_3533)
);

INVxp67_ASAP7_75t_L g3534 ( 
.A(n_3449),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3448),
.B(n_3452),
.Y(n_3535)
);

INVxp67_ASAP7_75t_SL g3536 ( 
.A(n_3473),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3463),
.B(n_3499),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3457),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3461),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3478),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3472),
.B(n_3404),
.Y(n_3541)
);

OAI221xp5_ASAP7_75t_L g3542 ( 
.A1(n_3466),
.A2(n_3401),
.B1(n_3396),
.B2(n_3434),
.C(n_3373),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3468),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3447),
.B(n_3355),
.Y(n_3544)
);

INVx1_ASAP7_75t_SL g3545 ( 
.A(n_3451),
.Y(n_3545)
);

HB1xp67_ASAP7_75t_L g3546 ( 
.A(n_3479),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3453),
.B(n_3416),
.Y(n_3547)
);

XNOR2xp5_ASAP7_75t_L g3548 ( 
.A(n_3497),
.B(n_3427),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3513),
.B(n_3429),
.Y(n_3549)
);

AOI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_3525),
.A2(n_3378),
.B1(n_3428),
.B2(n_3421),
.Y(n_3550)
);

OR2x2_ASAP7_75t_L g3551 ( 
.A(n_3454),
.B(n_3433),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3515),
.B(n_3431),
.Y(n_3552)
);

INVx1_ASAP7_75t_SL g3553 ( 
.A(n_3455),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3467),
.Y(n_3554)
);

NOR2x1_ASAP7_75t_L g3555 ( 
.A(n_3459),
.B(n_3387),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3444),
.Y(n_3556)
);

NAND4xp25_ASAP7_75t_L g3557 ( 
.A(n_3496),
.B(n_174),
.C(n_171),
.D(n_172),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3458),
.B(n_177),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3505),
.B(n_177),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3460),
.Y(n_3560)
);

HB1xp67_ASAP7_75t_L g3561 ( 
.A(n_3476),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3445),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3450),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3474),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3501),
.B(n_178),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3465),
.B(n_180),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3469),
.B(n_182),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3495),
.Y(n_3568)
);

OAI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3470),
.A2(n_184),
.B(n_185),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3475),
.B(n_184),
.Y(n_3570)
);

INVxp67_ASAP7_75t_L g3571 ( 
.A(n_3502),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3480),
.B(n_186),
.Y(n_3572)
);

INVx1_ASAP7_75t_SL g3573 ( 
.A(n_3520),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3481),
.B(n_186),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3482),
.B(n_187),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3484),
.B(n_188),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3486),
.B(n_190),
.Y(n_3577)
);

AOI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_3456),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3500),
.B(n_3504),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3462),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3471),
.Y(n_3581)
);

NOR3xp33_ASAP7_75t_SL g3582 ( 
.A(n_3509),
.B(n_195),
.C(n_196),
.Y(n_3582)
);

INVxp33_ASAP7_75t_L g3583 ( 
.A(n_3516),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3506),
.Y(n_3584)
);

NAND3xp33_ASAP7_75t_L g3585 ( 
.A(n_3483),
.B(n_195),
.C(n_197),
.Y(n_3585)
);

OR2x2_ASAP7_75t_L g3586 ( 
.A(n_3477),
.B(n_199),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3511),
.B(n_201),
.Y(n_3587)
);

NAND2x1_ASAP7_75t_L g3588 ( 
.A(n_3512),
.B(n_201),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3493),
.B(n_204),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3507),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3491),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3494),
.B(n_205),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3488),
.B(n_205),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3489),
.B(n_206),
.Y(n_3594)
);

OAI21xp5_ASAP7_75t_SL g3595 ( 
.A1(n_3510),
.A2(n_207),
.B(n_208),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3503),
.B(n_209),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3490),
.B(n_210),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3492),
.B(n_211),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3508),
.Y(n_3599)
);

NOR2x1_ASAP7_75t_L g3600 ( 
.A(n_3485),
.B(n_212),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3498),
.B(n_215),
.Y(n_3601)
);

INVx4_ASAP7_75t_L g3602 ( 
.A(n_3514),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3527),
.B(n_215),
.Y(n_3603)
);

OR2x2_ASAP7_75t_L g3604 ( 
.A(n_3523),
.B(n_216),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3517),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3521),
.B(n_217),
.Y(n_3606)
);

OR2x2_ASAP7_75t_L g3607 ( 
.A(n_3522),
.B(n_3530),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3524),
.B(n_220),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3519),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3526),
.B(n_221),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3518),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3528),
.B(n_222),
.Y(n_3612)
);

XOR2x2_ASAP7_75t_L g3613 ( 
.A(n_3464),
.B(n_225),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3448),
.B(n_225),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3464),
.B(n_226),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3448),
.B(n_226),
.Y(n_3616)
);

AND2x4_ASAP7_75t_L g3617 ( 
.A(n_3446),
.B(n_228),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3446),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3464),
.B(n_229),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3448),
.B(n_232),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3446),
.Y(n_3621)
);

NOR3xp33_ASAP7_75t_L g3622 ( 
.A(n_3446),
.B(n_233),
.C(n_234),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3446),
.Y(n_3623)
);

O2A1O1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3447),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3464),
.B(n_235),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3464),
.B(n_236),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3446),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3446),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3446),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3446),
.Y(n_3630)
);

OR2x2_ASAP7_75t_L g3631 ( 
.A(n_3446),
.B(n_238),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3446),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3464),
.B(n_238),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3448),
.B(n_239),
.Y(n_3634)
);

OAI221xp5_ASAP7_75t_L g3635 ( 
.A1(n_3466),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.C(n_244),
.Y(n_3635)
);

NAND3xp33_ASAP7_75t_L g3636 ( 
.A(n_3534),
.B(n_3590),
.C(n_3535),
.Y(n_3636)
);

AO21x1_ASAP7_75t_L g3637 ( 
.A1(n_3588),
.A2(n_243),
.B(n_245),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3537),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_SL g3639 ( 
.A(n_3546),
.B(n_3536),
.Y(n_3639)
);

OAI21xp33_ASAP7_75t_SL g3640 ( 
.A1(n_3555),
.A2(n_250),
.B(n_251),
.Y(n_3640)
);

NOR2xp67_ASAP7_75t_L g3641 ( 
.A(n_3602),
.B(n_252),
.Y(n_3641)
);

NAND3xp33_ASAP7_75t_SL g3642 ( 
.A(n_3624),
.B(n_255),
.C(n_258),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3634),
.A2(n_259),
.B(n_260),
.Y(n_3643)
);

INVxp67_ASAP7_75t_SL g3644 ( 
.A(n_3600),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3561),
.Y(n_3645)
);

OR2x2_ASAP7_75t_L g3646 ( 
.A(n_3557),
.B(n_261),
.Y(n_3646)
);

INVxp67_ASAP7_75t_L g3647 ( 
.A(n_3615),
.Y(n_3647)
);

NOR3x1_ASAP7_75t_L g3648 ( 
.A(n_3595),
.B(n_262),
.C(n_263),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3549),
.A2(n_264),
.B(n_265),
.Y(n_3649)
);

INVx2_ASAP7_75t_SL g3650 ( 
.A(n_3617),
.Y(n_3650)
);

INVx2_ASAP7_75t_SL g3651 ( 
.A(n_3617),
.Y(n_3651)
);

AOI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3579),
.A2(n_268),
.B(n_270),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3540),
.B(n_272),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_3619),
.B(n_273),
.Y(n_3654)
);

AOI221x1_ASAP7_75t_SL g3655 ( 
.A1(n_3531),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.C(n_282),
.Y(n_3655)
);

NOR2xp67_ASAP7_75t_SL g3656 ( 
.A(n_3602),
.B(n_278),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3631),
.Y(n_3657)
);

OAI21xp33_ASAP7_75t_L g3658 ( 
.A1(n_3583),
.A2(n_282),
.B(n_283),
.Y(n_3658)
);

CKINVDCx6p67_ASAP7_75t_R g3659 ( 
.A(n_3625),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3573),
.B(n_284),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3553),
.B(n_287),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3626),
.Y(n_3662)
);

OAI21xp33_ASAP7_75t_L g3663 ( 
.A1(n_3613),
.A2(n_3544),
.B(n_3532),
.Y(n_3663)
);

AOI221xp5_ASAP7_75t_L g3664 ( 
.A1(n_3543),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_3664)
);

NAND3xp33_ASAP7_75t_L g3665 ( 
.A(n_3585),
.B(n_292),
.C(n_294),
.Y(n_3665)
);

NAND3xp33_ASAP7_75t_SL g3666 ( 
.A(n_3545),
.B(n_292),
.C(n_294),
.Y(n_3666)
);

CKINVDCx5p33_ASAP7_75t_R g3667 ( 
.A(n_3582),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3621),
.B(n_295),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3618),
.B(n_296),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3623),
.B(n_297),
.Y(n_3670)
);

NAND2x1p5_ASAP7_75t_L g3671 ( 
.A(n_3564),
.B(n_3560),
.Y(n_3671)
);

HB1xp67_ASAP7_75t_L g3672 ( 
.A(n_3614),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3627),
.B(n_298),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3628),
.B(n_299),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3633),
.A2(n_302),
.B(n_303),
.Y(n_3675)
);

NAND4xp25_ASAP7_75t_L g3676 ( 
.A(n_3533),
.B(n_305),
.C(n_303),
.D(n_304),
.Y(n_3676)
);

NOR3xp33_ASAP7_75t_L g3677 ( 
.A(n_3542),
.B(n_304),
.C(n_305),
.Y(n_3677)
);

NAND3xp33_ASAP7_75t_L g3678 ( 
.A(n_3629),
.B(n_306),
.C(n_307),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3616),
.Y(n_3679)
);

NAND3xp33_ASAP7_75t_SL g3680 ( 
.A(n_3622),
.B(n_306),
.C(n_308),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3630),
.B(n_309),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3632),
.B(n_311),
.Y(n_3682)
);

NOR3xp33_ASAP7_75t_L g3683 ( 
.A(n_3571),
.B(n_313),
.C(n_314),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3620),
.B(n_315),
.Y(n_3684)
);

NAND3xp33_ASAP7_75t_L g3685 ( 
.A(n_3584),
.B(n_315),
.C(n_316),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3608),
.B(n_318),
.Y(n_3686)
);

NAND3xp33_ASAP7_75t_SL g3687 ( 
.A(n_3550),
.B(n_321),
.C(n_323),
.Y(n_3687)
);

INVx1_ASAP7_75t_SL g3688 ( 
.A(n_3565),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3568),
.B(n_324),
.Y(n_3689)
);

NOR2x1_ASAP7_75t_L g3690 ( 
.A(n_3559),
.B(n_325),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3554),
.B(n_3596),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3601),
.B(n_325),
.Y(n_3692)
);

NOR3x1_ASAP7_75t_L g3693 ( 
.A(n_3541),
.B(n_328),
.C(n_332),
.Y(n_3693)
);

NOR3xp33_ASAP7_75t_SL g3694 ( 
.A(n_3552),
.B(n_333),
.C(n_335),
.Y(n_3694)
);

NAND3xp33_ASAP7_75t_L g3695 ( 
.A(n_3548),
.B(n_335),
.C(n_336),
.Y(n_3695)
);

OAI321xp33_ASAP7_75t_L g3696 ( 
.A1(n_3636),
.A2(n_3547),
.A3(n_3611),
.B1(n_3539),
.B2(n_3538),
.C(n_3607),
.Y(n_3696)
);

O2A1O1Ixp33_ASAP7_75t_L g3697 ( 
.A1(n_3666),
.A2(n_3566),
.B(n_3570),
.C(n_3567),
.Y(n_3697)
);

OAI211xp5_ASAP7_75t_L g3698 ( 
.A1(n_3640),
.A2(n_3556),
.B(n_3558),
.C(n_3562),
.Y(n_3698)
);

OAI211xp5_ASAP7_75t_SL g3699 ( 
.A1(n_3663),
.A2(n_3563),
.B(n_3581),
.C(n_3580),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3637),
.Y(n_3700)
);

NOR4xp75_ASAP7_75t_L g3701 ( 
.A(n_3691),
.B(n_3650),
.C(n_3651),
.D(n_3642),
.Y(n_3701)
);

OAI211xp5_ASAP7_75t_L g3702 ( 
.A1(n_3644),
.A2(n_3599),
.B(n_3551),
.C(n_3605),
.Y(n_3702)
);

OAI221xp5_ASAP7_75t_L g3703 ( 
.A1(n_3639),
.A2(n_3574),
.B1(n_3576),
.B2(n_3575),
.C(n_3572),
.Y(n_3703)
);

AOI221xp5_ASAP7_75t_L g3704 ( 
.A1(n_3638),
.A2(n_3645),
.B1(n_3649),
.B2(n_3677),
.C(n_3667),
.Y(n_3704)
);

AOI221xp5_ASAP7_75t_L g3705 ( 
.A1(n_3687),
.A2(n_3676),
.B1(n_3655),
.B2(n_3680),
.C(n_3647),
.Y(n_3705)
);

AOI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3659),
.A2(n_3591),
.B1(n_3609),
.B2(n_3612),
.Y(n_3706)
);

AOI21xp33_ASAP7_75t_L g3707 ( 
.A1(n_3672),
.A2(n_3604),
.B(n_3577),
.Y(n_3707)
);

OAI221xp5_ASAP7_75t_L g3708 ( 
.A1(n_3671),
.A2(n_3569),
.B1(n_3594),
.B2(n_3597),
.C(n_3593),
.Y(n_3708)
);

OAI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3646),
.A2(n_3587),
.B1(n_3586),
.B2(n_3589),
.Y(n_3709)
);

AOI222xp33_ASAP7_75t_L g3710 ( 
.A1(n_3688),
.A2(n_3598),
.B1(n_3592),
.B2(n_3635),
.C1(n_3610),
.C2(n_3606),
.Y(n_3710)
);

OAI32xp33_ASAP7_75t_L g3711 ( 
.A1(n_3660),
.A2(n_3603),
.A3(n_3578),
.B1(n_339),
.B2(n_336),
.Y(n_3711)
);

AOI221xp5_ASAP7_75t_L g3712 ( 
.A1(n_3679),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.C(n_341),
.Y(n_3712)
);

INVx1_ASAP7_75t_SL g3713 ( 
.A(n_3684),
.Y(n_3713)
);

A2O1A1Ixp33_ASAP7_75t_L g3714 ( 
.A1(n_3641),
.A2(n_345),
.B(n_342),
.C(n_343),
.Y(n_3714)
);

AOI211xp5_ASAP7_75t_L g3715 ( 
.A1(n_3665),
.A2(n_345),
.B(n_342),
.C(n_343),
.Y(n_3715)
);

OAI311xp33_ASAP7_75t_L g3716 ( 
.A1(n_3657),
.A2(n_348),
.A3(n_346),
.B1(n_347),
.C1(n_349),
.Y(n_3716)
);

AOI221xp5_ASAP7_75t_L g3717 ( 
.A1(n_3662),
.A2(n_350),
.B1(n_346),
.B2(n_347),
.C(n_351),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3656),
.B(n_351),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3661),
.A2(n_352),
.B(n_355),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3690),
.Y(n_3720)
);

NAND2x1_ASAP7_75t_L g3721 ( 
.A(n_3694),
.B(n_357),
.Y(n_3721)
);

AOI221xp5_ASAP7_75t_L g3722 ( 
.A1(n_3652),
.A2(n_363),
.B1(n_357),
.B2(n_359),
.C(n_364),
.Y(n_3722)
);

OAI221xp5_ASAP7_75t_L g3723 ( 
.A1(n_3668),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.C(n_369),
.Y(n_3723)
);

CKINVDCx16_ASAP7_75t_R g3724 ( 
.A(n_3654),
.Y(n_3724)
);

AOI21xp33_ASAP7_75t_L g3725 ( 
.A1(n_3689),
.A2(n_372),
.B(n_374),
.Y(n_3725)
);

OAI21xp33_ASAP7_75t_L g3726 ( 
.A1(n_3653),
.A2(n_378),
.B(n_379),
.Y(n_3726)
);

OAI221xp5_ASAP7_75t_SL g3727 ( 
.A1(n_3658),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.C(n_382),
.Y(n_3727)
);

NAND4xp25_ASAP7_75t_L g3728 ( 
.A(n_3648),
.B(n_3693),
.C(n_3643),
.D(n_3675),
.Y(n_3728)
);

OAI222xp33_ASAP7_75t_L g3729 ( 
.A1(n_3681),
.A2(n_384),
.B1(n_387),
.B2(n_382),
.C1(n_383),
.C2(n_385),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3686),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3692),
.Y(n_3731)
);

O2A1O1Ixp33_ASAP7_75t_L g3732 ( 
.A1(n_3682),
.A2(n_392),
.B(n_389),
.C(n_391),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_SL g3733 ( 
.A1(n_3669),
.A2(n_393),
.B(n_394),
.Y(n_3733)
);

NAND4xp75_ASAP7_75t_L g3734 ( 
.A(n_3670),
.B(n_396),
.C(n_394),
.D(n_395),
.Y(n_3734)
);

AO22x2_ASAP7_75t_L g3735 ( 
.A1(n_3700),
.A2(n_3695),
.B1(n_3685),
.B2(n_3678),
.Y(n_3735)
);

AOI221xp5_ASAP7_75t_L g3736 ( 
.A1(n_3711),
.A2(n_3674),
.B1(n_3673),
.B2(n_3683),
.C(n_3664),
.Y(n_3736)
);

AO22x2_ASAP7_75t_L g3737 ( 
.A1(n_3720),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_3737)
);

AOI21xp33_ASAP7_75t_L g3738 ( 
.A1(n_3721),
.A2(n_397),
.B(n_398),
.Y(n_3738)
);

AOI221xp5_ASAP7_75t_L g3739 ( 
.A1(n_3696),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.C(n_402),
.Y(n_3739)
);

AOI211xp5_ASAP7_75t_L g3740 ( 
.A1(n_3707),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_3740)
);

OAI21xp33_ASAP7_75t_L g3741 ( 
.A1(n_3728),
.A2(n_3713),
.B(n_3704),
.Y(n_3741)
);

AO221x1_ASAP7_75t_L g3742 ( 
.A1(n_3709),
.A2(n_407),
.B1(n_404),
.B2(n_405),
.C(n_408),
.Y(n_3742)
);

NOR3x1_ASAP7_75t_L g3743 ( 
.A(n_3702),
.B(n_404),
.C(n_405),
.Y(n_3743)
);

HB1xp67_ASAP7_75t_L g3744 ( 
.A(n_3734),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3718),
.Y(n_3745)
);

AOI222xp33_ASAP7_75t_L g3746 ( 
.A1(n_3705),
.A2(n_412),
.B1(n_415),
.B2(n_410),
.C1(n_411),
.C2(n_414),
.Y(n_3746)
);

AOI211xp5_ASAP7_75t_SL g3747 ( 
.A1(n_3698),
.A2(n_3708),
.B(n_3703),
.C(n_3733),
.Y(n_3747)
);

AOI211xp5_ASAP7_75t_L g3748 ( 
.A1(n_3699),
.A2(n_421),
.B(n_416),
.C(n_419),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3724),
.B(n_422),
.Y(n_3749)
);

OAI222xp33_ASAP7_75t_L g3750 ( 
.A1(n_3706),
.A2(n_424),
.B1(n_427),
.B2(n_422),
.C1(n_423),
.C2(n_426),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3714),
.B(n_423),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3710),
.B(n_432),
.Y(n_3752)
);

HB1xp67_ASAP7_75t_L g3753 ( 
.A(n_3701),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3749),
.B(n_3742),
.Y(n_3754)
);

AOI221xp5_ASAP7_75t_L g3755 ( 
.A1(n_3739),
.A2(n_3697),
.B1(n_3716),
.B2(n_3731),
.C(n_3730),
.Y(n_3755)
);

OAI21xp33_ASAP7_75t_L g3756 ( 
.A1(n_3741),
.A2(n_3726),
.B(n_3727),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3752),
.B(n_3719),
.Y(n_3757)
);

AND3x1_ASAP7_75t_L g3758 ( 
.A(n_3748),
.B(n_3715),
.C(n_3722),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3753),
.B(n_3725),
.Y(n_3759)
);

AOI221xp5_ASAP7_75t_L g3760 ( 
.A1(n_3738),
.A2(n_3732),
.B1(n_3729),
.B2(n_3723),
.C(n_3712),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3746),
.B(n_3717),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3737),
.Y(n_3762)
);

A2O1A1Ixp33_ASAP7_75t_L g3763 ( 
.A1(n_3747),
.A2(n_440),
.B(n_438),
.C(n_439),
.Y(n_3763)
);

A2O1A1Ixp33_ASAP7_75t_SL g3764 ( 
.A1(n_3745),
.A2(n_443),
.B(n_440),
.C(n_441),
.Y(n_3764)
);

OR3x1_ASAP7_75t_L g3765 ( 
.A(n_3743),
.B(n_444),
.C(n_447),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3762),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3763),
.B(n_3740),
.Y(n_3767)
);

BUFx2_ASAP7_75t_L g3768 ( 
.A(n_3754),
.Y(n_3768)
);

INVx2_ASAP7_75t_SL g3769 ( 
.A(n_3759),
.Y(n_3769)
);

NOR3xp33_ASAP7_75t_SL g3770 ( 
.A(n_3756),
.B(n_3736),
.C(n_3750),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3758),
.B(n_3735),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3765),
.Y(n_3772)
);

AND2x4_ASAP7_75t_L g3773 ( 
.A(n_3757),
.B(n_3744),
.Y(n_3773)
);

BUFx2_ASAP7_75t_L g3774 ( 
.A(n_3772),
.Y(n_3774)
);

CKINVDCx5p33_ASAP7_75t_R g3775 ( 
.A(n_3770),
.Y(n_3775)
);

CKINVDCx5p33_ASAP7_75t_R g3776 ( 
.A(n_3768),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_3771),
.Y(n_3777)
);

CKINVDCx16_ASAP7_75t_R g3778 ( 
.A(n_3773),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_3769),
.Y(n_3779)
);

HB1xp67_ASAP7_75t_L g3780 ( 
.A(n_3766),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3780),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3779),
.Y(n_3782)
);

AO21x2_ASAP7_75t_L g3783 ( 
.A1(n_3778),
.A2(n_3764),
.B(n_3751),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3782),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3783),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3784),
.Y(n_3786)
);

OAI22xp33_ASAP7_75t_L g3787 ( 
.A1(n_3786),
.A2(n_3777),
.B1(n_3775),
.B2(n_3776),
.Y(n_3787)
);

OAI22xp33_ASAP7_75t_L g3788 ( 
.A1(n_3787),
.A2(n_3781),
.B1(n_3761),
.B2(n_3767),
.Y(n_3788)
);

NAND5xp2_ASAP7_75t_L g3789 ( 
.A(n_3788),
.B(n_3755),
.C(n_3774),
.D(n_3785),
.E(n_3760),
.Y(n_3789)
);

AOI222xp33_ASAP7_75t_L g3790 ( 
.A1(n_3789),
.A2(n_450),
.B1(n_452),
.B2(n_447),
.C1(n_449),
.C2(n_451),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3790),
.A2(n_452),
.B1(n_449),
.B2(n_450),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3791),
.A2(n_458),
.B(n_459),
.Y(n_3792)
);

AOI221xp5_ASAP7_75t_L g3793 ( 
.A1(n_3792),
.A2(n_464),
.B1(n_460),
.B2(n_461),
.C(n_465),
.Y(n_3793)
);

AOI211xp5_ASAP7_75t_L g3794 ( 
.A1(n_3793),
.A2(n_468),
.B(n_465),
.C(n_467),
.Y(n_3794)
);


endmodule