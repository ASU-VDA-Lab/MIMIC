module fake_jpeg_3248_n_391 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_391);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_391;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_5),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_46),
.B(n_50),
.Y(n_107)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_51),
.Y(n_136)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx12f_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_12),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_61),
.B(n_88),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_29),
.B(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_0),
.C(n_1),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_80),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_83),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

CKINVDCx6p67_ASAP7_75t_R g138 ( 
.A(n_82),
.Y(n_138)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_11),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_91),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_32),
.B(n_11),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_94),
.B(n_95),
.Y(n_144)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_40),
.B1(n_23),
.B2(n_15),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_153),
.B1(n_86),
.B2(n_63),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_18),
.C(n_33),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_123),
.C(n_103),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_46),
.A2(n_97),
.B1(n_92),
.B2(n_88),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_119),
.B1(n_133),
.B2(n_134),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_39),
.B1(n_26),
.B2(n_41),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_64),
.A2(n_20),
.B1(n_39),
.B2(n_26),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_70),
.B1(n_66),
.B2(n_67),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_18),
.C(n_28),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_18),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_131),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_40),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_39),
.B1(n_26),
.B2(n_35),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_78),
.A2(n_39),
.B1(n_26),
.B2(n_35),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_71),
.A2(n_84),
.B(n_28),
.C(n_22),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_137),
.A2(n_140),
.B(n_141),
.C(n_114),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_89),
.A2(n_41),
.B1(n_35),
.B2(n_36),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_149),
.B1(n_133),
.B2(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_49),
.A2(n_36),
.B1(n_33),
.B2(n_41),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_57),
.A2(n_31),
.B1(n_27),
.B2(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_155),
.B(n_164),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_27),
.B1(n_82),
.B2(n_80),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_158),
.A2(n_172),
.B1(n_162),
.B2(n_169),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_60),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_175),
.Y(n_204)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_181),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_174),
.B1(n_100),
.B2(n_146),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_109),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_5),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_7),
.B1(n_8),
.B2(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_8),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_105),
.A2(n_129),
.B1(n_150),
.B2(n_148),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_150),
.B1(n_148),
.B2(n_138),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_180),
.B1(n_190),
.B2(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_107),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_183),
.Y(n_225)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_103),
.B(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_134),
.A2(n_122),
.B1(n_143),
.B2(n_125),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_193),
.B1(n_151),
.B2(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_192),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_99),
.B(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_125),
.A2(n_132),
.B1(n_145),
.B2(n_117),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_130),
.B(n_188),
.C(n_187),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_116),
.B(n_113),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_179),
.C(n_159),
.Y(n_226)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_114),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_132),
.B1(n_145),
.B2(n_121),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_206),
.B1(n_221),
.B2(n_229),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_121),
.B1(n_151),
.B2(n_152),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_141),
.B(n_114),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_223),
.B(n_224),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_173),
.A2(n_152),
.B1(n_130),
.B2(n_100),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_130),
.B(n_175),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_224),
.A2(n_195),
.B(n_154),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_157),
.B(n_168),
.C(n_167),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_235),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_189),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_238),
.A2(n_240),
.B(n_251),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_186),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_241),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_195),
.B(n_167),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_167),
.B1(n_163),
.B2(n_181),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_214),
.B1(n_205),
.B2(n_206),
.Y(n_256)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_203),
.B(n_165),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_226),
.C(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_183),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_193),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_203),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_265),
.C(n_276),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_214),
.B1(n_213),
.B2(n_211),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_214),
.B1(n_211),
.B2(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_231),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_217),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_207),
.B1(n_220),
.B2(n_200),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_272),
.B1(n_247),
.B2(n_242),
.Y(n_286)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

AO21x2_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_221),
.B(n_200),
.Y(n_270)
);

AO22x1_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_225),
.B1(n_179),
.B2(n_198),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_228),
.B1(n_222),
.B2(n_166),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_228),
.B(n_222),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_244),
.B(n_243),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_202),
.B1(n_218),
.B2(n_209),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_232),
.B(n_225),
.C(n_198),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_239),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_279),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_235),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_283),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_287),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_291),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_257),
.A2(n_254),
.B1(n_232),
.B2(n_238),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_290),
.A2(n_293),
.B1(n_270),
.B2(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_273),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_267),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_248),
.B1(n_245),
.B2(n_241),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_297),
.B(n_258),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_253),
.C(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_276),
.C(n_278),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_266),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

NAND2x1_ASAP7_75t_SL g297 ( 
.A(n_270),
.B(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_265),
.B(n_227),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_302),
.B(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_261),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_317),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_309),
.B(n_271),
.Y(n_328)
);

NOR4xp25_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_261),
.C(n_266),
.D(n_275),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_321),
.B(n_294),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_315),
.C(n_318),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_260),
.C(n_264),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_270),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_264),
.C(n_278),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_293),
.B1(n_280),
.B2(n_283),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_268),
.B(n_259),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_290),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_332),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_325),
.A2(n_297),
.B(n_298),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_310),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_327),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_304),
.B1(n_305),
.B2(n_303),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_301),
.B(n_281),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_296),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_335),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_285),
.C(n_282),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_318),
.C(n_314),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_259),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_316),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_319),
.B1(n_304),
.B2(n_320),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_338),
.A2(n_306),
.B1(n_286),
.B2(n_303),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_343),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_312),
.B(n_306),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_342),
.A2(n_344),
.B1(n_338),
.B2(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_306),
.C(n_317),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_331),
.B(n_311),
.CI(n_297),
.CON(n_345),
.SN(n_345)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_345),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_347),
.A2(n_350),
.B1(n_329),
.B2(n_323),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_337),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_348),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_353),
.B(n_361),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_355),
.B1(n_358),
.B2(n_359),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_350),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_335),
.B(n_298),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_346),
.A2(n_323),
.B1(n_332),
.B2(n_274),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_336),
.B1(n_256),
.B2(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_343),
.Y(n_363)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_339),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_344),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_362),
.B(n_347),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_345),
.B1(n_309),
.B2(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_358),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_369),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_368),
.A2(n_322),
.B(n_340),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_313),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_341),
.C(n_333),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_371),
.C(n_331),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_340),
.C(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_373),
.A2(n_378),
.B(n_371),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_377),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_345),
.B1(n_300),
.B2(n_271),
.Y(n_377)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_269),
.B(n_161),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_364),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_380),
.A2(n_382),
.B(n_376),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_385),
.B(n_202),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_202),
.C(n_269),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_383),
.B(n_160),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_387),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_388),
.B(n_196),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_182),
.Y(n_391)
);


endmodule