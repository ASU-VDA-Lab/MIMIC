module fake_netlist_1_1718_n_611 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_611);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_611;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_65;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_67;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_446;
wire n_195;
wire n_420;
wire n_165;
wire n_285;
wire n_342;
wire n_423;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_64;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g63 ( .A(n_38), .Y(n_63) );
INVx2_ASAP7_75t_L g64 ( .A(n_27), .Y(n_64) );
CKINVDCx5p33_ASAP7_75t_R g65 ( .A(n_2), .Y(n_65) );
CKINVDCx5p33_ASAP7_75t_R g66 ( .A(n_42), .Y(n_66) );
INVx2_ASAP7_75t_L g67 ( .A(n_55), .Y(n_67) );
NOR2xp67_ASAP7_75t_L g68 ( .A(n_20), .B(n_52), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_2), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_17), .Y(n_70) );
INVxp67_ASAP7_75t_SL g71 ( .A(n_22), .Y(n_71) );
INVxp33_ASAP7_75t_SL g72 ( .A(n_19), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_35), .Y(n_73) );
INVxp33_ASAP7_75t_SL g74 ( .A(n_57), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_10), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_46), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_44), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_60), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_29), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_11), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_5), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_23), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_9), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_47), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_32), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_41), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_59), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_16), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_49), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_50), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_61), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_7), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_16), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_84), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_108), .B(n_0), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_64), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_93), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_64), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_73), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_87), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_81), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_67), .Y(n_122) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_67), .A2(n_36), .B(n_62), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_91), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_107), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_94), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_94), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_101), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_101), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_96), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_69), .B(n_1), .Y(n_137) );
NOR2xp33_ASAP7_75t_R g138 ( .A(n_66), .B(n_34), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_69), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_70), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_63), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_72), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_70), .B(n_3), .Y(n_150) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_123), .A2(n_109), .B(n_92), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_113), .B(n_85), .Y(n_153) );
OR2x2_ASAP7_75t_L g154 ( .A(n_142), .B(n_98), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_145), .B(n_74), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_117), .B(n_78), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_131), .B(n_98), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_142), .B(n_75), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_115), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_120), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_124), .B(n_100), .Y(n_168) );
OAI221xp5_ASAP7_75t_L g169 ( .A1(n_150), .A2(n_75), .B1(n_100), .B2(n_80), .C(n_104), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_112), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_113), .B(n_95), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_124), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_129), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_115), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_124), .B(n_80), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_112), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_111), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_112), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_116), .B(n_118), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_110), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_116), .B(n_118), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_122), .Y(n_189) );
CKINVDCx11_ASAP7_75t_R g190 ( .A(n_135), .Y(n_190) );
OR2x2_ASAP7_75t_SL g191 ( .A(n_150), .B(n_90), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_122), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_114), .Y(n_195) );
BUFx4f_ASAP7_75t_L g196 ( .A(n_121), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_119), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_135), .Y(n_198) );
OAI221xp5_ASAP7_75t_L g199 ( .A1(n_121), .A2(n_104), .B1(n_90), .B2(n_86), .C(n_71), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_135), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_125), .B(n_103), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_122), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_137), .B(n_109), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_119), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_119), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_127), .Y(n_208) );
INVx5_ASAP7_75t_L g209 ( .A(n_206), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_203), .B(n_143), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_137), .B1(n_143), .B2(n_83), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_185), .B(n_130), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_181), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_185), .B(n_130), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_185), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_190), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_181), .Y(n_217) );
NAND2xp33_ASAP7_75t_R g218 ( .A(n_200), .B(n_138), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_185), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_205), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_160), .B(n_143), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_196), .B(n_139), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_161), .B(n_132), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_196), .B(n_159), .Y(n_226) );
INVxp67_ASAP7_75t_SL g227 ( .A(n_205), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_198), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_168), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_196), .B(n_139), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_163), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_161), .B(n_132), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_167), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_174), .A2(n_125), .B1(n_148), .B2(n_147), .Y(n_237) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_168), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_154), .B(n_136), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_159), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_163), .B(n_147), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_184), .Y(n_242) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_183), .B(n_136), .C(n_148), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_184), .Y(n_244) );
NOR2x1_ASAP7_75t_L g245 ( .A(n_155), .B(n_144), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_174), .B(n_144), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_154), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_168), .A2(n_157), .B1(n_179), .B2(n_196), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_199), .B(n_186), .C(n_169), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_168), .A2(n_141), .B1(n_127), .B2(n_133), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_179), .B(n_141), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_202), .B(n_105), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_157), .B(n_127), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_184), .B(n_105), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_189), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_159), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_189), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_189), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_195), .B(n_87), .Y(n_262) );
O2A1O1Ixp5_ASAP7_75t_L g263 ( .A1(n_188), .A2(n_133), .B(n_128), .C(n_106), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_153), .B(n_133), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_153), .B(n_128), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_156), .B(n_171), .C(n_92), .Y(n_266) );
NOR3xp33_ASAP7_75t_SL g267 ( .A(n_171), .B(n_97), .C(n_99), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_191), .B(n_102), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_191), .B(n_97), .C(n_99), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_192), .B1(n_170), .B2(n_204), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g272 ( .A(n_221), .B(n_192), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_263), .A2(n_164), .B(n_180), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_216), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_240), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_227), .B(n_164), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_233), .B(n_175), .Y(n_279) );
NAND2xp33_ASAP7_75t_SL g280 ( .A(n_222), .B(n_159), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_226), .A2(n_164), .B(n_159), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_226), .A2(n_159), .B(n_151), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_170), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g284 ( .A(n_230), .B(n_170), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_227), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_210), .B(n_170), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_217), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_223), .B(n_204), .Y(n_290) );
OR2x6_ASAP7_75t_L g291 ( .A(n_262), .B(n_87), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_240), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_249), .A2(n_204), .B1(n_151), .B2(n_102), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_239), .B(n_204), .Y(n_294) );
INVxp33_ASAP7_75t_SL g295 ( .A(n_236), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_254), .B(n_151), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_254), .B(n_128), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_262), .B(n_68), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_230), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_215), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_259), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_238), .B(n_151), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_228), .A2(n_119), .B(n_140), .C(n_149), .Y(n_303) );
OAI22xp5_ASAP7_75t_SL g304 ( .A1(n_211), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_257), .B(n_206), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_224), .A2(n_177), .B(n_173), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_257), .B(n_140), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_213), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_220), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_219), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_225), .B(n_4), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_265), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_209), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_259), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_212), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_242), .Y(n_317) );
OR2x6_ASAP7_75t_L g318 ( .A(n_247), .B(n_235), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_286), .B(n_243), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_293), .B(n_267), .C(n_266), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_318), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_295), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_311), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_291), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_295), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_318), .A2(n_237), .B1(n_214), .B2(n_252), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_304), .A2(n_268), .B1(n_255), .B2(n_256), .Y(n_330) );
INVx4_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_318), .A2(n_268), .B1(n_245), .B2(n_255), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_278), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_313), .B(n_251), .Y(n_335) );
CKINVDCx14_ASAP7_75t_R g336 ( .A(n_274), .Y(n_336) );
NAND2xp33_ASAP7_75t_R g337 ( .A(n_274), .B(n_250), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_277), .Y(n_338) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_296), .A2(n_218), .B(n_224), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_313), .B(n_316), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_316), .B(n_250), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_279), .Y(n_342) );
NAND2xp33_ASAP7_75t_R g343 ( .A(n_291), .B(n_270), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_281), .A2(n_259), .B(n_232), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_232), .B1(n_252), .B2(n_229), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_275), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_308), .B(n_253), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_330), .A2(n_298), .B1(n_312), .B2(n_283), .Y(n_350) );
AO221x2_ASAP7_75t_L g351 ( .A1(n_320), .A2(n_267), .B1(n_270), .B2(n_10), .C(n_11), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g353 ( .A1(n_343), .A2(n_298), .B(n_275), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_345), .A2(n_298), .B1(n_308), .B2(n_275), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_344), .A2(n_282), .B(n_273), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_329), .A2(n_308), .B1(n_266), .B2(n_271), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_341), .B(n_290), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_340), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_345), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_342), .A2(n_307), .B1(n_297), .B2(n_271), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_332), .B(n_299), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_272), .B1(n_264), .B2(n_246), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_325), .A2(n_272), .B1(n_234), .B2(n_231), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_348), .B(n_284), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_338), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_319), .A2(n_322), .B1(n_349), .B2(n_325), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_337), .A2(n_218), .B(n_303), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_319), .A2(n_288), .B1(n_289), .B2(n_310), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_326), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_263), .B1(n_280), .B2(n_261), .C(n_260), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_352), .B(n_334), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_361), .B(n_324), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_355), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g381 ( .A1(n_350), .A2(n_328), .B1(n_324), .B2(n_319), .C1(n_349), .C2(n_334), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_359), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
INVx5_ASAP7_75t_SL g384 ( .A(n_375), .Y(n_384) );
BUFx10_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_321), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_357), .A2(n_349), .B1(n_321), .B2(n_331), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_368), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_374), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_339), .B(n_292), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_351), .A2(n_319), .B1(n_349), .B2(n_331), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_362), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_374), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_336), .B(n_328), .C(n_347), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_276), .B(n_315), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_375), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
NOR4xp25_ASAP7_75t_SL g403 ( .A(n_353), .B(n_280), .C(n_305), .D(n_326), .Y(n_403) );
OAI22xp5_ASAP7_75t_SL g404 ( .A1(n_366), .A2(n_284), .B1(n_333), .B2(n_346), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_367), .B(n_354), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_358), .B(n_333), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_351), .A2(n_289), .B1(n_288), .B2(n_314), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_356), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_357), .A2(n_305), .B1(n_317), .B2(n_269), .C(n_314), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_381), .A2(n_365), .B1(n_354), .B2(n_364), .C(n_371), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_383), .B(n_356), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_408), .B(n_351), .C(n_376), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_389), .B(n_351), .Y(n_416) );
OAI222xp33_ASAP7_75t_L g417 ( .A1(n_405), .A2(n_367), .B1(n_369), .B2(n_373), .C1(n_314), .C2(n_14), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_394), .B(n_140), .C(n_149), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_409), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_405), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_405), .A2(n_356), .B1(n_310), .B2(n_309), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_385), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_405), .A2(n_309), .B1(n_317), .B2(n_259), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_315), .B(n_292), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_384), .B(n_301), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g432 ( .A(n_378), .B(n_140), .C(n_149), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_383), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_391), .B(n_6), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_380), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_401), .B(n_9), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_149), .B1(n_306), .B2(n_182), .C(n_152), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_392), .B(n_12), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_382), .Y(n_440) );
NOR3xp33_ASAP7_75t_SL g441 ( .A(n_388), .B(n_180), .C(n_162), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_400), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_400), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_407), .B(n_12), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_402), .A2(n_13), .B(n_14), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_15), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_398), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_390), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_377), .B(n_15), .Y(n_451) );
NAND2x1p5_ASAP7_75t_SL g452 ( .A(n_396), .B(n_276), .Y(n_452) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_398), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_387), .B(n_17), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_387), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_406), .B(n_18), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_384), .B(n_21), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_440), .B(n_396), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_456), .B(n_384), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
NAND2xp33_ASAP7_75t_SL g463 ( .A(n_424), .B(n_404), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_456), .B(n_393), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_414), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_453), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_413), .B(n_393), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_413), .B(n_393), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_421), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_444), .B(n_395), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_414), .B(n_403), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_435), .B(n_410), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_419), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_420), .B(n_152), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_436), .B(n_152), .Y(n_477) );
NAND2xp33_ASAP7_75t_R g478 ( .A(n_425), .B(n_24), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_165), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_446), .B(n_162), .C(n_173), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_447), .B(n_182), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_411), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_429), .B(n_165), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_428), .A2(n_431), .B(n_450), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_421), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_433), .B(n_165), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_425), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_447), .B(n_182), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_422), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_411), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_422), .B(n_172), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_436), .B(n_172), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_427), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_426), .B(n_448), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_439), .B(n_172), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_426), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_424), .Y(n_499) );
NOR4xp25_ASAP7_75t_SL g500 ( .A(n_446), .B(n_194), .C(n_178), .D(n_177), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_426), .B(n_193), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_442), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_442), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_425), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_427), .B(n_301), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_412), .A2(n_301), .B1(n_277), .B2(n_285), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_427), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_439), .B(n_187), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_448), .B(n_193), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_463), .A2(n_415), .B1(n_432), .B2(n_416), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_503), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_505), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_473), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_473), .B(n_437), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_460), .B(n_445), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_480), .A2(n_415), .B1(n_418), .B2(n_423), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_475), .B(n_437), .Y(n_521) );
NAND3xp33_ASAP7_75t_SL g522 ( .A(n_500), .B(n_458), .C(n_441), .Y(n_522) );
OAI22xp33_ASAP7_75t_SL g523 ( .A1(n_495), .A2(n_459), .B1(n_454), .B2(n_455), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_475), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_484), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_466), .B(n_443), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_478), .A2(n_505), .B1(n_495), .B2(n_482), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_484), .B(n_451), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_474), .A2(n_417), .B1(n_434), .B2(n_418), .C(n_438), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_472), .A2(n_458), .B1(n_457), .B2(n_449), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_471), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_470), .A2(n_449), .B1(n_430), .B2(n_452), .C(n_457), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_510), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_491), .B(n_452), .Y(n_534) );
AOI221x1_ASAP7_75t_L g535 ( .A1(n_472), .A2(n_452), .B1(n_158), .B2(n_194), .C(n_178), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_485), .B(n_193), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_496), .B(n_187), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_489), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_509), .A2(n_158), .B(n_176), .Y(n_539) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_461), .B(n_301), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_499), .A2(n_176), .B1(n_187), .B2(n_285), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_496), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_498), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_507), .A2(n_176), .B1(n_277), .B2(n_244), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_461), .A2(n_277), .B1(n_209), .B2(n_258), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_486), .A2(n_207), .B(n_197), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_477), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_504), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_492), .A2(n_209), .B1(n_37), .B2(n_39), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_467), .B(n_31), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_467), .B(n_45), .Y(n_552) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_527), .A2(n_468), .A3(n_506), .B1(n_502), .B2(n_493), .C1(n_494), .C2(n_490), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_542), .B(n_502), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_519), .B(n_481), .Y(n_555) );
NAND2xp33_ASAP7_75t_L g556 ( .A(n_515), .B(n_502), .Y(n_556) );
NOR3xp33_ASAP7_75t_SL g557 ( .A(n_522), .B(n_511), .C(n_497), .Y(n_557) );
OAI211xp5_ASAP7_75t_L g558 ( .A1(n_513), .A2(n_464), .B(n_493), .C(n_508), .Y(n_558) );
NAND2xp33_ASAP7_75t_SL g559 ( .A(n_515), .B(n_464), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_520), .A2(n_462), .B1(n_469), .B2(n_487), .C(n_494), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_517), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_526), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_525), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_514), .B(n_512), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_548), .B(n_512), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_547), .Y(n_568) );
NOR3xp33_ASAP7_75t_SL g569 ( .A(n_550), .B(n_483), .C(n_479), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_531), .B(n_483), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g571 ( .A(n_530), .B(n_479), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_549), .B(n_476), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
NOR4xp25_ASAP7_75t_SL g574 ( .A(n_532), .B(n_476), .C(n_501), .D(n_488), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_534), .B(n_518), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_528), .B(n_488), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_555), .A2(n_523), .B1(n_529), .B2(n_521), .C(n_538), .Y(n_577) );
AOI22x1_ASAP7_75t_L g578 ( .A1(n_564), .A2(n_546), .B1(n_533), .B2(n_551), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_575), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_568), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_569), .A2(n_550), .B(n_546), .Y(n_581) );
OAI332xp33_ASAP7_75t_L g582 ( .A1(n_561), .A2(n_552), .A3(n_537), .B1(n_536), .B2(n_545), .B3(n_501), .C1(n_540), .C2(n_535), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_553), .B(n_539), .C(n_541), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_567), .B(n_544), .Y(n_584) );
INVxp33_ASAP7_75t_SL g585 ( .A(n_571), .Y(n_585) );
XNOR2x1_ASAP7_75t_L g586 ( .A(n_576), .B(n_51), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_573), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_556), .B(n_54), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_577), .A2(n_557), .B1(n_559), .B2(n_554), .Y(n_589) );
NAND4xp25_ASAP7_75t_SL g590 ( .A(n_577), .B(n_559), .C(n_570), .D(n_554), .Y(n_590) );
NAND2xp33_ASAP7_75t_SL g591 ( .A(n_586), .B(n_574), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_579), .B(n_572), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_585), .A2(n_572), .B1(n_566), .B2(n_556), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_582), .B(n_565), .C(n_563), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_581), .A2(n_566), .B1(n_562), .B2(n_560), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_580), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g597 ( .A1(n_588), .A2(n_583), .B1(n_578), .B2(n_584), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_588), .Y(n_598) );
AOI211x1_ASAP7_75t_L g599 ( .A1(n_587), .A2(n_581), .B(n_558), .C(n_583), .Y(n_599) );
OAI22xp5_ASAP7_75t_SL g600 ( .A1(n_585), .A2(n_167), .B1(n_588), .B2(n_581), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_598), .B(n_589), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_596), .Y(n_602) );
NAND4xp25_ASAP7_75t_SL g603 ( .A(n_593), .B(n_595), .C(n_594), .D(n_599), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_602), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_601), .A2(n_597), .B1(n_600), .B2(n_592), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_603), .B(n_590), .C(n_591), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_604), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_605), .Y(n_608) );
INVx4_ASAP7_75t_L g609 ( .A(n_607), .Y(n_609) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_609), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_610), .A2(n_608), .B(n_606), .Y(n_611) );
endmodule