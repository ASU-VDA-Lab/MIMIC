module fake_jpeg_29884_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_8),
.B(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_21),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_12),
.B1(n_15),
.B2(n_11),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_18),
.B(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_27),
.B1(n_3),
.B2(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_29),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_11),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_52),
.B1(n_39),
.B2(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_22),
.B1(n_12),
.B2(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.C(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_28),
.C(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_58),
.C(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_53),
.B1(n_59),
.B2(n_41),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_41),
.C(n_40),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_66),
.C(n_63),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.C(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_72),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_70),
.B1(n_71),
.B2(n_48),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_21),
.C(n_10),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_21),
.B(n_10),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_80),
.B(n_10),
.C(n_30),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_40),
.Y(n_84)
);


endmodule