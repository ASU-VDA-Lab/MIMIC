module fake_jpeg_1956_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_62),
.Y(n_89)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_54),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_59),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_67),
.Y(n_90)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_29),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_22),
.B(n_27),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_75),
.Y(n_103)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_101),
.B1(n_108),
.B2(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_26),
.B1(n_41),
.B2(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_41),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_54),
.Y(n_97)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_115),
.B1(n_102),
.B2(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_31),
.B1(n_35),
.B2(n_42),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_57),
.A2(n_42),
.B1(n_8),
.B2(n_10),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_43),
.A2(n_10),
.B1(n_58),
.B2(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_45),
.B(n_46),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_73),
.B1(n_79),
.B2(n_55),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_43),
.B1(n_111),
.B2(n_64),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_101),
.B(n_103),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_127),
.B(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_137),
.B1(n_138),
.B2(n_122),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_105),
.B(n_108),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_132),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_105),
.B(n_110),
.C(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_82),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_133),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_119),
.B1(n_118),
.B2(n_106),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_138),
.B1(n_147),
.B2(n_120),
.Y(n_157)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_114),
.B1(n_109),
.B2(n_99),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_85),
.C(n_109),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_135),
.C(n_129),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_149),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_89),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_148),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_93),
.A2(n_87),
.B1(n_101),
.B2(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_112),
.B(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_90),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_89),
.B(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_130),
.Y(n_155)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_126),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_141),
.B1(n_142),
.B2(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_132),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_127),
.B(n_123),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_170),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_152),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_172),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_157),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_181),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_172),
.Y(n_200)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_191),
.B1(n_169),
.B2(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_192),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_142),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_193),
.C(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_168),
.C(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_202),
.C(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_158),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_199),
.B(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_175),
.C(n_165),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_165),
.C(n_156),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_180),
.C(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_211),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

AO221x1_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_185),
.B1(n_154),
.B2(n_173),
.C(n_177),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_191),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_225),
.B(n_217),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_203),
.C(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_207),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_180),
.B(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_231),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_217),
.CI(n_219),
.CON(n_229),
.SN(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_218),
.B(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_214),
.B1(n_212),
.B2(n_219),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_204),
.B(n_213),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_232),
.C(n_187),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_216),
.A3(n_191),
.B1(n_210),
.B2(n_178),
.C1(n_220),
.C2(n_184),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_237),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_240),
.B(n_210),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_220),
.Y(n_242)
);


endmodule