module real_aes_9024_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_713, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_713;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g172 ( .A1(n_0), .A2(n_173), .B(n_174), .C(n_178), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_1), .B(n_167), .Y(n_180) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_3), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_4), .A2(n_141), .B(n_158), .C(n_465), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_161), .B(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_6), .A2(n_161), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_7), .B(n_167), .Y(n_492) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_8), .A2(n_133), .B(n_220), .Y(n_219) );
AND2x6_ASAP7_75t_L g158 ( .A(n_9), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_10), .A2(n_141), .B(n_158), .C(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g457 ( .A(n_11), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_40), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_13), .B(n_177), .Y(n_467) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_15), .B(n_152), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_16), .A2(n_153), .B(n_476), .C(n_478), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_17), .B(n_167), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_18), .A2(n_66), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_18), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_19), .B(n_210), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_141), .B(n_204), .C(n_209), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_21), .A2(n_176), .B(n_228), .C(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_22), .B(n_177), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_23), .B(n_177), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_24), .Y(n_495) );
INVx1_ASAP7_75t_L g507 ( .A(n_25), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_26), .A2(n_141), .B(n_209), .C(n_223), .Y(n_222) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_28), .Y(n_463) );
INVx1_ASAP7_75t_L g524 ( .A(n_29), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_30), .A2(n_161), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g143 ( .A(n_31), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_32), .A2(n_156), .B(n_188), .C(n_189), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_33), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_34), .A2(n_176), .B(n_489), .C(n_491), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_35), .A2(n_122), .B1(n_417), .B2(n_418), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_35), .Y(n_417) );
INVxp67_ASAP7_75t_L g525 ( .A(n_36), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_37), .B(n_225), .Y(n_224) );
CKINVDCx14_ASAP7_75t_R g487 ( .A(n_38), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_39), .A2(n_141), .B(n_209), .C(n_506), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_41), .A2(n_429), .B1(n_697), .B2(n_698), .C1(n_704), .C2(n_708), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_42), .A2(n_178), .B(n_455), .C(n_456), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_43), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_44), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_45), .B(n_152), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_46), .B(n_161), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_47), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_48), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_49), .A2(n_104), .B1(n_115), .B2(n_711), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_50), .A2(n_156), .B(n_188), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g175 ( .A(n_51), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_52), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_52), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_53), .A2(n_84), .B1(n_702), .B2(n_703), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_53), .Y(n_703) );
INVx1_ASAP7_75t_L g250 ( .A(n_54), .Y(n_250) );
INVx1_ASAP7_75t_L g445 ( .A(n_55), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_56), .B(n_161), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_57), .Y(n_213) );
CKINVDCx14_ASAP7_75t_R g453 ( .A(n_58), .Y(n_453) );
INVx1_ASAP7_75t_L g159 ( .A(n_59), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_60), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_61), .B(n_167), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_62), .A2(n_148), .B(n_208), .C(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
INVx1_ASAP7_75t_SL g490 ( .A(n_64), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_66), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_67), .B(n_152), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_68), .B(n_167), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_69), .B(n_153), .Y(n_239) );
INVx1_ASAP7_75t_L g498 ( .A(n_70), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_71), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_72), .B(n_192), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_73), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_74), .Y(n_264) );
INVx1_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_76), .A2(n_161), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_77), .B(n_424), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_78), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_79), .A2(n_161), .B(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_80), .A2(n_202), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g474 ( .A(n_81), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_82), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_83), .B(n_191), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_84), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_85), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_86), .A2(n_161), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g477 ( .A(n_87), .Y(n_477) );
INVx2_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx1_ASAP7_75t_L g466 ( .A(n_89), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_90), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_91), .B(n_177), .Y(n_240) );
INVx2_ASAP7_75t_L g110 ( .A(n_92), .Y(n_110) );
OR2x2_ASAP7_75t_L g422 ( .A(n_92), .B(n_111), .Y(n_422) );
OR2x2_ASAP7_75t_L g432 ( .A(n_92), .B(n_112), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_93), .A2(n_141), .B(n_156), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_94), .B(n_161), .Y(n_186) );
INVx1_ASAP7_75t_L g190 ( .A(n_95), .Y(n_190) );
INVxp67_ASAP7_75t_L g267 ( .A(n_96), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_97), .B(n_133), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
INVx1_ASAP7_75t_L g235 ( .A(n_100), .Y(n_235) );
INVx2_ASAP7_75t_L g448 ( .A(n_101), .Y(n_448) );
AND2x2_ASAP7_75t_L g252 ( .A(n_102), .B(n_195), .Y(n_252) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g711 ( .A(n_105), .Y(n_711) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g708 ( .A(n_108), .Y(n_708) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g435 ( .A(n_110), .B(n_112), .Y(n_435) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_427), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g710 ( .A(n_118), .Y(n_710) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_419), .B(n_423), .Y(n_120) );
INVx1_ASAP7_75t_L g418 ( .A(n_122), .Y(n_418) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx2_ASAP7_75t_L g433 ( .A(n_126), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_126), .A2(n_431), .B1(n_706), .B2(n_707), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_360), .Y(n_126) );
AND4x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_300), .C(n_315), .D(n_340), .Y(n_127) );
NOR2xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_273), .Y(n_128) );
OAI21xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_181), .B(n_253), .Y(n_129) );
AND2x2_ASAP7_75t_L g303 ( .A(n_130), .B(n_199), .Y(n_303) );
AND2x2_ASAP7_75t_L g316 ( .A(n_130), .B(n_198), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_130), .B(n_182), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_130), .Y(n_370) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
INVx2_ASAP7_75t_L g287 ( .A(n_131), .Y(n_287) );
BUFx2_ASAP7_75t_L g314 ( .A(n_131), .Y(n_314) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_164), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_132), .B(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_132), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_132), .A2(n_234), .B(n_241), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_132), .B(n_470), .Y(n_469) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_132), .A2(n_494), .B(n_500), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_132), .B(n_510), .Y(n_509) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_222), .Y(n_220) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_133), .Y(n_261) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g243 ( .A(n_134), .Y(n_243) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_135), .B(n_136), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_160), .Y(n_139) );
INVx5_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
BUFx3_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx1_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_145), .B(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
INVx1_ASAP7_75t_L g225 ( .A(n_145), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_149), .B(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_149), .B(n_477), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_149), .A2(n_152), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
INVx2_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_152), .B(n_267), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_152), .A2(n_207), .B(n_507), .C(n_508), .Y(n_506) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_153), .B(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g491 ( .A(n_155), .Y(n_491) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_157), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_157), .A2(n_171), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g444 ( .A1(n_157), .A2(n_171), .B(n_445), .C(n_446), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_157), .A2(n_171), .B(n_453), .C(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_157), .A2(n_171), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_157), .A2(n_171), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_157), .A2(n_171), .B(n_521), .C(n_522), .Y(n_520) );
INVx4_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g161 ( .A(n_158), .B(n_162), .Y(n_161) );
BUFx3_ASAP7_75t_L g209 ( .A(n_158), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_158), .B(n_162), .Y(n_236) );
BUFx2_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx1_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
AND2x2_ASAP7_75t_L g254 ( .A(n_166), .B(n_199), .Y(n_254) );
INVx2_ASAP7_75t_L g270 ( .A(n_166), .Y(n_270) );
AND2x2_ASAP7_75t_L g279 ( .A(n_166), .B(n_198), .Y(n_279) );
AND2x2_ASAP7_75t_L g358 ( .A(n_166), .B(n_287), .Y(n_358) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_180), .Y(n_166) );
INVx2_ASAP7_75t_L g188 ( .A(n_171), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_176), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g455 ( .A(n_177), .Y(n_455) );
INVx2_ASAP7_75t_L g468 ( .A(n_178), .Y(n_468) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
INVx1_ASAP7_75t_L g478 ( .A(n_179), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_215), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_182), .B(n_285), .Y(n_323) );
INVx1_ASAP7_75t_L g411 ( .A(n_182), .Y(n_411) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
AND2x2_ASAP7_75t_L g269 ( .A(n_183), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g283 ( .A(n_183), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_183), .Y(n_312) );
OR2x2_ASAP7_75t_L g344 ( .A(n_183), .B(n_286), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_183), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g385 ( .A(n_183), .B(n_354), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_183), .B(n_254), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_183), .B(n_314), .Y(n_410) );
AND2x2_ASAP7_75t_L g416 ( .A(n_183), .B(n_303), .Y(n_416) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx2_ASAP7_75t_L g276 ( .A(n_184), .Y(n_276) );
AND2x2_ASAP7_75t_L g306 ( .A(n_184), .B(n_286), .Y(n_306) );
AND2x2_ASAP7_75t_L g339 ( .A(n_184), .B(n_299), .Y(n_339) );
AND2x2_ASAP7_75t_L g359 ( .A(n_184), .B(n_199), .Y(n_359) );
AND2x2_ASAP7_75t_L g393 ( .A(n_184), .B(n_259), .Y(n_393) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_196), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_195), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .C(n_194), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_191), .A2(n_194), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_191), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_191), .A2(n_468), .B(n_498), .C(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g211 ( .A(n_195), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_195), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_195), .A2(n_247), .B(n_248), .Y(n_246) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_195), .A2(n_451), .B(n_458), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_195), .A2(n_236), .B(n_504), .C(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g299 ( .A(n_198), .B(n_270), .Y(n_299) );
AND2x2_ASAP7_75t_L g310 ( .A(n_198), .B(n_306), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_198), .B(n_286), .Y(n_349) );
INVx2_ASAP7_75t_L g364 ( .A(n_198), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_198), .B(n_298), .Y(n_387) );
AND2x2_ASAP7_75t_L g406 ( .A(n_198), .B(n_358), .Y(n_406) );
INVx5_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_199), .Y(n_305) );
AND2x2_ASAP7_75t_L g313 ( .A(n_199), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g354 ( .A(n_199), .B(n_270), .Y(n_354) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_212), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_210), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_208), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_211), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_214), .A2(n_462), .B(n_469), .Y(n_461) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_230), .Y(n_216) );
AND2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_260), .Y(n_277) );
INVx1_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_218), .B(n_233), .Y(n_257) );
OR2x2_ASAP7_75t_L g290 ( .A(n_218), .B(n_260), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_218), .B(n_260), .Y(n_295) );
AND2x2_ASAP7_75t_L g322 ( .A(n_218), .B(n_259), .Y(n_322) );
AND2x2_ASAP7_75t_L g374 ( .A(n_218), .B(n_232), .Y(n_374) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_219), .B(n_244), .Y(n_282) );
AND2x2_ASAP7_75t_L g318 ( .A(n_219), .B(n_233), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_226), .B(n_227), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_227), .A2(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_230), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g308 ( .A(n_231), .B(n_290), .Y(n_308) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_244), .Y(n_231) );
OAI322xp33_ASAP7_75t_L g273 ( .A1(n_232), .A2(n_274), .A3(n_278), .B1(n_280), .B2(n_283), .C1(n_288), .C2(n_296), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_232), .B(n_259), .Y(n_281) );
OR2x2_ASAP7_75t_L g291 ( .A(n_232), .B(n_245), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_232), .B(n_245), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_232), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_232), .B(n_260), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_232), .B(n_389), .Y(n_388) );
INVx5_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_233), .B(n_277), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_236), .A2(n_463), .B(n_464), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_236), .A2(n_495), .B(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g518 ( .A(n_243), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_244), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g271 ( .A(n_244), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_244), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g333 ( .A(n_244), .B(n_260), .Y(n_333) );
AOI211xp5_ASAP7_75t_SL g361 ( .A1(n_244), .A2(n_362), .B(n_365), .C(n_377), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_244), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g399 ( .A(n_244), .B(n_374), .Y(n_399) );
INVx5_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g327 ( .A(n_245), .B(n_260), .Y(n_327) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_245), .Y(n_336) );
AND2x2_ASAP7_75t_L g376 ( .A(n_245), .B(n_374), .Y(n_376) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_245), .B(n_277), .Y(n_407) );
AND2x2_ASAP7_75t_L g414 ( .A(n_245), .B(n_373), .Y(n_414) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_252), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B1(n_269), .B2(n_271), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_254), .B(n_276), .Y(n_324) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
OR2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_333), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g380 ( .A1(n_257), .A2(n_381), .B1(n_383), .B2(n_384), .C(n_386), .Y(n_380) );
INVx2_ASAP7_75t_L g319 ( .A(n_258), .Y(n_319) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g382 ( .A(n_259), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_259), .B(n_374), .Y(n_395) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_L g337 ( .A(n_260), .Y(n_337) );
AND2x2_ASAP7_75t_L g373 ( .A(n_260), .B(n_374), .Y(n_373) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_268), .Y(n_260) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_261), .A2(n_443), .B(n_449), .Y(n_442) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_261), .A2(n_472), .B(n_479), .Y(n_471) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_261), .A2(n_485), .B(n_492), .Y(n_484) );
AND2x2_ASAP7_75t_L g375 ( .A(n_269), .B(n_314), .Y(n_375) );
AND2x2_ASAP7_75t_L g285 ( .A(n_270), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_270), .B(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_SL g356 ( .A(n_272), .B(n_319), .Y(n_356) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g362 ( .A(n_275), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g348 ( .A(n_276), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g413 ( .A(n_276), .B(n_358), .Y(n_413) );
INVx2_ASAP7_75t_L g346 ( .A(n_277), .Y(n_346) );
NAND4xp25_ASAP7_75t_SL g409 ( .A(n_278), .B(n_410), .C(n_411), .D(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_279), .B(n_343), .Y(n_378) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_SL g415 ( .A(n_282), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_SL g377 ( .A1(n_283), .A2(n_346), .B(n_350), .C(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g372 ( .A(n_285), .B(n_364), .Y(n_372) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_286), .Y(n_298) );
INVx1_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_292), .C(n_294), .Y(n_288) );
AND2x2_ASAP7_75t_L g309 ( .A(n_289), .B(n_293), .Y(n_309) );
OAI322xp33_ASAP7_75t_SL g347 ( .A1(n_289), .A2(n_348), .A3(n_350), .B1(n_351), .B2(n_355), .C1(n_356), .C2(n_357), .Y(n_347) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g369 ( .A(n_291), .B(n_295), .Y(n_369) );
INVx1_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
INVx1_ASAP7_75t_SL g368 ( .A(n_295), .Y(n_368) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AOI222xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B1(n_309), .B2(n_310), .C1(n_311), .C2(n_713), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
OAI322xp33_ASAP7_75t_L g390 ( .A1(n_302), .A2(n_364), .A3(n_369), .B1(n_391), .B2(n_392), .C1(n_394), .C2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_303), .A2(n_317), .B1(n_341), .B2(n_345), .C(n_347), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OAI222xp33_ASAP7_75t_L g320 ( .A1(n_308), .A2(n_321), .B1(n_323), .B2(n_324), .C1(n_325), .C2(n_328), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_310), .A2(n_317), .B1(n_387), .B2(n_388), .Y(n_386) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_320), .C(n_331), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_317), .A2(n_354), .B(n_397), .C(n_400), .Y(n_396) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_318), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g389 ( .A(n_322), .Y(n_389) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_329), .B(n_354), .Y(n_383) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_338), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_332), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_404), .Y(n_400) );
INVxp33_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_336), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_343), .B(n_354), .Y(n_394) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g405 ( .A(n_358), .B(n_364), .Y(n_405) );
AND4x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_379), .C(n_396), .D(n_408), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B1(n_369), .B2(n_370), .C(n_371), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_375), .B2(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
INVx1_ASAP7_75t_SL g391 ( .A(n_376), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_390), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_392), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_399), .A2(n_405), .B1(n_406), .B2(n_407), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g426 ( .A(n_422), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_423), .A2(n_428), .B(n_709), .Y(n_427) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_434), .B2(n_436), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx6_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g706 ( .A(n_435), .Y(n_706) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g707 ( .A(n_437), .Y(n_707) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_623), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_565), .C(n_595), .D(n_605), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_480), .B(n_528), .C(n_555), .Y(n_439) );
OAI222xp33_ASAP7_75t_L g650 ( .A1(n_440), .A2(n_570), .B1(n_651), .B2(n_652), .C1(n_653), .C2(n_654), .Y(n_650) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_459), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g576 ( .A1(n_441), .A2(n_563), .A3(n_564), .B1(n_577), .B2(n_582), .B3(n_584), .Y(n_576) );
OAI211xp5_ASAP7_75t_SL g633 ( .A1(n_441), .A2(n_634), .B(n_636), .C(n_638), .Y(n_633) );
OR2x2_ASAP7_75t_L g649 ( .A(n_441), .B(n_635), .Y(n_649) );
INVx1_ASAP7_75t_L g682 ( .A(n_441), .Y(n_682) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_450), .Y(n_441) );
INVx2_ASAP7_75t_L g559 ( .A(n_442), .Y(n_559) );
AND2x2_ASAP7_75t_L g575 ( .A(n_442), .B(n_471), .Y(n_575) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_442), .Y(n_610) );
AND2x2_ASAP7_75t_L g639 ( .A(n_442), .B(n_450), .Y(n_639) );
INVx2_ASAP7_75t_L g539 ( .A(n_450), .Y(n_539) );
BUFx3_ASAP7_75t_L g547 ( .A(n_450), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_450), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g558 ( .A(n_450), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_450), .B(n_460), .Y(n_587) );
AND2x2_ASAP7_75t_L g656 ( .A(n_450), .B(n_590), .Y(n_656) );
INVx2_ASAP7_75t_SL g550 ( .A(n_459), .Y(n_550) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_460), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g592 ( .A(n_460), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_460), .B(n_559), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_460), .B(n_588), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_460), .B(n_590), .Y(n_635) );
AND2x2_ASAP7_75t_L g694 ( .A(n_460), .B(n_639), .Y(n_694) );
INVx4_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g564 ( .A(n_461), .B(n_471), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_461), .B(n_575), .Y(n_574) );
BUFx3_ASAP7_75t_L g596 ( .A(n_461), .Y(n_596) );
AND3x2_ASAP7_75t_L g655 ( .A(n_461), .B(n_656), .C(n_657), .Y(n_655) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_471), .Y(n_546) );
INVx1_ASAP7_75t_SL g590 ( .A(n_471), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_471), .B(n_539), .C(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_511), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_481), .A2(n_574), .B(n_626), .C(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_483), .B(n_502), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_483), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_SL g642 ( .A(n_483), .Y(n_642) );
AND2x2_ASAP7_75t_L g663 ( .A(n_483), .B(n_513), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_483), .B(n_572), .Y(n_691) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
AND2x2_ASAP7_75t_L g536 ( .A(n_484), .B(n_527), .Y(n_536) );
INVx2_ASAP7_75t_L g543 ( .A(n_484), .Y(n_543) );
AND2x2_ASAP7_75t_L g563 ( .A(n_484), .B(n_513), .Y(n_563) );
AND2x2_ASAP7_75t_L g613 ( .A(n_484), .B(n_502), .Y(n_613) );
INVx1_ASAP7_75t_L g617 ( .A(n_484), .Y(n_617) );
INVx2_ASAP7_75t_SL g527 ( .A(n_493), .Y(n_527) );
BUFx2_ASAP7_75t_L g553 ( .A(n_493), .Y(n_553) );
AND2x2_ASAP7_75t_L g680 ( .A(n_493), .B(n_502), .Y(n_680) );
INVx3_ASAP7_75t_SL g513 ( .A(n_502), .Y(n_513) );
AND2x2_ASAP7_75t_L g535 ( .A(n_502), .B(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g542 ( .A(n_502), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g572 ( .A(n_502), .B(n_532), .Y(n_572) );
OR2x2_ASAP7_75t_L g581 ( .A(n_502), .B(n_527), .Y(n_581) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_502), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_502), .B(n_557), .Y(n_604) );
AND2x2_ASAP7_75t_L g632 ( .A(n_502), .B(n_515), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_502), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g670 ( .A(n_502), .B(n_514), .Y(n_670) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_L g594 ( .A(n_513), .B(n_543), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_513), .B(n_536), .Y(n_622) );
AND2x2_ASAP7_75t_L g640 ( .A(n_513), .B(n_557), .Y(n_640) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_527), .Y(n_514) );
AND2x2_ASAP7_75t_L g541 ( .A(n_515), .B(n_527), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_515), .B(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g579 ( .A(n_515), .Y(n_579) );
OR2x2_ASAP7_75t_L g627 ( .A(n_515), .B(n_547), .Y(n_627) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_519), .B(n_526), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_517), .A2(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g533 ( .A(n_519), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_526), .Y(n_534) );
AND2x2_ASAP7_75t_L g562 ( .A(n_527), .B(n_532), .Y(n_562) );
INVx1_ASAP7_75t_L g570 ( .A(n_527), .Y(n_570) );
AND2x2_ASAP7_75t_L g665 ( .A(n_527), .B(n_543), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_537), .B1(n_540), .B2(n_544), .C1(n_548), .C2(n_551), .Y(n_528) );
INVx1_ASAP7_75t_L g660 ( .A(n_529), .Y(n_660) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AND2x2_ASAP7_75t_L g556 ( .A(n_530), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g567 ( .A(n_530), .B(n_536), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_530), .B(n_558), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g605 ( .A1(n_530), .A2(n_606), .B1(n_611), .B2(n_612), .C1(n_620), .C2(n_622), .Y(n_605) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g593 ( .A(n_532), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_532), .B(n_613), .Y(n_653) );
AND2x2_ASAP7_75t_L g664 ( .A(n_532), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g672 ( .A(n_535), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_537), .B(n_588), .Y(n_651) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_539), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx3_ASAP7_75t_L g554 ( .A(n_542), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_542), .A2(n_645), .B(n_648), .C(n_650), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_542), .B(n_579), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_542), .B(n_562), .Y(n_684) );
AND2x2_ASAP7_75t_L g557 ( .A(n_543), .B(n_553), .Y(n_557) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g584 ( .A(n_546), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_547), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g636 ( .A(n_547), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g675 ( .A(n_547), .B(n_575), .Y(n_675) );
INVx1_ASAP7_75t_L g687 ( .A(n_547), .Y(n_687) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_550), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g668 ( .A(n_553), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_558), .B(n_560), .C(n_564), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_556), .A2(n_586), .B1(n_601), .B2(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_557), .B(n_571), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_557), .B(n_579), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_558), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g621 ( .A(n_558), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_558), .B(n_608), .Y(n_628) );
INVx2_ASAP7_75t_L g589 ( .A(n_559), .Y(n_589) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NOR4xp25_ASAP7_75t_L g566 ( .A(n_563), .B(n_567), .C(n_568), .D(n_571), .Y(n_566) );
INVx1_ASAP7_75t_SL g637 ( .A(n_564), .Y(n_637) );
AND2x2_ASAP7_75t_L g681 ( .A(n_564), .B(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_573), .B(n_576), .C(n_585), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_572), .B(n_642), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_574), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_SL g647 ( .A(n_575), .Y(n_647) );
AND2x2_ASAP7_75t_L g686 ( .A(n_575), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_579), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_583), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_584), .B(n_609), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_591), .B(n_593), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g661 ( .A(n_588), .Y(n_661) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g689 ( .A(n_589), .Y(n_689) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_590), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_600), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_596), .Y(n_608) );
OR2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI21xp33_ASAP7_75t_SL g641 ( .A1(n_599), .A2(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_603), .A2(n_630), .B1(n_633), .B2(n_640), .C(n_641), .Y(n_629) );
INVx1_ASAP7_75t_SL g673 ( .A(n_604), .Y(n_673) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g620 ( .A(n_608), .B(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g657 ( .A(n_610), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_617), .B2(n_618), .Y(n_612) );
INVx1_ASAP7_75t_L g652 ( .A(n_613), .Y(n_652) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_616), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_658), .C(n_671), .D(n_683), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_629), .C(n_644), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_627), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_634), .B(n_639), .Y(n_643) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI221xp5_ASAP7_75t_SL g671 ( .A1(n_646), .A2(n_672), .B1(n_673), .B2(n_674), .C(n_676), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_648), .A2(n_663), .B(n_664), .C(n_666), .Y(n_662) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_649), .A2(n_667), .B1(n_669), .B2(n_670), .Y(n_666) );
INVx2_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_661), .C(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g677 ( .A(n_670), .Y(n_677) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_685), .B1(n_688), .B2(n_690), .C(n_692), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
endmodule