module fake_netlist_6_2138_n_1820 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1820);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1820;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_924;
wire n_475;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_172),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_20),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_35),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_106),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_26),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_174),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_131),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_96),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_34),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_85),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_31),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_4),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_83),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_40),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_155),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_7),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_135),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_23),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_145),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_27),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_0),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_18),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_66),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_20),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_43),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_151),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_28),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_56),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_77),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_60),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_53),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_56),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_87),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_22),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_150),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_12),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_89),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_108),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_137),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_86),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_95),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_29),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_104),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_52),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_162),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_94),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_110),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_156),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_147),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_139),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_158),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_173),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_115),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_175),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_112),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_59),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_93),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_82),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_65),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_142),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_138),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_134),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_80),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_18),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_2),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_101),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_24),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_8),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_148),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_21),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_116),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_11),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_75),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_149),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_0),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_5),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_88),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_98),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_120),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_9),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_40),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_132),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_130),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_64),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_141),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_49),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_57),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_50),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_128),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_63),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_38),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_67),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_19),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_68),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_31),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_69),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_46),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_28),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_92),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_127),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_43),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_146),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_126),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_16),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_84),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_121),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_14),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_9),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_160),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_15),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_105),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_129),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_114),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_154),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_100),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_27),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_17),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_240),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_206),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_245),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_206),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_198),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_198),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_206),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_201),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_206),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_180),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_206),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_206),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_237),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_237),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_237),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_184),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_237),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_237),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_237),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_237),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_263),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_263),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_263),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_263),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_182),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_263),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_263),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_211),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_263),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_196),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_184),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_201),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_261),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_231),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_212),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_178),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_185),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_214),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_202),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_234),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_238),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_220),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_221),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_248),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_189),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_231),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_258),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_268),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_274),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_192),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_312),
.Y(n_415)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_261),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_186),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_281),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_288),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_183),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_303),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_308),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_186),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_311),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_288),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_183),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_225),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_227),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_189),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_229),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_265),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_231),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_266),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_265),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_230),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_231),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_328),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_205),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_205),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_181),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_188),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_301),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_183),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_207),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_232),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_209),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_344),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_301),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_239),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_246),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_353),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_254),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_361),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_416),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_197),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_197),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_339),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_339),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_190),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_360),
.A2(n_335),
.B1(n_226),
.B2(n_276),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_190),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_416),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_415),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_440),
.B(n_191),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_223),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_417),
.B(n_223),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_390),
.B(n_236),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_364),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_367),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_305),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_455),
.B(n_177),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_380),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_381),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_382),
.B(n_236),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_370),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_369),
.B(n_191),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_414),
.B(n_314),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_382),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_383),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_372),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_373),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_383),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_384),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_397),
.B(n_292),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_384),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_385),
.B(n_193),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_365),
.B(n_226),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_366),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_388),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_396),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_399),
.B(n_292),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_438),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_441),
.B(n_305),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_362),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_370),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_410),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_432),
.B(n_307),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_432),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_368),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_437),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_391),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_459),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_459),
.Y(n_538)
);

CKINVDCx6p67_ASAP7_75t_R g539 ( 
.A(n_531),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_457),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_491),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_461),
.B(n_386),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_461),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_479),
.B(n_394),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_492),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_486),
.B(n_377),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_500),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_519),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_484),
.B(n_393),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_484),
.B(n_395),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_486),
.B(n_392),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_394),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_465),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_469),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_495),
.B(n_446),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_495),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_469),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_478),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_458),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_458),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_519),
.B(n_389),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_504),
.B(n_449),
.C(n_398),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_504),
.B(n_389),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_488),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_491),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_514),
.B(n_406),
.C(n_402),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_501),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_487),
.B(n_431),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_526),
.B(n_307),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_458),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_502),
.B(n_473),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_518),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_527),
.B(n_406),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_473),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_500),
.A2(n_409),
.B1(n_451),
.B2(n_429),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_487),
.B(n_431),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_489),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_495),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_527),
.B(n_407),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_481),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_496),
.B(n_400),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_491),
.B(n_231),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_490),
.B(n_434),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_502),
.B(n_407),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_489),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_498),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_526),
.B(n_362),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_427),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_528),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_498),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_525),
.B(n_428),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_528),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_482),
.B(n_419),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_528),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_531),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_499),
.B(n_428),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_518),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_522),
.B(n_420),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_506),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_500),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_490),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_530),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_530),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_526),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_517),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_496),
.A2(n_250),
.B1(n_283),
.B2(n_218),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_500),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_458),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_515),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_462),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_500),
.A2(n_314),
.B1(n_334),
.B2(n_401),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_462),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_462),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_480),
.B(n_430),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_490),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_529),
.A2(n_334),
.B(n_215),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_493),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_477),
.B(n_434),
.Y(n_657)
);

CKINVDCx11_ASAP7_75t_R g658 ( 
.A(n_517),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_477),
.B(n_403),
.Y(n_659)
);

AO22x2_ASAP7_75t_L g660 ( 
.A1(n_477),
.A2(n_351),
.B1(n_222),
.B2(n_228),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_480),
.B(n_430),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_493),
.B(n_435),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_534),
.Y(n_663)
);

BUFx4f_ASAP7_75t_L g664 ( 
.A(n_492),
.Y(n_664)
);

AO22x2_ASAP7_75t_L g665 ( 
.A1(n_529),
.A2(n_290),
.B1(n_256),
.B2(n_309),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_483),
.B(n_435),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_529),
.A2(n_253),
.B1(n_355),
.B2(n_259),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_510),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_492),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_491),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_534),
.Y(n_673)
);

NOR2x1p5_ASAP7_75t_L g674 ( 
.A(n_483),
.B(n_363),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_512),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_462),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_462),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_510),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_493),
.B(n_448),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_494),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_562),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_540),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_555),
.B(n_453),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_561),
.B(n_453),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_557),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_618),
.B(n_454),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_584),
.B(n_231),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_562),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_600),
.B(n_492),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_548),
.B(n_529),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_596),
.B(n_266),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_550),
.B(n_276),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_548),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_559),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_574),
.B(n_454),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_666),
.B(n_456),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_639),
.B(n_675),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_574),
.B(n_456),
.Y(n_698)
);

O2A1O1Ixp5_ASAP7_75t_L g699 ( 
.A1(n_540),
.A2(n_529),
.B(n_466),
.C(n_476),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_660),
.A2(n_523),
.B1(n_512),
.B2(n_347),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_594),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_594),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_606),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_675),
.B(n_497),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_606),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_549),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_547),
.A2(n_503),
.B(n_494),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_615),
.B(n_497),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_615),
.B(n_497),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_611),
.B(n_271),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_627),
.B(n_647),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_624),
.B(n_324),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_654),
.B(n_193),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_627),
.B(n_497),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_570),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_617),
.Y(n_719)
);

BUFx8_ASAP7_75t_L g720 ( 
.A(n_551),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_554),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_647),
.B(n_497),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_570),
.B(n_517),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_636),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_617),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_497),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_660),
.A2(n_523),
.B1(n_512),
.B2(n_347),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_556),
.B(n_507),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_558),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_591),
.B(n_194),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_507),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_586),
.A2(n_252),
.B1(n_523),
.B2(n_445),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_566),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_567),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_568),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_569),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_569),
.B(n_507),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_578),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_578),
.B(n_597),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_657),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_633),
.A2(n_604),
.B1(n_614),
.B2(n_558),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_607),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_607),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_585),
.B(n_426),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_613),
.B(n_507),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_638),
.B(n_507),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_620),
.B(n_507),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_620),
.B(n_516),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_614),
.A2(n_318),
.B1(n_297),
.B2(n_247),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_635),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_635),
.B(n_516),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_557),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_657),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_636),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_614),
.A2(n_295),
.B1(n_294),
.B2(n_291),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_557),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_547),
.A2(n_664),
.B(n_662),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_637),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_679),
.B(n_179),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_571),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_543),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_537),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_628),
.B(n_476),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_573),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_482),
.C(n_405),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_544),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_550),
.B(n_335),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_537),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_638),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_563),
.B(n_516),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_659),
.B(n_194),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_571),
.B(n_582),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_653),
.A2(n_425),
.B1(n_452),
.B2(n_282),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_645),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_588),
.B(n_516),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_538),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_661),
.B(n_195),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_582),
.B(n_552),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_538),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_659),
.B(n_195),
.Y(n_782)
);

NAND3x1_ASAP7_75t_L g783 ( 
.A(n_658),
.B(n_408),
.C(n_404),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_603),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_541),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_547),
.A2(n_503),
.B(n_494),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_552),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_659),
.B(n_645),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_645),
.B(n_266),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_542),
.B(n_266),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_542),
.B(n_590),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_669),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_542),
.B(n_293),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_SL g794 ( 
.A(n_674),
.B(n_348),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_546),
.B(n_199),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_545),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_199),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_650),
.B(n_524),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_642),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_511),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_623),
.B(n_200),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_671),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_602),
.B(n_200),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_612),
.B(n_656),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_587),
.B(n_280),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_587),
.B(n_593),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_587),
.B(n_280),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_573),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_SL g809 ( 
.A(n_642),
.B(n_348),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_545),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_573),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_671),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_542),
.B(n_293),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_630),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_634),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_678),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_680),
.B(n_513),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_580),
.B(n_513),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_564),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_575),
.B(n_343),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_580),
.B(n_513),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_595),
.B(n_503),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_576),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_564),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_565),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_576),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_575),
.B(n_343),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_565),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_572),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_575),
.B(n_345),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_572),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_595),
.B(n_508),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_579),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_593),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_682),
.Y(n_835)
);

AO22x1_ASAP7_75t_L g836 ( 
.A1(n_684),
.A2(n_643),
.B1(n_632),
.B2(n_349),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_682),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_710),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_774),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_694),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_684),
.B(n_632),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_714),
.B(n_660),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_714),
.B(n_660),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_718),
.B(n_576),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_699),
.A2(n_664),
.B(n_655),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_710),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_741),
.B(n_524),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_693),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_693),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_724),
.B(n_581),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_716),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_720),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_706),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_533),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_712),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_707),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_697),
.B(n_579),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_707),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_721),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_665),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_776),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_681),
.B(n_533),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_721),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_733),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_733),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_691),
.B(n_542),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_720),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_826),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_735),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_691),
.A2(n_667),
.B1(n_665),
.B2(n_616),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_823),
.B(n_634),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_735),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_R g875 ( 
.A(n_809),
.B(n_601),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_736),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_692),
.A2(n_665),
.B1(n_667),
.B2(n_349),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_737),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_765),
.B(n_589),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_698),
.B(n_560),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_688),
.B(n_411),
.Y(n_882)
);

AO22x1_ASAP7_75t_L g883 ( 
.A1(n_767),
.A2(n_269),
.B1(n_279),
.B2(n_262),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_765),
.B(n_589),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_685),
.Y(n_885)
);

INVx5_ASAP7_75t_L g886 ( 
.A(n_776),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_712),
.B(n_592),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_737),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_762),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_739),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_739),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_729),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_756),
.B(n_581),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_683),
.B(n_695),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_745),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_745),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_776),
.B(n_605),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_695),
.B(n_701),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_599),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_752),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_744),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_719),
.B(n_539),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_760),
.B(n_599),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_740),
.B(n_621),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_690),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_743),
.A2(n_804),
.B1(n_788),
.B2(n_746),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_826),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_792),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_787),
.A2(n_667),
.B1(n_630),
.B2(n_293),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_802),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_771),
.B(n_590),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_812),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_799),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_686),
.B(n_539),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_SL g915 ( 
.A1(n_769),
.A2(n_177),
.B1(n_316),
.B2(n_323),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_816),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_685),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_702),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_763),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_758),
.B(n_412),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_768),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_689),
.B(n_621),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_784),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_703),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_705),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_815),
.Y(n_926)
);

AND2x4_ASAP7_75t_SL g927 ( 
.A(n_754),
.B(n_601),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_713),
.B(n_622),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_725),
.B(n_622),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_764),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_798),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_804),
.B(n_625),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_754),
.B(n_213),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_746),
.A2(n_553),
.B1(n_670),
.B2(n_577),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_704),
.B(n_625),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_770),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_779),
.A2(n_795),
.B1(n_696),
.B2(n_797),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_723),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_798),
.B(n_773),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_770),
.Y(n_940)
);

AND2x2_ASAP7_75t_SL g941 ( 
.A(n_700),
.B(n_293),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_778),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_820),
.B(n_626),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_814),
.B(n_413),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_779),
.A2(n_553),
.B1(n_670),
.B2(n_577),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_820),
.B(n_827),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_758),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_827),
.B(n_629),
.Y(n_948)
);

AND2x6_ASAP7_75t_L g949 ( 
.A(n_811),
.B(n_605),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_811),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_SL g951 ( 
.A(n_794),
.B(n_287),
.C(n_285),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_811),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_700),
.A2(n_243),
.B1(n_242),
.B2(n_304),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_830),
.B(n_795),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_782),
.B(n_418),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_727),
.B(n_233),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_715),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_830),
.B(n_629),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_508),
.B(n_509),
.C(n_289),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_781),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_775),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_803),
.B(n_631),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_785),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_803),
.B(n_421),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_727),
.A2(n_277),
.B1(n_241),
.B2(n_244),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_732),
.B(n_577),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_766),
.B(n_631),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_730),
.B(n_422),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_796),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_758),
.B(n_424),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_810),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_808),
.B(n_640),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_757),
.A2(n_267),
.B1(n_272),
.B2(n_350),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_759),
.B(n_672),
.Y(n_974)
);

AO22x1_ASAP7_75t_L g975 ( 
.A1(n_801),
.A2(n_321),
.B1(n_326),
.B2(n_300),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_709),
.B(n_672),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_711),
.B(n_672),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_810),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_687),
.A2(n_509),
.B(n_313),
.C(n_354),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_717),
.B(n_664),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_824),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_824),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_SL g983 ( 
.A(n_805),
.B(n_352),
.C(n_345),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_828),
.B(n_640),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_722),
.B(n_573),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_807),
.B(n_439),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_833),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_806),
.Y(n_988)
);

AO22x1_ASAP7_75t_L g989 ( 
.A1(n_783),
.A2(n_302),
.B1(n_320),
.B2(n_306),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_726),
.B(n_553),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_772),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_819),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_777),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_825),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_789),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_947),
.B(n_748),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_SL g997 ( 
.A(n_961),
.B(n_315),
.C(n_310),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_855),
.B(n_761),
.Y(n_998)
);

BUFx4_ASAP7_75t_SL g999 ( 
.A(n_852),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_861),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_839),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_941),
.A2(n_747),
.B1(n_749),
.B2(n_731),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_886),
.A2(n_786),
.B(n_708),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_855),
.B(n_728),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_861),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_SL g1007 ( 
.A(n_983),
.B(n_333),
.C(n_319),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_937),
.A2(n_753),
.B1(n_750),
.B2(n_738),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_941),
.A2(n_956),
.B1(n_894),
.B2(n_939),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_886),
.B(n_829),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_835),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_841),
.B(n_338),
.C(n_337),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_834),
.B(n_439),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_886),
.A2(n_946),
.B(n_943),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_846),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_889),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_842),
.A2(n_329),
.B(n_346),
.C(n_299),
.Y(n_1017)
);

AND2x2_ASAP7_75t_SL g1018 ( 
.A(n_953),
.B(n_336),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_948),
.A2(n_791),
.B(n_818),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_958),
.A2(n_791),
.B(n_821),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_841),
.A2(n_358),
.B1(n_359),
.B2(n_352),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_922),
.A2(n_832),
.B(n_822),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_898),
.B(n_831),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_906),
.A2(n_843),
.B(n_966),
.C(n_965),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_964),
.B(n_800),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_938),
.B(n_817),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_953),
.A2(n_340),
.B1(n_342),
.B2(n_790),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_944),
.B(n_790),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_859),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_861),
.B(n_793),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_889),
.B(n_838),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_840),
.B(n_203),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_965),
.A2(n_813),
.B1(n_793),
.B2(n_655),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_879),
.A2(n_652),
.B(n_648),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_931),
.B(n_641),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_931),
.B(n_649),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_859),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_884),
.A2(n_652),
.B(n_648),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_846),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_947),
.B(n_813),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_845),
.A2(n_619),
.B(n_609),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_864),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_881),
.B(n_316),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_867),
.Y(n_1044)
);

CKINVDCx6p67_ASAP7_75t_R g1045 ( 
.A(n_885),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_983),
.A2(n_663),
.B(n_649),
.C(n_673),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_861),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_904),
.A2(n_608),
.B(n_583),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_844),
.B(n_598),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_844),
.B(n_646),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_885),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_850),
.B(n_646),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_870),
.Y(n_1053)
);

BUFx5_ASAP7_75t_L g1054 ( 
.A(n_897),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_918),
.A2(n_673),
.B(n_668),
.C(n_609),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_868),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_957),
.A2(n_210),
.B1(n_357),
.B2(n_356),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_967),
.A2(n_608),
.B(n_652),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_850),
.B(n_893),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_866),
.A2(n_980),
.B(n_977),
.C(n_976),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_901),
.B(n_887),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_991),
.B(n_668),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_993),
.B(n_610),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_918),
.A2(n_610),
.B(n_619),
.C(n_535),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_924),
.B(n_677),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_869),
.B(n_204),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_870),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_SL g1069 ( 
.A1(n_956),
.A2(n_316),
.B1(n_323),
.B2(n_330),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_871),
.A2(n_677),
.B1(n_676),
.B2(n_651),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_917),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_925),
.B(n_677),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_926),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_966),
.A2(n_676),
.B(n_646),
.C(n_651),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_939),
.A2(n_676),
.B(n_651),
.C(n_298),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_847),
.B(n_208),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_995),
.A2(n_296),
.B(n_216),
.C(n_217),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_972),
.A2(n_652),
.B(n_648),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_950),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_875),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_935),
.A2(n_491),
.B(n_505),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_907),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_848),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_836),
.B(n_219),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_902),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_848),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_986),
.A2(n_535),
.B(n_475),
.C(n_505),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_988),
.A2(n_919),
.B1(n_923),
.B2(n_921),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_927),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_920),
.B(n_583),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_873),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_980),
.A2(n_652),
.B(n_648),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_875),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_908),
.A2(n_322),
.B(n_235),
.C(n_249),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_932),
.A2(n_608),
.B(n_583),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_910),
.A2(n_325),
.B(n_251),
.C(n_255),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_915),
.A2(n_317),
.B(n_257),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_912),
.B(n_535),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_916),
.B(n_224),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_876),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_913),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_962),
.A2(n_985),
.B(n_928),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_847),
.B(n_260),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_955),
.A2(n_332),
.B(n_270),
.C(n_273),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_915),
.B(n_264),
.C(n_275),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_985),
.A2(n_532),
.B(n_521),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_955),
.A2(n_278),
.B1(n_284),
.B2(n_286),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_876),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_914),
.B(n_323),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_973),
.A2(n_536),
.B(n_521),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_974),
.A2(n_977),
.B(n_976),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_920),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_984),
.A2(n_475),
.B(n_521),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_950),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_857),
.A2(n_532),
.B(n_521),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_890),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_968),
.A2(n_505),
.B(n_475),
.C(n_536),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_890),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_854),
.B(n_330),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_849),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_900),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_900),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_SL g1123 ( 
.A1(n_990),
.A2(n_475),
.B(n_505),
.C(n_330),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_871),
.A2(n_505),
.B1(n_536),
.B2(n_532),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_968),
.B(n_862),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_849),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_909),
.A2(n_536),
.B1(n_532),
.B2(n_475),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_837),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_882),
.A2(n_491),
.B1(n_536),
.B2(n_470),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_909),
.B(n_470),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_SL g1131 ( 
.A1(n_877),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_877),
.B(n_462),
.Y(n_1132)
);

BUFx4_ASAP7_75t_SL g1133 ( 
.A(n_920),
.Y(n_1133)
);

AO32x2_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_951),
.A3(n_883),
.B1(n_860),
.B2(n_973),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1001),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1024),
.A2(n_903),
.B(n_899),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1128),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1102),
.A2(n_1020),
.B(n_1019),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1025),
.B(n_882),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_927),
.Y(n_1140)
);

NAND2x1_ASAP7_75t_L g1141 ( 
.A(n_1006),
.B(n_897),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1062),
.B(n_929),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1011),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1074),
.A2(n_856),
.B(n_853),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_1031),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1022),
.A2(n_911),
.B(n_945),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1026),
.B(n_992),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1015),
.B(n_970),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1037),
.Y(n_1149)
);

AO32x2_ASAP7_75t_L g1150 ( 
.A1(n_1003),
.A2(n_951),
.A3(n_860),
.B1(n_975),
.B2(n_895),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1003),
.A2(n_878),
.B(n_896),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1109),
.A2(n_933),
.B(n_863),
.C(n_865),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_1041),
.A2(n_888),
.B(n_891),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1008),
.A2(n_874),
.A3(n_858),
.B(n_987),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1005),
.B(n_880),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_L g1156 ( 
.A(n_996),
.B(n_905),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1125),
.B(n_880),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1009),
.A2(n_892),
.B1(n_934),
.B2(n_994),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1042),
.Y(n_1159)
);

NAND3x1_ASAP7_75t_L g1160 ( 
.A(n_1012),
.B(n_989),
.C(n_872),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_998),
.A2(n_860),
.B1(n_952),
.B2(n_963),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1088),
.B(n_1018),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1017),
.A2(n_959),
.B(n_979),
.C(n_981),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1105),
.A2(n_960),
.B(n_940),
.C(n_978),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1069),
.B(n_969),
.C(n_942),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1044),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1028),
.B(n_970),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1061),
.A2(n_936),
.B(n_930),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1007),
.A2(n_971),
.B(n_982),
.C(n_963),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1034),
.A2(n_982),
.B(n_897),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1089),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1038),
.A2(n_1048),
.B(n_1059),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1106),
.A2(n_952),
.B(n_897),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1085),
.B(n_8),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1078),
.A2(n_897),
.B(n_949),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1084),
.A2(n_949),
.B(n_470),
.C(n_467),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1095),
.A2(n_949),
.B(n_491),
.Y(n_1177)
);

BUFx2_ASAP7_75t_R g1178 ( 
.A(n_1051),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1043),
.B(n_949),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1097),
.A2(n_462),
.B(n_467),
.C(n_13),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1119),
.B(n_10),
.C(n_11),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1132),
.A2(n_491),
.B(n_61),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1033),
.A2(n_1075),
.A3(n_1117),
.B(n_1124),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1085),
.B(n_467),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1023),
.B(n_10),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1016),
.B(n_467),
.Y(n_1186)
);

BUFx10_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1041),
.A2(n_171),
.B(n_166),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_1082),
.B(n_13),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_996),
.A2(n_1049),
.B1(n_1050),
.B2(n_1052),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1115),
.A2(n_1081),
.B(n_1098),
.Y(n_1191)
);

AO22x2_ASAP7_75t_L g1192 ( 
.A1(n_1033),
.A2(n_14),
.B1(n_19),
.B2(n_21),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1055),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_996),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1063),
.B(n_30),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1039),
.B(n_32),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1055),
.B(n_118),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1046),
.A2(n_1065),
.B(n_1056),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1087),
.A2(n_90),
.B(n_81),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1124),
.A2(n_32),
.A3(n_37),
.B(n_38),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1002),
.B(n_37),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1053),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1071),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1029),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1104),
.A2(n_1094),
.B(n_1096),
.C(n_1077),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1073),
.B(n_39),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_1090),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1080),
.B(n_41),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1071),
.B(n_74),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_R g1210 ( 
.A(n_1093),
.B(n_71),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1032),
.B(n_42),
.C(n_44),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1099),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_R g1213 ( 
.A(n_1112),
.B(n_70),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1070),
.A2(n_62),
.B(n_47),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1057),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1130),
.A2(n_45),
.B(n_48),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_51),
.B(n_52),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1101),
.B(n_51),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1035),
.A2(n_53),
.B(n_54),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1057),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1036),
.A2(n_54),
.B(n_58),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1127),
.A2(n_1129),
.B(n_1110),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_1027),
.A2(n_1127),
.A3(n_1123),
.B1(n_1021),
.B2(n_1058),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1027),
.A2(n_1121),
.A3(n_1068),
.B(n_1108),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1103),
.B(n_1064),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1091),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1071),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1118),
.A2(n_1072),
.B(n_1066),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1010),
.A2(n_1122),
.B(n_1100),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1010),
.A2(n_1116),
.B(n_1030),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1076),
.A2(n_1040),
.B(n_1126),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1030),
.A2(n_1083),
.B(n_1126),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1086),
.A2(n_1120),
.B(n_1047),
.C(n_1000),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1079),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1067),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1079),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1045),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_1090),
.B(n_1114),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1054),
.A2(n_1107),
.B(n_1114),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_997),
.A2(n_1054),
.B(n_1114),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_1133),
.A2(n_1090),
.B1(n_999),
.B2(n_1054),
.Y(n_1241)
);

NOR3xp33_ASAP7_75t_SL g1242 ( 
.A(n_1054),
.B(n_593),
.C(n_632),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1009),
.A2(n_937),
.B1(n_954),
.B2(n_691),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1113),
.A2(n_1092),
.B(n_1111),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1060),
.B(n_684),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1109),
.A2(n_954),
.B(n_946),
.C(n_684),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1109),
.A2(n_684),
.B(n_714),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1055),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1024),
.A2(n_776),
.B(n_954),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1001),
.Y(n_1250)
);

AOI221x1_ASAP7_75t_L g1251 ( 
.A1(n_1024),
.A2(n_954),
.B1(n_946),
.B2(n_1109),
.C(n_1014),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1089),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1060),
.B(n_684),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1004),
.A2(n_946),
.B(n_886),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1128),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1109),
.A2(n_769),
.B1(n_692),
.B2(n_937),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1015),
.B(n_846),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1060),
.B(n_855),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

CKINVDCx8_ASAP7_75t_R g1261 ( 
.A(n_1055),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1245),
.B(n_1253),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1214),
.A2(n_1192),
.B1(n_1247),
.B2(n_1243),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1143),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1261),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1258),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1207),
.B(n_1156),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1207),
.B(n_1156),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1142),
.B(n_1162),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1259),
.B(n_1155),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1251),
.A2(n_1172),
.A3(n_1176),
.B(n_1146),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1204),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1254),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1147),
.B(n_1139),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1258),
.B(n_1203),
.Y(n_1275)
);

NOR2x1_ASAP7_75t_SL g1276 ( 
.A(n_1207),
.B(n_1190),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1214),
.A2(n_1246),
.B(n_1222),
.C(n_1217),
.Y(n_1277)
);

AOI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1192),
.A2(n_1136),
.B(n_1158),
.Y(n_1278)
);

INVx3_ASAP7_75t_SL g1279 ( 
.A(n_1171),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1148),
.B(n_1227),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1255),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1168),
.A2(n_1163),
.A3(n_1152),
.B(n_1164),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1225),
.B(n_1157),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1249),
.A2(n_1136),
.B(n_1198),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1170),
.A2(n_1173),
.B(n_1177),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1260),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1228),
.A2(n_1199),
.B(n_1188),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1167),
.B(n_1195),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1187),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1222),
.A2(n_1180),
.B1(n_1181),
.B2(n_1256),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1232),
.A2(n_1239),
.B(n_1230),
.Y(n_1291)
);

AOI222xp33_ASAP7_75t_L g1292 ( 
.A1(n_1211),
.A2(n_1189),
.B1(n_1206),
.B2(n_1218),
.C1(n_1201),
.C2(n_1194),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1149),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1231),
.A2(n_1238),
.B(n_1216),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1159),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1166),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1240),
.B(n_1141),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1185),
.A2(n_1174),
.B1(n_1212),
.B2(n_1160),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1205),
.A2(n_1169),
.B(n_1228),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1165),
.A2(n_1219),
.B(n_1221),
.C(n_1161),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1202),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1229),
.A2(n_1144),
.B(n_1191),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1135),
.B(n_1250),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1144),
.A2(n_1191),
.B(n_1153),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1189),
.A2(n_1241),
.B1(n_1182),
.B2(n_1179),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1197),
.A2(n_1209),
.B(n_1242),
.C(n_1134),
.Y(n_1307)
);

BUFx4_ASAP7_75t_SL g1308 ( 
.A(n_1215),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1186),
.A2(n_1184),
.B(n_1134),
.C(n_1236),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1240),
.B(n_1227),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1227),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1224),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1233),
.A2(n_1150),
.B(n_1223),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1248),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1224),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1145),
.B(n_1235),
.Y(n_1316)
);

OAI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1208),
.A2(n_1196),
.B1(n_1237),
.B2(n_1248),
.C(n_1223),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1200),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_SL g1319 ( 
.A(n_1210),
.B(n_1252),
.C(n_1220),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1187),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1193),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1183),
.B(n_1200),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1248),
.A2(n_1209),
.B1(n_1197),
.B2(n_1213),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1193),
.B(n_1200),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1178),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1223),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1227),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1138),
.A2(n_1172),
.B(n_1151),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1258),
.B(n_1203),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1137),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1258),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1151),
.A2(n_1175),
.B(n_1254),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1245),
.B(n_1253),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1258),
.Y(n_1334)
);

AO21x1_ASAP7_75t_L g1335 ( 
.A1(n_1247),
.A2(n_1253),
.B(n_1245),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1147),
.B(n_840),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1245),
.B(n_1253),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1234),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1138),
.A2(n_1249),
.B(n_946),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1175),
.A2(n_1113),
.B(n_1244),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1138),
.A2(n_1172),
.B(n_1151),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1137),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1175),
.A2(n_1113),
.B(n_1244),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1245),
.B(n_1253),
.Y(n_1345)
);

AO22x2_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_1214),
.B1(n_1251),
.B2(n_1190),
.Y(n_1346)
);

BUFx4f_ASAP7_75t_L g1347 ( 
.A(n_1260),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1137),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1137),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1140),
.B(n_1013),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1246),
.A2(n_1247),
.B(n_1253),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_941),
.B2(n_965),
.Y(n_1352)
);

AOI221x1_ASAP7_75t_L g1353 ( 
.A1(n_1247),
.A2(n_1245),
.B1(n_1253),
.B2(n_1192),
.C(n_1214),
.Y(n_1353)
);

INVx4_ASAP7_75t_SL g1354 ( 
.A(n_1200),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1138),
.A2(n_1249),
.B(n_946),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1137),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_1247),
.B2(n_941),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1251),
.A2(n_1172),
.A3(n_1176),
.B(n_1243),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1137),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1245),
.A2(n_941),
.B1(n_1253),
.B2(n_366),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1258),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_961),
.B2(n_841),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1260),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1251),
.A2(n_1138),
.B(n_1172),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1247),
.A2(n_1253),
.B(n_1245),
.C(n_1257),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1137),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1140),
.B(n_1013),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_941),
.B2(n_965),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1137),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1251),
.A2(n_1138),
.B(n_1172),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1260),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_1247),
.B2(n_941),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1175),
.A2(n_1113),
.B(n_1244),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1259),
.B(n_1147),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1207),
.B(n_886),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1265),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1274),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1284),
.A2(n_1304),
.B(n_1302),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1362),
.B(n_1262),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1279),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1284),
.A2(n_1355),
.B(n_1340),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1263),
.A2(n_1277),
.B(n_1278),
.C(n_1351),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1293),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1366),
.A2(n_1352),
.B(n_1369),
.C(n_1263),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1366),
.A2(n_1352),
.B(n_1369),
.C(n_1277),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1303),
.B(n_1288),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1265),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1321),
.Y(n_1391)
);

CKINVDCx6p67_ASAP7_75t_R g1392 ( 
.A(n_1279),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1283),
.B(n_1351),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1360),
.A2(n_1357),
.B1(n_1373),
.B2(n_1337),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1357),
.B(n_1373),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1331),
.B(n_1334),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1278),
.A2(n_1335),
.B(n_1299),
.C(n_1290),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1308),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1316),
.B(n_1319),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1361),
.B(n_1266),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1328),
.A2(n_1342),
.B(n_1273),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1290),
.A2(n_1313),
.B(n_1305),
.C(n_1307),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1262),
.B(n_1333),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1280),
.B(n_1272),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1323),
.A2(n_1376),
.B(n_1353),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1333),
.B(n_1337),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1298),
.A2(n_1345),
.B(n_1300),
.C(n_1292),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1295),
.B(n_1296),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1360),
.A2(n_1345),
.B1(n_1336),
.B2(n_1323),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1317),
.A2(n_1346),
.B1(n_1316),
.B2(n_1325),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1292),
.A2(n_1294),
.B(n_1319),
.C(n_1309),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1309),
.A2(n_1356),
.B(n_1339),
.C(n_1343),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1281),
.A2(n_1359),
.B(n_1349),
.C(n_1348),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1275),
.B(n_1329),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1326),
.A2(n_1318),
.B(n_1315),
.C(n_1312),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1330),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1346),
.B(n_1306),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1346),
.B(n_1301),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1276),
.B(n_1367),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1321),
.A2(n_1267),
.B1(n_1268),
.B2(n_1370),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1365),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1338),
.B(n_1314),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1321),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1338),
.B(n_1314),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1341),
.A2(n_1344),
.B(n_1374),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1364),
.B(n_1371),
.Y(n_1426)
);

OA22x2_ASAP7_75t_L g1427 ( 
.A1(n_1289),
.A2(n_1320),
.B1(n_1291),
.B2(n_1285),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1267),
.A2(n_1268),
.B(n_1310),
.C(n_1371),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1358),
.B(n_1354),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1311),
.Y(n_1430)
);

INVx6_ASAP7_75t_SL g1431 ( 
.A(n_1308),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1347),
.A2(n_1376),
.B1(n_1297),
.B2(n_1327),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1311),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1314),
.B(n_1327),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1327),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1347),
.A2(n_1297),
.B1(n_1287),
.B2(n_1286),
.Y(n_1436)
);

CKINVDCx12_ASAP7_75t_R g1437 ( 
.A(n_1372),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1358),
.B(n_1271),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1358),
.B(n_1282),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1287),
.A2(n_1363),
.B1(n_1332),
.B2(n_1282),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1366),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1444)
);

INVx5_ASAP7_75t_L g1445 ( 
.A(n_1324),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1340),
.A2(n_1355),
.B(n_1284),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1263),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1360),
.A2(n_1245),
.B1(n_1253),
.B2(n_1362),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1366),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1450)
);

O2A1O1Ixp5_ASAP7_75t_L g1451 ( 
.A1(n_1263),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1265),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1266),
.B(n_1280),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1366),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1264),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1360),
.A2(n_1245),
.B1(n_1253),
.B2(n_1362),
.Y(n_1458)
);

OAI211xp5_ASAP7_75t_L g1459 ( 
.A1(n_1360),
.A2(n_1245),
.B(n_1253),
.C(n_1247),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1340),
.A2(n_1355),
.B(n_1284),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1263),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1360),
.A2(n_1245),
.B1(n_1253),
.B2(n_1362),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1274),
.B(n_1375),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1324),
.A2(n_954),
.B(n_1322),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1360),
.A2(n_1245),
.B1(n_1253),
.B2(n_1362),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_SL g1468 ( 
.A1(n_1324),
.A2(n_954),
.B(n_1322),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1366),
.A2(n_1247),
.B(n_1253),
.C(n_1245),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1360),
.A2(n_1245),
.B1(n_1253),
.B2(n_1362),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1415),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1379),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1421),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1380),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1456),
.A2(n_1459),
.B1(n_1441),
.B2(n_1470),
.C(n_1448),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1417),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1378),
.B(n_1442),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1447),
.A2(n_1463),
.B(n_1451),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1442),
.B(n_1444),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1418),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1458),
.A2(n_1467),
.B1(n_1464),
.B2(n_1394),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1418),
.B(n_1438),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1446),
.A2(n_1462),
.B(n_1401),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1485)
);

OR2x6_ASAP7_75t_L g1486 ( 
.A(n_1446),
.B(n_1462),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1426),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1380),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1384),
.B(n_1389),
.Y(n_1489)
);

OAI321xp33_ASAP7_75t_L g1490 ( 
.A1(n_1459),
.A2(n_1407),
.A3(n_1449),
.B1(n_1469),
.B2(n_1387),
.C(n_1388),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1386),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1445),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1384),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1419),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1393),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1430),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1416),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1427),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1385),
.A2(n_1402),
.B(n_1397),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1430),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1425),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1440),
.A2(n_1388),
.B(n_1395),
.Y(n_1502)
);

INVxp33_ASAP7_75t_L g1503 ( 
.A(n_1396),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1419),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1413),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1413),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1449),
.A2(n_1469),
.B(n_1407),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1412),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1428),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1408),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1381),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1395),
.A2(n_1387),
.B(n_1393),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1411),
.A2(n_1409),
.B(n_1436),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1412),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1427),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1382),
.A2(n_1410),
.B1(n_1399),
.B2(n_1392),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1443),
.A2(n_1450),
.B1(n_1452),
.B2(n_1461),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1420),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1403),
.A2(n_1406),
.B1(n_1460),
.B2(n_1437),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1405),
.A2(n_1468),
.B(n_1466),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_L g1521 ( 
.A(n_1432),
.B(n_1457),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1501),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1497),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1404),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1489),
.B(n_1406),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1501),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1486),
.B(n_1434),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1486),
.B(n_1422),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1424),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1476),
.B(n_1403),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1493),
.B(n_1484),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1489),
.B(n_1435),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1471),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1476),
.B(n_1400),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_R g1538 ( 
.A(n_1496),
.B(n_1398),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1473),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1484),
.B(n_1414),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1480),
.B(n_1433),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1492),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1480),
.B(n_1512),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1484),
.B(n_1455),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1485),
.B(n_1391),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1474),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1526),
.A2(n_1475),
.B1(n_1482),
.B2(n_1490),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1525),
.A2(n_1507),
.B1(n_1512),
.B2(n_1478),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1523),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1535),
.B(n_1498),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_R g1551 ( 
.A(n_1545),
.B(n_1383),
.Y(n_1551)
);

AOI33xp33_ASAP7_75t_L g1552 ( 
.A1(n_1533),
.A2(n_1516),
.A3(n_1517),
.B1(n_1519),
.B2(n_1483),
.B3(n_1505),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1523),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1523),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1524),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1525),
.A2(n_1512),
.B1(n_1478),
.B2(n_1502),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1522),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1534),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1536),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1535),
.B(n_1515),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1534),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1542),
.B(n_1494),
.Y(n_1562)
);

OR2x6_ASAP7_75t_SL g1563 ( 
.A(n_1526),
.B(n_1495),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1535),
.B(n_1515),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1538),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

INVx5_ASAP7_75t_L g1569 ( 
.A(n_1542),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1543),
.A2(n_1490),
.B1(n_1513),
.B2(n_1509),
.C(n_1504),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1525),
.A2(n_1512),
.B1(n_1502),
.B2(n_1518),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1538),
.Y(n_1572)
);

AOI31xp33_ASAP7_75t_L g1573 ( 
.A1(n_1530),
.A2(n_1519),
.A3(n_1503),
.B(n_1531),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_R g1574 ( 
.A(n_1542),
.B(n_1431),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1545),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1543),
.A2(n_1513),
.B1(n_1472),
.B2(n_1511),
.C(n_1506),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1534),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1525),
.A2(n_1502),
.B1(n_1518),
.B2(n_1499),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1546),
.A2(n_1474),
.B(n_1488),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1471),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1545),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1530),
.A2(n_1502),
.B1(n_1499),
.B2(n_1520),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1530),
.A2(n_1520),
.B1(n_1499),
.B2(n_1506),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1532),
.A2(n_1495),
.B1(n_1477),
.B2(n_1479),
.C(n_1481),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1542),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1529),
.B(n_1494),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1529),
.B(n_1494),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1533),
.B(n_1499),
.C(n_1521),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1527),
.Y(n_1590)
);

NOR4xp25_ASAP7_75t_SL g1591 ( 
.A(n_1539),
.B(n_1508),
.C(n_1514),
.D(n_1505),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1541),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1579),
.A2(n_1589),
.B(n_1533),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1551),
.B(n_1492),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1567),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1549),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1563),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1580),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1547),
.A2(n_1521),
.B(n_1514),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1563),
.B(n_1544),
.Y(n_1603)
);

INVx4_ASAP7_75t_SL g1604 ( 
.A(n_1562),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1553),
.Y(n_1606)
);

AND2x6_ASAP7_75t_SL g1607 ( 
.A(n_1562),
.B(n_1431),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1550),
.B(n_1544),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1570),
.A2(n_1508),
.B(n_1533),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1550),
.B(n_1544),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1569),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1569),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

INVx4_ASAP7_75t_SL g1616 ( 
.A(n_1562),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1590),
.Y(n_1617)
);

AND2x4_ASAP7_75t_SL g1618 ( 
.A(n_1585),
.B(n_1492),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1554),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1546),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1576),
.A2(n_1544),
.B(n_1540),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1569),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1555),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1555),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1568),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1560),
.B(n_1540),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1624),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1594),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1600),
.B(n_1560),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1611),
.A2(n_1548),
.B1(n_1556),
.B2(n_1571),
.C(n_1578),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1594),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1597),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1611),
.B(n_1552),
.C(n_1565),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1564),
.Y(n_1634)
);

NAND2x1_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1573),
.Y(n_1635)
);

NAND2x1_ASAP7_75t_L g1636 ( 
.A(n_1614),
.B(n_1613),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1564),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1587),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1594),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1587),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1602),
.B(n_1593),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1646)
);

NAND2x1_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1575),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1599),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1583),
.C(n_1582),
.D(n_1540),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1605),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1605),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1591),
.C(n_1540),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1624),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1604),
.B(n_1616),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1603),
.B(n_1575),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1607),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1614),
.B(n_1569),
.C(n_1491),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1616),
.B(n_1558),
.Y(n_1665)
);

AND2x4_ASAP7_75t_SL g1666 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1605),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1616),
.B(n_1561),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1606),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1596),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1616),
.B(n_1577),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1603),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1601),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1661),
.B(n_1616),
.Y(n_1675)
);

AND3x1_ASAP7_75t_L g1676 ( 
.A(n_1661),
.B(n_1622),
.C(n_1613),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1614),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1616),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1663),
.B(n_1645),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_L g1680 ( 
.A(n_1646),
.B(n_1572),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1635),
.A2(n_1614),
.B1(n_1622),
.B2(n_1613),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1628),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1627),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1635),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1650),
.B(n_1601),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1628),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1636),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1632),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_1633),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1631),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1608),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1377),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1629),
.B(n_1616),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1634),
.B(n_1626),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1662),
.B(n_1655),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1636),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1659),
.B(n_1609),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1631),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1609),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1640),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1627),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1666),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1664),
.B(n_1610),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1640),
.B(n_1581),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1641),
.B(n_1643),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1642),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1688),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1682),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1679),
.B(n_1693),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1709),
.B(n_1666),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1673),
.B(n_1609),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1678),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1686),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1690),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1674),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1612),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1702),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1709),
.B(n_1641),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1687),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1694),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1695),
.B(n_1642),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1704),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1687),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1697),
.B(n_1647),
.C(n_1614),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1695),
.B(n_1648),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1698),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1706),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1677),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1674),
.B(n_1648),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1737),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1681),
.B(n_1680),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1737),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1711),
.A2(n_1680),
.B1(n_1694),
.B2(n_1676),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1731),
.A2(n_1701),
.B1(n_1699),
.B2(n_1707),
.C(n_1677),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1720),
.A2(n_1707),
.B1(n_1614),
.B2(n_1685),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1730),
.Y(n_1746)
);

OAI322xp33_ASAP7_75t_L g1747 ( 
.A1(n_1735),
.A2(n_1685),
.A3(n_1696),
.B1(n_1691),
.B2(n_1703),
.C1(n_1708),
.C2(n_1683),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1714),
.A2(n_1675),
.B1(n_1637),
.B2(n_1656),
.Y(n_1748)
);

OAI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1716),
.A2(n_1691),
.B(n_1698),
.Y(n_1749)
);

OAI322xp33_ASAP7_75t_L g1750 ( 
.A1(n_1721),
.A2(n_1708),
.A3(n_1705),
.B1(n_1683),
.B2(n_1652),
.C1(n_1657),
.C2(n_1658),
.Y(n_1750)
);

AOI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1713),
.A2(n_1700),
.B1(n_1665),
.B2(n_1672),
.C1(n_1668),
.C2(n_1651),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1656),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1712),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1730),
.Y(n_1754)
);

AOI222xp33_ASAP7_75t_L g1755 ( 
.A1(n_1715),
.A2(n_1700),
.B1(n_1668),
.B2(n_1665),
.C1(n_1651),
.C2(n_1637),
.Y(n_1755)
);

AOI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1736),
.A2(n_1622),
.B(n_1613),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1723),
.A2(n_1622),
.B(n_1651),
.Y(n_1757)
);

OR4x1_ASAP7_75t_L g1758 ( 
.A(n_1712),
.B(n_1657),
.C(n_1669),
.D(n_1667),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1740),
.A2(n_1734),
.B1(n_1729),
.B2(n_1725),
.C(n_1723),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1739),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1743),
.B(n_1734),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1746),
.B(n_1725),
.Y(n_1762)
);

INVxp67_ASAP7_75t_SL g1763 ( 
.A(n_1745),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1738),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1744),
.A2(n_1651),
.B1(n_1729),
.B2(n_1595),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1754),
.B(n_1717),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1749),
.B(n_1717),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1753),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1748),
.B(n_1727),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1766),
.A2(n_1742),
.B(n_1744),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1763),
.A2(n_1745),
.B(n_1756),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1759),
.A2(n_1747),
.B1(n_1750),
.B2(n_1758),
.C(n_1752),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1757),
.Y(n_1774)
);

AOI211x1_ASAP7_75t_SL g1775 ( 
.A1(n_1768),
.A2(n_1767),
.B(n_1705),
.C(n_1770),
.Y(n_1775)
);

O2A1O1Ixp5_ASAP7_75t_L g1776 ( 
.A1(n_1762),
.A2(n_1728),
.B(n_1718),
.C(n_1733),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1761),
.A2(n_1751),
.B1(n_1755),
.B2(n_1770),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1762),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1760),
.A2(n_1733),
.B(n_1728),
.C(n_1722),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1764),
.B(n_1761),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1760),
.A2(n_1722),
.B1(n_1718),
.B2(n_1732),
.C(n_1727),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1778),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1780),
.Y(n_1783)
);

AO22x1_ASAP7_75t_SL g1784 ( 
.A1(n_1775),
.A2(n_1769),
.B1(n_1620),
.B2(n_1669),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1777),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1776),
.Y(n_1786)
);

AO22x2_ASAP7_75t_L g1787 ( 
.A1(n_1772),
.A2(n_1732),
.B1(n_1658),
.B2(n_1667),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1779),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1781),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1782),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1785),
.B(n_1773),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1786),
.B(n_1774),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1788),
.B(n_1771),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1783),
.B(n_1612),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1787),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1789),
.B(n_1595),
.C(n_1671),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1791),
.A2(n_1784),
.B(n_1787),
.C(n_1390),
.Y(n_1797)
);

BUFx12f_ASAP7_75t_L g1798 ( 
.A(n_1790),
.Y(n_1798)
);

AOI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1792),
.A2(n_1793),
.B(n_1795),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1794),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1796),
.A2(n_1784),
.B1(n_1595),
.B2(n_1454),
.C(n_1671),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1794),
.B(n_1620),
.Y(n_1802)
);

OAI311xp33_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1652),
.A3(n_1592),
.B1(n_1612),
.C1(n_1541),
.Y(n_1803)
);

NAND5xp2_ASAP7_75t_L g1804 ( 
.A(n_1797),
.B(n_1574),
.C(n_1529),
.D(n_1531),
.E(n_1530),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1800),
.B(n_1639),
.Y(n_1805)
);

NAND4xp25_ASAP7_75t_L g1806 ( 
.A(n_1799),
.B(n_1423),
.C(n_1586),
.D(n_1620),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1802),
.Y(n_1807)
);

AOI322xp5_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1798),
.A3(n_1805),
.B1(n_1806),
.B2(n_1803),
.C1(n_1625),
.C2(n_1639),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1808),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1808),
.A2(n_1660),
.B1(n_1644),
.B2(n_1595),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1809),
.Y(n_1811)
);

AOI22x1_ASAP7_75t_L g1812 ( 
.A1(n_1810),
.A2(n_1660),
.B1(n_1644),
.B2(n_1625),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1620),
.B1(n_1618),
.B2(n_1623),
.C(n_1619),
.Y(n_1813)
);

INVx4_ASAP7_75t_L g1814 ( 
.A(n_1812),
.Y(n_1814)
);

XNOR2xp5_ASAP7_75t_L g1815 ( 
.A(n_1813),
.B(n_1618),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1814),
.B1(n_1620),
.B2(n_1595),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1816),
.B(n_1620),
.Y(n_1817)
);

AOI22x1_ASAP7_75t_L g1818 ( 
.A1(n_1817),
.A2(n_1598),
.B1(n_1617),
.B2(n_1615),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1595),
.B1(n_1618),
.B2(n_1596),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1574),
.B(n_1496),
.C(n_1500),
.Y(n_1820)
);


endmodule