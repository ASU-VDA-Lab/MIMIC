module fake_netlist_1_3175_n_557 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_557);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_557;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_70), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_47), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_31), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_2), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_58), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_71), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_53), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_68), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_21), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_51), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_5), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_10), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_76), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_41), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_54), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_28), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_46), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_43), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_35), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_89), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_85), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_85), .Y(n_115) );
NAND2xp33_ASAP7_75t_L g116 ( .A(n_91), .B(n_30), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_86), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_111), .B(n_0), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_78), .Y(n_121) );
INVx2_ASAP7_75t_SL g122 ( .A(n_90), .Y(n_122) );
AND2x6_ASAP7_75t_L g123 ( .A(n_87), .B(n_27), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_90), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_98), .B(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_99), .Y(n_129) );
AND3x2_ASAP7_75t_L g130 ( .A(n_112), .B(n_1), .C(n_2), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_99), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_83), .B(n_3), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
INVx5_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_105), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_125), .B(n_110), .Y(n_138) );
OAI22xp33_ASAP7_75t_L g139 ( .A1(n_127), .A2(n_79), .B1(n_93), .B2(n_101), .Y(n_139) );
NOR2xp33_ASAP7_75t_SL g140 ( .A(n_123), .B(n_79), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_114), .B(n_93), .Y(n_141) );
INVx6_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_129), .B(n_114), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_116), .B(n_95), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_115), .B(n_101), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_123), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_120), .B(n_95), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_115), .B(n_109), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_137), .A2(n_108), .B1(n_107), .B2(n_104), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_117), .B(n_103), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_117), .B(n_88), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
AND3x1_ASAP7_75t_L g164 ( .A(n_131), .B(n_100), .C(n_97), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_132), .B(n_96), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_163), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_141), .B(n_118), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_164), .B(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_143), .B(n_118), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_138), .B(n_132), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_139), .B(n_128), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_149), .B(n_120), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_147), .B(n_133), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_154), .B(n_120), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_154), .B(n_120), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_147), .B(n_122), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_140), .A2(n_123), .B1(n_135), .B2(n_122), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_156), .B(n_121), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_147), .B(n_113), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_152), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_160), .B(n_135), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_161), .B(n_113), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_165), .B(n_123), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_154), .B(n_84), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_167), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_168), .B(n_140), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_171), .B(n_158), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_196), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_198), .A2(n_158), .B(n_148), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_172), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_179), .A2(n_123), .B1(n_158), .B2(n_134), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_186), .A2(n_134), .B(n_126), .C(n_80), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_194), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_169), .B(n_158), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_177), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_181), .A2(n_148), .B(n_145), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
AND3x1_ASAP7_75t_SL g221 ( .A(n_200), .B(n_130), .C(n_82), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_126), .B(n_134), .C(n_92), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_194), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_173), .B(n_148), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_148), .B1(n_94), .B2(n_81), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_188), .B(n_126), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_200), .B(n_148), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_169), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_124), .B(n_148), .C(n_157), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_146), .B(n_145), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_169), .A2(n_142), .B1(n_136), .B2(n_124), .Y(n_232) );
BUFx8_ASAP7_75t_L g233 ( .A(n_175), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_167), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_230), .A2(n_201), .B(n_174), .C(n_180), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_236), .A2(n_192), .B1(n_197), .B2(n_187), .C(n_136), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_230), .A2(n_199), .B(n_195), .C(n_180), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_214), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
NAND2x1p5_ASAP7_75t_L g242 ( .A(n_217), .B(n_177), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_209), .A2(n_199), .B(n_195), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_235), .A2(n_191), .B1(n_193), .B2(n_194), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_214), .Y(n_246) );
AO31x2_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_146), .A3(n_157), .B(n_155), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_208), .B(n_193), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_214), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_207), .A2(n_191), .B(n_182), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_213), .A2(n_162), .B(n_155), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_216), .B(n_177), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_214), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_232), .A2(n_162), .B(n_190), .Y(n_257) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_166), .B(n_190), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_205), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_194), .B1(n_178), .B2(n_183), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_222), .A2(n_185), .B(n_182), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_227), .B(n_177), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_207), .A2(n_124), .B1(n_136), .B2(n_178), .C(n_183), .Y(n_263) );
INVx6_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_226), .B(n_217), .C(n_220), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_238), .A2(n_210), .B1(n_203), .B2(n_233), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_241), .B(n_205), .Y(n_267) );
AOI22xp33_ASAP7_75t_SL g268 ( .A1(n_249), .A2(n_233), .B1(n_210), .B2(n_203), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_254), .A2(n_234), .B1(n_215), .B2(n_211), .Y(n_270) );
OR2x6_ASAP7_75t_SL g271 ( .A(n_244), .B(n_221), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_259), .B(n_211), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_237), .A2(n_212), .B1(n_234), .B2(n_215), .C(n_204), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_248), .B(n_212), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_248), .B(n_225), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_239), .A2(n_224), .B(n_231), .Y(n_279) );
NOR2x1_ASAP7_75t_SL g280 ( .A(n_255), .B(n_223), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_245), .B(n_253), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_262), .A2(n_124), .B1(n_221), .B2(n_136), .C(n_219), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_252), .A2(n_185), .B(n_166), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_250), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_258), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_282), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_282), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_276), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_272), .B(n_257), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_266), .B(n_253), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_286), .Y(n_295) );
INVxp33_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_272), .B(n_257), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_271), .B(n_242), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_285), .A2(n_252), .B(n_261), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_287), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_273), .B(n_246), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_267), .B(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_267), .B(n_246), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_256), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_278), .B(n_256), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
OAI31xp33_ASAP7_75t_L g311 ( .A1(n_296), .A2(n_265), .A3(n_277), .B(n_278), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_309), .B(n_277), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_309), .B(n_284), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_309), .B(n_284), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_303), .B(n_281), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_307), .B(n_276), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_307), .B(n_257), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
NOR2xp33_ASAP7_75t_SL g322 ( .A(n_291), .B(n_282), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_308), .B(n_271), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g324 ( .A(n_297), .B(n_283), .C(n_275), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_307), .B(n_280), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_297), .B(n_257), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_289), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_305), .B(n_280), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_305), .B(n_282), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_305), .B(n_282), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_291), .B(n_250), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_296), .B(n_255), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_306), .B(n_285), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_285), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_306), .B(n_285), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_293), .B(n_247), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_295), .B(n_255), .Y(n_342) );
NAND3xp33_ASAP7_75t_SL g343 ( .A(n_311), .B(n_299), .C(n_291), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_314), .B(n_308), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_337), .B(n_293), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_327), .B(n_291), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_332), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_327), .B(n_295), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_337), .B(n_298), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_327), .B(n_291), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_332), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
AOI211x1_ASAP7_75t_L g354 ( .A1(n_323), .A2(n_298), .B(n_304), .C(n_5), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_314), .B(n_304), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_313), .B(n_304), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_321), .B(n_294), .Y(n_360) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_311), .A2(n_299), .B(n_294), .C(n_302), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_339), .B(n_288), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_339), .B(n_292), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_325), .B(n_289), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_340), .B(n_292), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_340), .B(n_292), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_320), .B(n_301), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_316), .B(n_302), .Y(n_371) );
AND4x1_ASAP7_75t_L g372 ( .A(n_322), .B(n_3), .C(n_4), .D(n_6), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_335), .B(n_302), .Y(n_374) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_329), .B(n_289), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_322), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_324), .B(n_136), .C(n_270), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_324), .B(n_310), .C(n_289), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_320), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_319), .B(n_301), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
INVx6_ASAP7_75t_L g384 ( .A(n_325), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_319), .B(n_289), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_318), .B(n_310), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_310), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_326), .B(n_310), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_367), .B(n_326), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_388), .B(n_341), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_367), .B(n_325), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_381), .B(n_325), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_381), .B(n_328), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
AOI221x1_ASAP7_75t_L g399 ( .A1(n_380), .A2(n_310), .B1(n_335), .B2(n_279), .C(n_334), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_386), .B(n_316), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_388), .B(n_317), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_384), .Y(n_402) );
NOR2xp67_ASAP7_75t_SL g403 ( .A(n_378), .B(n_379), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_344), .B(n_317), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
OAI32xp33_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_336), .A3(n_342), .B1(n_330), .B2(n_333), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_357), .B(n_334), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_345), .B(n_333), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_369), .B(n_335), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_345), .B(n_335), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_387), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_387), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_347), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_350), .B(n_247), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_350), .B(n_247), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_359), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_352), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_352), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_376), .B(n_4), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_358), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_358), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
AND3x1_ASAP7_75t_L g428 ( .A(n_361), .B(n_6), .C(n_7), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_247), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_360), .B(n_8), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_363), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_343), .A2(n_389), .B1(n_371), .B2(n_364), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_365), .B(n_9), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_365), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_364), .A2(n_264), .B1(n_258), .B2(n_240), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_384), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_354), .B(n_263), .C(n_260), .D(n_11), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_366), .B(n_9), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_366), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g441 ( .A(n_374), .B(n_240), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_382), .B(n_389), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_397), .B(n_384), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_420), .B(n_382), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_422), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_397), .B(n_384), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_391), .B(n_385), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_428), .A2(n_375), .B1(n_349), .B2(n_346), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_430), .A2(n_385), .B1(n_364), .B2(n_377), .C(n_159), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
AOI31xp33_ASAP7_75t_L g453 ( .A1(n_433), .A2(n_351), .A3(n_346), .B(n_372), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_391), .B(n_351), .Y(n_454) );
OAI31xp33_ASAP7_75t_L g455 ( .A1(n_438), .A2(n_242), .A3(n_256), .B(n_12), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_433), .B(n_263), .C(n_11), .D(n_12), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_407), .A2(n_258), .B(n_252), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_441), .A2(n_255), .B1(n_264), .B2(n_242), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_414), .B(n_10), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_415), .B(n_13), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_264), .B1(n_258), .B2(n_261), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_439), .A2(n_264), .B1(n_251), .B2(n_225), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_423), .A2(n_264), .B1(n_251), .B2(n_225), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_394), .Y(n_468) );
AOI32xp33_ASAP7_75t_L g469 ( .A1(n_394), .A2(n_13), .A3(n_243), .B1(n_218), .B2(n_17), .Y(n_469) );
NAND2x1_ASAP7_75t_SL g470 ( .A(n_395), .B(n_15), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_395), .B(n_247), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_410), .Y(n_472) );
OAI322xp33_ASAP7_75t_L g473 ( .A1(n_434), .A2(n_159), .A3(n_247), .B1(n_225), .B2(n_223), .C1(n_23), .C2(n_24), .Y(n_473) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_412), .B(n_159), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_413), .B(n_16), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_399), .A2(n_243), .B(n_218), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_393), .B(n_19), .C(n_20), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_416), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_396), .Y(n_479) );
AOI211xp5_ASAP7_75t_L g480 ( .A1(n_402), .A2(n_159), .B(n_25), .C(n_36), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_417), .A2(n_159), .B1(n_142), .B2(n_40), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_417), .A2(n_142), .B1(n_38), .B2(n_42), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_424), .B(n_22), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_437), .B(n_177), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_398), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_392), .B(n_45), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_455), .A2(n_442), .B(n_400), .C(n_405), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_465), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_472), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_453), .B(n_429), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_479), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_485), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_450), .A2(n_419), .B(n_429), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_446), .B(n_440), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_467), .Y(n_496) );
AOI322xp5_ASAP7_75t_L g497 ( .A1(n_447), .A2(n_435), .A3(n_431), .B1(n_427), .B2(n_419), .C1(n_409), .C2(n_425), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_471), .B(n_408), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_464), .B(n_401), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_449), .B(n_432), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_468), .B(n_436), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_471), .B(n_432), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_445), .B(n_458), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_478), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_478), .B(n_425), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_454), .B(n_421), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_456), .A2(n_421), .B(n_418), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_443), .B(n_418), .Y(n_509) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_457), .A2(n_416), .B(n_50), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_448), .B(n_49), .Y(n_511) );
XNOR2x1_ASAP7_75t_L g512 ( .A(n_486), .B(n_52), .Y(n_512) );
XOR2xp5_ASAP7_75t_L g513 ( .A(n_460), .B(n_55), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_459), .B(n_177), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_498), .B(n_451), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_488), .Y(n_517) );
OAI211xp5_ASAP7_75t_SL g518 ( .A1(n_487), .A2(n_469), .B(n_481), .C(n_482), .Y(n_518) );
BUFx2_ASAP7_75t_SL g519 ( .A(n_512), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_515), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_497), .A2(n_470), .B(n_480), .C(n_477), .Y(n_521) );
XNOR2x1_ASAP7_75t_L g522 ( .A(n_513), .B(n_482), .Y(n_522) );
AOI211xp5_ASAP7_75t_L g523 ( .A1(n_491), .A2(n_463), .B(n_466), .C(n_475), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_498), .B(n_462), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_494), .A2(n_473), .B1(n_483), .B2(n_481), .C(n_476), .Y(n_525) );
O2A1O1Ixp5_ASAP7_75t_L g526 ( .A1(n_502), .A2(n_474), .B(n_484), .C(n_59), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_495), .Y(n_527) );
AOI21x1_ASAP7_75t_L g528 ( .A1(n_514), .A2(n_56), .B(n_57), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_499), .A2(n_61), .B1(n_62), .B2(n_63), .C(n_64), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g530 ( .A(n_500), .B(n_65), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_497), .B(n_508), .C(n_496), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_503), .B(n_183), .Y(n_532) );
AOI211xp5_ASAP7_75t_SL g533 ( .A1(n_518), .A2(n_511), .B(n_505), .C(n_503), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_531), .B(n_490), .C(n_492), .D(n_493), .Y(n_534) );
AOI21xp33_ASAP7_75t_SL g535 ( .A1(n_522), .A2(n_510), .B(n_489), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g536 ( .A1(n_516), .A2(n_507), .B1(n_501), .B2(n_509), .C1(n_504), .C2(n_506), .Y(n_536) );
AOI211xp5_ASAP7_75t_L g537 ( .A1(n_521), .A2(n_510), .B(n_69), .C(n_72), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_519), .A2(n_142), .B1(n_73), .B2(n_75), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g539 ( .A1(n_523), .A2(n_66), .B(n_77), .C(n_178), .Y(n_539) );
NOR4xp25_ASAP7_75t_L g540 ( .A(n_520), .B(n_527), .C(n_517), .D(n_525), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_524), .A2(n_525), .B1(n_526), .B2(n_529), .C(n_530), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_540), .B(n_532), .Y(n_542) );
NOR2xp67_ASAP7_75t_L g543 ( .A(n_535), .B(n_528), .Y(n_543) );
AOI21x1_ASAP7_75t_L g544 ( .A1(n_539), .A2(n_529), .B(n_533), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_538), .B(n_536), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_546), .B(n_534), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_542), .B(n_537), .C(n_545), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_545), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_549), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_547), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_550), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_550), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_552), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_554), .Y(n_555) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_553), .B(n_551), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_556), .A2(n_548), .B1(n_543), .B2(n_544), .Y(n_557) );
endmodule