module real_aes_8244_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_85), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g455 ( .A(n_0), .Y(n_455) );
INVx1_ASAP7_75t_L g505 ( .A(n_1), .Y(n_505) );
INVx1_ASAP7_75t_L g201 ( .A(n_2), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_3), .A2(n_77), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_3), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_4), .A2(n_38), .B1(n_157), .B2(n_521), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g181 ( .A1(n_5), .A2(n_138), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_6), .B(n_131), .Y(n_496) );
AND2x6_ASAP7_75t_L g143 ( .A(n_7), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_8), .A2(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_9), .B(n_39), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_10), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g188 ( .A(n_11), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_12), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g500 ( .A(n_13), .Y(n_500) );
INVx1_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
INVx1_ASAP7_75t_L g246 ( .A(n_15), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_16), .B(n_169), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_17), .B(n_132), .Y(n_477) );
AO32x2_ASAP7_75t_L g529 ( .A1(n_18), .A2(n_131), .A3(n_166), .B1(n_483), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_19), .B(n_157), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_20), .B(n_152), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_21), .B(n_132), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_22), .A2(n_50), .B1(n_157), .B2(n_521), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_23), .B(n_138), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_24), .A2(n_74), .B1(n_157), .B2(n_169), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_25), .B(n_157), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_26), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_27), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_29), .B(n_190), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_30), .B(n_186), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_31), .A2(n_42), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_31), .Y(n_748) );
INVx1_ASAP7_75t_L g175 ( .A(n_32), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_33), .B(n_190), .Y(n_544) );
INVx2_ASAP7_75t_L g141 ( .A(n_34), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_35), .B(n_157), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_36), .B(n_190), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_37), .A2(n_143), .B(n_147), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g173 ( .A(n_40), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_41), .B(n_186), .Y(n_256) );
CKINVDCx14_ASAP7_75t_R g749 ( .A(n_42), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_43), .B(n_157), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_44), .A2(n_86), .B1(n_219), .B2(n_521), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_45), .B(n_157), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_46), .B(n_157), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_47), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_48), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_49), .B(n_138), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_51), .A2(n_60), .B1(n_157), .B2(n_169), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_52), .A2(n_147), .B1(n_169), .B2(n_171), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_53), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_54), .B(n_157), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_55), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_56), .B(n_157), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_57), .A2(n_156), .B(n_185), .C(n_187), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_58), .Y(n_260) );
INVx1_ASAP7_75t_L g183 ( .A(n_59), .Y(n_183) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_62), .B(n_157), .Y(n_506) );
INVx1_ASAP7_75t_L g135 ( .A(n_63), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
AO32x2_ASAP7_75t_L g524 ( .A1(n_65), .A2(n_131), .A3(n_226), .B1(n_483), .B2(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g563 ( .A(n_66), .Y(n_563) );
INVx1_ASAP7_75t_L g539 ( .A(n_67), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_SL g151 ( .A1(n_68), .A2(n_152), .B(n_153), .C(n_156), .Y(n_151) );
INVxp67_ASAP7_75t_L g154 ( .A(n_69), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_70), .B(n_169), .Y(n_540) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_72), .Y(n_179) );
INVx1_ASAP7_75t_L g253 ( .A(n_73), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_75), .A2(n_143), .B(n_147), .C(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_76), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_77), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_78), .B(n_169), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_79), .B(n_202), .Y(n_215) );
INVx2_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_81), .B(n_152), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_82), .A2(n_102), .B1(n_111), .B2(n_758), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_83), .B(n_169), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_84), .A2(n_143), .B(n_147), .C(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g452 ( .A(n_85), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g464 ( .A(n_85), .B(n_454), .Y(n_464) );
INVx2_ASAP7_75t_L g468 ( .A(n_85), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_87), .A2(n_100), .B1(n_169), .B2(n_170), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_88), .A2(n_461), .B1(n_747), .B2(n_750), .C1(n_752), .C2(n_753), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_89), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_90), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_91), .A2(n_143), .B(n_147), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_92), .Y(n_236) );
INVx1_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_94), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_95), .B(n_202), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_96), .B(n_169), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_97), .B(n_131), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_99), .A2(n_138), .B(n_145), .Y(n_137) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g760 ( .A(n_104), .Y(n_760) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g454 ( .A(n_105), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_459), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g757 ( .A(n_115), .Y(n_757) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_449), .B(n_456), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B1(n_123), .B2(n_448), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g448 ( .A(n_123), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_123), .A2(n_462), .B1(n_465), .B2(n_469), .Y(n_461) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_385), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_315), .C(n_346), .D(n_365), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_273), .C(n_288), .D(n_306), .Y(n_125) );
AOI222xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_208), .B1(n_249), .B2(n_261), .C1(n_266), .C2(n_268), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_191), .Y(n_127) );
INVx1_ASAP7_75t_L g329 ( .A(n_128), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_162), .Y(n_128) );
AND2x2_ASAP7_75t_L g192 ( .A(n_129), .B(n_180), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_129), .B(n_195), .Y(n_358) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g265 ( .A(n_130), .B(n_164), .Y(n_265) );
AND2x2_ASAP7_75t_L g274 ( .A(n_130), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g300 ( .A(n_130), .Y(n_300) );
AND2x2_ASAP7_75t_L g321 ( .A(n_130), .B(n_164), .Y(n_321) );
BUFx2_ASAP7_75t_L g344 ( .A(n_130), .Y(n_344) );
AND2x2_ASAP7_75t_L g368 ( .A(n_130), .B(n_165), .Y(n_368) );
AND2x2_ASAP7_75t_L g432 ( .A(n_130), .B(n_180), .Y(n_432) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_137), .B(n_159), .Y(n_130) );
INVx4_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_131), .A2(n_488), .B(n_496), .Y(n_487) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_133), .B(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g240 ( .A(n_138), .Y(n_240) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_139), .B(n_143), .Y(n_177) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g495 ( .A(n_140), .Y(n_495) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
INVx1_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx1_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
INVx4_ASAP7_75t_SL g158 ( .A(n_143), .Y(n_158) );
BUFx3_ASAP7_75t_L g483 ( .A(n_143), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_143), .A2(n_489), .B(n_492), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_143), .A2(n_499), .B(n_503), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_143), .A2(n_514), .B(n_518), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_143), .A2(n_538), .B(n_541), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B(n_151), .C(n_158), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_146), .A2(n_158), .B(n_183), .C(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_146), .A2(n_158), .B(n_242), .C(n_243), .Y(n_241) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx3_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
INVx1_ASAP7_75t_L g521 ( .A(n_148), .Y(n_521) );
INVx1_ASAP7_75t_L g517 ( .A(n_152), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_155), .B(n_188), .Y(n_187) );
INVx5_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g525 ( .A1(n_155), .A2(n_186), .B1(n_526), .B2(n_527), .Y(n_525) );
O2A1O1Ixp5_ASAP7_75t_SL g538 ( .A1(n_156), .A2(n_202), .B(n_539), .C(n_540), .Y(n_538) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g167 ( .A1(n_158), .A2(n_168), .B1(n_176), .B2(n_177), .Y(n_167) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_160), .A2(n_181), .B(n_189), .Y(n_180) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g221 ( .A(n_161), .B(n_222), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_161), .B(n_479), .C(n_483), .Y(n_478) );
AO21x1_ASAP7_75t_L g571 ( .A1(n_161), .A2(n_479), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g333 ( .A(n_162), .B(n_264), .Y(n_333) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_163), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
OR2x2_ASAP7_75t_L g293 ( .A(n_164), .B(n_196), .Y(n_293) );
AND2x2_ASAP7_75t_L g305 ( .A(n_164), .B(n_264), .Y(n_305) );
BUFx2_ASAP7_75t_L g437 ( .A(n_164), .Y(n_437) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g194 ( .A(n_165), .B(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g287 ( .A(n_165), .B(n_196), .Y(n_287) );
AND2x2_ASAP7_75t_L g340 ( .A(n_165), .B(n_180), .Y(n_340) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_165), .Y(n_376) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_178), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_166), .B(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_166), .A2(n_197), .B(n_205), .Y(n_196) );
INVx2_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
INVx2_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g174 ( .A(n_172), .Y(n_174) );
INVx4_ASAP7_75t_L g244 ( .A(n_172), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_177), .A2(n_198), .B(n_199), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_177), .A2(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g263 ( .A(n_180), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g275 ( .A(n_180), .Y(n_275) );
INVx2_ASAP7_75t_L g286 ( .A(n_180), .Y(n_286) );
BUFx2_ASAP7_75t_L g310 ( .A(n_180), .Y(n_310) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_180), .B(n_368), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_185), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_L g562 ( .A1(n_185), .A2(n_504), .B(n_563), .C(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx4_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_186), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_186), .A2(n_481), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g207 ( .A(n_190), .Y(n_207) );
INVx2_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_190), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_190), .A2(n_513), .B(n_522), .Y(n_512) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_190), .A2(n_537), .B(n_544), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
AOI332xp33_ASAP7_75t_L g288 ( .A1(n_192), .A2(n_289), .A3(n_293), .B1(n_294), .B2(n_298), .B3(n_301), .C1(n_302), .C2(n_304), .Y(n_288) );
NAND2x1_ASAP7_75t_L g373 ( .A(n_192), .B(n_264), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_192), .B(n_278), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_SL g306 ( .A1(n_193), .A2(n_307), .B(n_310), .C(n_311), .Y(n_306) );
AND2x2_ASAP7_75t_L g445 ( .A(n_193), .B(n_286), .Y(n_445) );
INVx3_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g342 ( .A(n_194), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g347 ( .A(n_194), .B(n_344), .Y(n_347) );
INVx1_ASAP7_75t_L g278 ( .A(n_195), .Y(n_278) );
AND2x2_ASAP7_75t_L g381 ( .A(n_195), .B(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_195), .B(n_321), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_195), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_195), .B(n_299), .Y(n_407) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g264 ( .A(n_196), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_204), .Y(n_200) );
INVx2_ASAP7_75t_L g481 ( .A(n_202), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_202), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_202), .A2(n_560), .B(n_561), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_204), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_207), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_207), .B(n_260), .Y(n_259) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_208), .A2(n_367), .A3(n_374), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_223), .Y(n_208) );
AND2x2_ASAP7_75t_L g249 ( .A(n_209), .B(n_250), .Y(n_249) );
NAND2x1_ASAP7_75t_SL g269 ( .A(n_209), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_209), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_209), .B(n_272), .Y(n_361) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_210), .A2(n_274), .B(n_276), .C(n_279), .Y(n_273) );
OR2x2_ASAP7_75t_L g290 ( .A(n_210), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g303 ( .A(n_210), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_210), .B(n_251), .Y(n_309) );
INVx2_ASAP7_75t_L g327 ( .A(n_210), .Y(n_327) );
AND2x2_ASAP7_75t_L g338 ( .A(n_210), .B(n_292), .Y(n_338) );
AND2x2_ASAP7_75t_L g370 ( .A(n_210), .B(n_328), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_210), .B(n_297), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_210), .B(n_223), .Y(n_379) );
AND2x2_ASAP7_75t_L g413 ( .A(n_210), .B(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_210), .B(n_316), .Y(n_447) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g211 ( .A1(n_212), .A2(n_213), .B(n_220), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_217), .A2(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
INVx1_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_220), .A2(n_498), .B(n_507), .Y(n_497) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_220), .A2(n_558), .B(n_565), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_223), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g355 ( .A(n_223), .Y(n_355) );
AND2x2_ASAP7_75t_L g417 ( .A(n_223), .B(n_338), .Y(n_417) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
OR2x2_ASAP7_75t_L g271 ( .A(n_224), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g281 ( .A(n_224), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_224), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g389 ( .A(n_224), .Y(n_389) );
AND2x2_ASAP7_75t_L g406 ( .A(n_224), .B(n_251), .Y(n_406) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g297 ( .A(n_225), .B(n_237), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_225), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g337 ( .A(n_225), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_225), .B(n_292), .Y(n_428) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g250 ( .A(n_238), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g272 ( .A(n_238), .Y(n_272) );
AND2x2_ASAP7_75t_L g328 ( .A(n_238), .B(n_292), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g502 ( .A(n_244), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_244), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g430 ( .A(n_249), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_250), .Y(n_434) );
INVx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_258), .B(n_259), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_263), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_263), .B(n_368), .Y(n_426) );
OR2x2_ASAP7_75t_L g267 ( .A(n_264), .B(n_265), .Y(n_267) );
INVx1_ASAP7_75t_SL g319 ( .A(n_264), .Y(n_319) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_270), .A2(n_323), .B1(n_325), .B2(n_329), .C(n_330), .Y(n_322) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g350 ( .A(n_271), .B(n_314), .Y(n_350) );
INVx2_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_272), .B(n_292), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_272), .B(n_295), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_272), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_274), .B(n_278), .Y(n_324) );
AND2x4_ASAP7_75t_L g299 ( .A(n_275), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g412 ( .A(n_278), .B(n_368), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_281), .B(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g420 ( .A(n_282), .Y(n_420) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g320 ( .A(n_286), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g392 ( .A(n_286), .B(n_368), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_286), .B(n_305), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g352 ( .A1(n_287), .A2(n_321), .A3(n_328), .B1(n_353), .B2(n_356), .C1(n_357), .C2(n_359), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_287), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
INVx2_ASAP7_75t_L g295 ( .A(n_292), .Y(n_295) );
INVx1_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_293), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g390 ( .A(n_295), .B(n_303), .Y(n_390) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g302 ( .A(n_297), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g345 ( .A(n_297), .B(n_338), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_297), .B(n_309), .Y(n_349) );
OAI21xp33_ASAP7_75t_SL g359 ( .A1(n_298), .A2(n_360), .B(n_362), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_298), .A2(n_430), .B1(n_431), .B2(n_433), .Y(n_429) );
INVx3_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_299), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_299), .B(n_319), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_301), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g441 ( .A(n_308), .Y(n_441) );
INVx4_ASAP7_75t_L g314 ( .A(n_309), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_309), .B(n_336), .Y(n_384) );
INVx1_ASAP7_75t_SL g396 ( .A(n_310), .Y(n_396) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_314), .B(n_410), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B(n_322), .C(n_339), .Y(n_315) );
OAI221xp5_ASAP7_75t_SL g435 ( .A1(n_317), .A2(n_355), .B1(n_434), .B2(n_436), .C(n_438), .Y(n_435) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_319), .B(n_432), .Y(n_431) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_320), .A2(n_397), .A3(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g401 ( .A(n_326), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_328), .B(n_337), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_338), .B(n_441), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_348), .B1(n_350), .B2(n_351), .C(n_352), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_347), .A2(n_416), .B(n_418), .C(n_421), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_350), .B(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_361), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g405 ( .A(n_361), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B(n_371), .C(n_380), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_369), .A2(n_379), .B1(n_443), .B2(n_444), .C(n_446), .Y(n_442) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_375), .B2(n_378), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_382), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_SL g443 ( .A(n_382), .Y(n_443) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_415), .C(n_435), .D(n_442), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_391), .B(n_393), .C(n_411), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_399), .C(n_403), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g422 ( .A(n_400), .Y(n_422) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g433 ( .A(n_401), .B(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_427), .C(n_429), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_432), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22x1_ASAP7_75t_SL g750 ( .A1(n_448), .A2(n_467), .B1(n_470), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_452), .Y(n_458) );
NOR2x2_ASAP7_75t_L g755 ( .A(n_453), .B(n_468), .Y(n_755) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g467 ( .A(n_454), .B(n_468), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_456), .B(n_460), .C(n_756), .Y(n_459) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g751 ( .A(n_463), .Y(n_751) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_472), .B(n_681), .Y(n_471) );
NOR5xp2_ASAP7_75t_L g472 ( .A(n_473), .B(n_594), .C(n_640), .D(n_653), .E(n_665), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_508), .B(n_548), .C(n_575), .Y(n_473) );
INVx1_ASAP7_75t_SL g676 ( .A(n_474), .Y(n_676) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
AND2x2_ASAP7_75t_L g600 ( .A(n_475), .B(n_485), .Y(n_600) );
AND2x2_ASAP7_75t_L g628 ( .A(n_475), .B(n_574), .Y(n_628) );
AND2x2_ASAP7_75t_L g636 ( .A(n_475), .B(n_579), .Y(n_636) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g566 ( .A(n_476), .B(n_486), .Y(n_566) );
INVx2_ASAP7_75t_L g578 ( .A(n_476), .Y(n_578) );
AND2x2_ASAP7_75t_L g703 ( .A(n_476), .B(n_645), .Y(n_703) );
OR2x2_ASAP7_75t_L g705 ( .A(n_476), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g572 ( .A(n_477), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_481), .A2(n_493), .B(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_481), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_483), .A2(n_559), .B(n_562), .Y(n_558) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_588), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_485), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g730 ( .A(n_485), .B(n_570), .Y(n_730) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
AND2x2_ASAP7_75t_L g573 ( .A(n_486), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g620 ( .A(n_486), .Y(n_620) );
AND2x2_ASAP7_75t_L g645 ( .A(n_486), .B(n_557), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_486), .B(n_678), .Y(n_715) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g579 ( .A(n_487), .B(n_557), .Y(n_579) );
AND2x2_ASAP7_75t_L g593 ( .A(n_487), .B(n_556), .Y(n_593) );
AND2x2_ASAP7_75t_L g610 ( .A(n_487), .B(n_497), .Y(n_610) );
AND2x2_ASAP7_75t_L g667 ( .A(n_487), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_487), .B(n_574), .Y(n_680) );
AND2x2_ASAP7_75t_L g732 ( .A(n_487), .B(n_657), .Y(n_732) );
INVx2_ASAP7_75t_L g504 ( .A(n_495), .Y(n_504) );
AND2x2_ASAP7_75t_L g555 ( .A(n_497), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g574 ( .A(n_497), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_497), .B(n_557), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_533), .B(n_545), .Y(n_508) );
INVx1_ASAP7_75t_SL g664 ( .A(n_509), .Y(n_664) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_523), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_511), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g547 ( .A(n_512), .Y(n_547) );
INVx1_ASAP7_75t_L g584 ( .A(n_512), .Y(n_584) );
AND2x2_ASAP7_75t_L g605 ( .A(n_512), .B(n_528), .Y(n_605) );
AND2x2_ASAP7_75t_L g639 ( .A(n_512), .B(n_529), .Y(n_639) );
OR2x2_ASAP7_75t_L g658 ( .A(n_512), .B(n_535), .Y(n_658) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_512), .Y(n_672) );
AND2x2_ASAP7_75t_L g685 ( .A(n_512), .B(n_686), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_523), .A2(n_607), .B1(n_608), .B2(n_617), .Y(n_606) );
AND2x2_ASAP7_75t_L g690 ( .A(n_523), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
INVx1_ASAP7_75t_L g551 ( .A(n_524), .Y(n_551) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_524), .Y(n_588) );
INVx1_ASAP7_75t_L g599 ( .A(n_524), .Y(n_599) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_529), .Y(n_614) );
OR2x2_ASAP7_75t_L g568 ( .A(n_528), .B(n_553), .Y(n_568) );
AND2x2_ASAP7_75t_L g598 ( .A(n_528), .B(n_599), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_528), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g546 ( .A(n_529), .B(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g655 ( .A(n_529), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_533), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g633 ( .A(n_534), .B(n_599), .Y(n_633) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g545 ( .A(n_535), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g604 ( .A(n_535), .Y(n_604) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g553 ( .A(n_536), .Y(n_553) );
OR2x2_ASAP7_75t_L g583 ( .A(n_536), .B(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_536), .Y(n_638) );
AOI32xp33_ASAP7_75t_L g675 ( .A1(n_545), .A2(n_605), .A3(n_676), .B1(n_677), .B2(n_679), .Y(n_675) );
AND2x2_ASAP7_75t_L g601 ( .A(n_546), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_546), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_546), .B(n_633), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_546), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_554), .B1(n_567), .B2(n_569), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g654 ( .A(n_550), .B(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_551), .B(n_553), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_552), .A2(n_576), .B1(n_580), .B2(n_590), .Y(n_575) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_598), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_552), .A2(n_566), .B(n_614), .C(n_649), .Y(n_648) );
OAI332xp33_ASAP7_75t_L g653 ( .A1(n_552), .A2(n_654), .A3(n_656), .B1(n_658), .B2(n_659), .B3(n_661), .C1(n_662), .C2(n_664), .Y(n_653) );
INVx2_ASAP7_75t_L g694 ( .A(n_552), .Y(n_694) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
INVx1_ASAP7_75t_L g687 ( .A(n_553), .Y(n_687) );
AND2x2_ASAP7_75t_L g741 ( .A(n_553), .B(n_605), .Y(n_741) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_566), .Y(n_554) );
AND2x2_ASAP7_75t_L g621 ( .A(n_556), .B(n_571), .Y(n_621) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g570 ( .A(n_557), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g669 ( .A(n_557), .B(n_571), .Y(n_669) );
INVx1_ASAP7_75t_L g678 ( .A(n_557), .Y(n_678) );
INVx1_ASAP7_75t_L g652 ( .A(n_566), .Y(n_652) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g736 ( .A(n_568), .B(n_588), .Y(n_736) );
INVx1_ASAP7_75t_SL g647 ( .A(n_569), .Y(n_647) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
AND2x2_ASAP7_75t_L g674 ( .A(n_570), .B(n_632), .Y(n_674) );
INVx1_ASAP7_75t_L g693 ( .A(n_570), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_570), .B(n_660), .Y(n_695) );
INVx1_ASAP7_75t_L g592 ( .A(n_571), .Y(n_592) );
AND2x2_ASAP7_75t_L g596 ( .A(n_573), .B(n_577), .Y(n_596) );
AND2x2_ASAP7_75t_L g663 ( .A(n_573), .B(n_621), .Y(n_663) );
INVx2_ASAP7_75t_L g706 ( .A(n_573), .Y(n_706) );
INVx2_ASAP7_75t_L g589 ( .A(n_574), .Y(n_589) );
AND2x2_ASAP7_75t_L g591 ( .A(n_574), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g607 ( .A(n_577), .Y(n_607) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_578), .B(n_651), .Y(n_657) );
OR2x2_ASAP7_75t_L g721 ( .A(n_578), .B(n_680), .Y(n_721) );
INVx1_ASAP7_75t_L g745 ( .A(n_578), .Y(n_745) );
INVx1_ASAP7_75t_L g701 ( .A(n_579), .Y(n_701) );
AND2x2_ASAP7_75t_L g746 ( .A(n_579), .B(n_589), .Y(n_746) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_583), .A2(n_609), .B1(n_611), .B2(n_615), .Y(n_608) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI322xp33_ASAP7_75t_SL g692 ( .A1(n_586), .A2(n_693), .A3(n_694), .B1(n_695), .B2(n_696), .C1(n_699), .C2(n_701), .Y(n_692) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_L g689 ( .A(n_587), .B(n_605), .Y(n_689) );
OR2x2_ASAP7_75t_L g723 ( .A(n_587), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g726 ( .A(n_587), .B(n_658), .Y(n_726) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g671 ( .A(n_588), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g727 ( .A(n_588), .B(n_658), .Y(n_727) );
INVx3_ASAP7_75t_L g660 ( .A(n_589), .Y(n_660) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g716 ( .A(n_591), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_593), .A2(n_596), .B1(n_597), .B2(n_600), .C1(n_601), .C2(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
NAND3xp33_ASAP7_75t_SL g594 ( .A(n_595), .B(n_606), .C(n_623), .Y(n_594) );
AND2x2_ASAP7_75t_L g711 ( .A(n_598), .B(n_612), .Y(n_711) );
BUFx2_ASAP7_75t_L g602 ( .A(n_599), .Y(n_602) );
INVx1_ASAP7_75t_L g643 ( .A(n_599), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_600), .A2(n_636), .B1(n_689), .B2(n_690), .C(n_692), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_602), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_605), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_605), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_610), .B(n_621), .Y(n_622) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_612), .A2(n_618), .B(n_622), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_612), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g709 ( .A(n_614), .B(n_691), .Y(n_709) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g632 ( .A(n_620), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_621), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g738 ( .A(n_621), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_629), .B1(n_630), .B2(n_633), .C(n_634), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_625), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g734 ( .A(n_633), .B(n_639), .Y(n_734) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OAI31xp33_ASAP7_75t_SL g702 ( .A1(n_637), .A2(n_676), .A3(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g691 ( .A(n_638), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_639), .B(n_643), .Y(n_742) );
OAI221xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_644), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_640) );
INVx1_ASAP7_75t_L g646 ( .A(n_642), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_645), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g661 ( .A(n_654), .Y(n_661) );
INVx2_ASAP7_75t_L g697 ( .A(n_655), .Y(n_697) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g683 ( .A(n_660), .B(n_669), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g733 ( .A1(n_660), .A2(n_677), .B(n_734), .C(n_735), .Y(n_733) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_661), .A2(n_666), .B1(n_670), .B2(n_673), .C(n_675), .Y(n_665) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_664), .A2(n_729), .B(n_731), .C(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_667), .A2(n_718), .B1(n_720), .B2(n_722), .C(n_725), .Y(n_717) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NOR4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_707), .C(n_728), .D(n_739), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B(n_688), .C(n_702), .Y(n_682) );
INVx1_ASAP7_75t_SL g737 ( .A(n_689), .Y(n_737) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_SL g700 ( .A(n_698), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_705), .A2(n_714), .B1(n_726), .B2(n_727), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_712), .C(n_717), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI31xp33_ASAP7_75t_L g739 ( .A1(n_710), .A2(n_740), .A3(n_742), .B(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g752 ( .A(n_747), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule