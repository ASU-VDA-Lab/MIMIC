module fake_ibex_961_n_1393 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1393);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1393;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1115;
wire n_998;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g263 ( 
.A(n_119),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_95),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_78),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_82),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_85),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_64),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_162),
.B(n_215),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_122),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_153),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_161),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_242),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_14),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_205),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_125),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_132),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_118),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_29),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_33),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_31),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_156),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_142),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_240),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_157),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_31),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_52),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_103),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_207),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_10),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_124),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_151),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_86),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_137),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_203),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_143),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_110),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_252),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_88),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_166),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_104),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_147),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_174),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_185),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_55),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_24),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_97),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_149),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_182),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_152),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_68),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_71),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_211),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_128),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_84),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_169),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_229),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_232),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_208),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_217),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_6),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_214),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_67),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_131),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_65),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_244),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_114),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_123),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_254),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_101),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_231),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_98),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_243),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_18),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_224),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_148),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_12),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_68),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_102),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_17),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_126),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_112),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_92),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_219),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_49),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_29),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_188),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_25),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_184),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_51),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_241),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_167),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_36),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_176),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_255),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_30),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_170),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_258),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_33),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_164),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_163),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_212),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_93),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_0),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_23),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_223),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_155),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_13),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_178),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_94),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_9),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_175),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_225),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_139),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_187),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_79),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_70),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_9),
.B(n_165),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_19),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_30),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_8),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_228),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_67),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_186),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_199),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_234),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_189),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_28),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_50),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_80),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_168),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_194),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_190),
.B(n_108),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_11),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_42),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_89),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_70),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_81),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_76),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_115),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_140),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_50),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_12),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_47),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_210),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_35),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_260),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_121),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_69),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_179),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_5),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_48),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_26),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_117),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_318),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_361),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_284),
.A2(n_87),
.B(n_83),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_0),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_281),
.Y(n_449)
);

OAI22x1_ASAP7_75t_SL g450 ( 
.A1(n_314),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_284),
.A2(n_91),
.B(n_90),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_291),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_275),
.B(n_96),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_274),
.B(n_1),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_289),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_318),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_291),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_318),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_307),
.B(n_327),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_344),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_289),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_355),
.B(n_8),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_286),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_345),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_275),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_314),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_323),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_286),
.B(n_15),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_15),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_352),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_347),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_352),
.B(n_16),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_345),
.A2(n_383),
.B(n_356),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_347),
.B(n_19),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_375),
.B(n_20),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_278),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_270),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_356),
.A2(n_120),
.B(n_262),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_441),
.B(n_20),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_399),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_405),
.B(n_99),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g492 ( 
.A(n_405),
.B(n_100),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_21),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_278),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_363),
.B(n_24),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

OAI22x1_ASAP7_75t_SL g498 ( 
.A1(n_331),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_287),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_288),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_298),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_303),
.B(n_27),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_441),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_305),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_331),
.A2(n_372),
.B1(n_387),
.B2(n_336),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_404),
.B(n_32),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_337),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_412),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_336),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_278),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_373),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_407),
.B(n_32),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_363),
.B(n_398),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_407),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_398),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_420),
.A2(n_134),
.B(n_259),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_434),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_378),
.B(n_34),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_372),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_263),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_393),
.B(n_37),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_396),
.B(n_38),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_441),
.B(n_39),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_319),
.B(n_40),
.Y(n_531)
);

CKINVDCx11_ASAP7_75t_R g532 ( 
.A(n_387),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_264),
.Y(n_533)
);

CKINVDCx11_ASAP7_75t_R g534 ( 
.A(n_428),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_409),
.B(n_40),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_319),
.B(n_334),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_265),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_41),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_433),
.B(n_41),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_319),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_496),
.B(n_266),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_268),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_472),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_496),
.B(n_267),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_496),
.B(n_271),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_536),
.B(n_408),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_475),
.A2(n_417),
.B1(n_418),
.B2(n_408),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_478),
.Y(n_553)
);

NOR2x1p5_ASAP7_75t_L g554 ( 
.A(n_494),
.B(n_417),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_531),
.B(n_304),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_499),
.B(n_423),
.C(n_418),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_483),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_480),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_524),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_516),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_483),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_334),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_505),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_481),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_516),
.B(n_343),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_540),
.B(n_273),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_493),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_483),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_334),
.Y(n_573)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_461),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_524),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_540),
.B(n_277),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_483),
.B(n_279),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_471),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_540),
.B(n_282),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_499),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_540),
.B(n_283),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

AND3x2_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_465),
.C(n_531),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_521),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_542),
.B(n_304),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_528),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_528),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_529),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_532),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_540),
.B(n_293),
.Y(n_594)
);

BUFx6f_ASAP7_75t_SL g595 ( 
.A(n_529),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_521),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_521),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_499),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_519),
.Y(n_600)
);

INVxp33_ASAP7_75t_SL g601 ( 
.A(n_484),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_428),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_446),
.A2(n_317),
.B1(n_333),
.B2(n_315),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_535),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_527),
.B(n_533),
.Y(n_606)
);

AND3x2_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_349),
.C(n_440),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_535),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_527),
.B(n_294),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_445),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_445),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_519),
.B(n_279),
.Y(n_612)
);

BUFx6f_ASAP7_75t_SL g613 ( 
.A(n_535),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_453),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_458),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_494),
.B(n_295),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_539),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_448),
.A2(n_317),
.B1(n_333),
.B2(n_315),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

AND3x1_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_310),
.C(n_300),
.Y(n_622)
);

AND3x2_ASAP7_75t_L g623 ( 
.A(n_489),
.B(n_313),
.C(n_311),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_484),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_449),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_449),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_458),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_519),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_527),
.B(n_322),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_527),
.B(n_325),
.Y(n_631)
);

AO22x2_ASAP7_75t_L g632 ( 
.A1(n_455),
.A2(n_280),
.B1(n_350),
.B2(n_332),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_541),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_537),
.B(n_285),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_458),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_466),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_530),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_533),
.B(n_326),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_453),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_448),
.A2(n_370),
.B1(n_368),
.B2(n_414),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_453),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_453),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_530),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_532),
.Y(n_644)
);

INVxp67_ASAP7_75t_R g645 ( 
.A(n_450),
.Y(n_645)
);

INVx6_ASAP7_75t_L g646 ( 
.A(n_469),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_449),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_520),
.A2(n_419),
.B1(n_370),
.B2(n_368),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_534),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_477),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_500),
.B(n_340),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_474),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_534),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_491),
.B(n_285),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_456),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_474),
.B(n_342),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_501),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_452),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_518),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_492),
.B(n_346),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_457),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_456),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_454),
.B(n_296),
.C(n_292),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_503),
.B(n_290),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_504),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_456),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_457),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_459),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_459),
.B(n_348),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_507),
.B(n_354),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_456),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_462),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_504),
.A2(n_419),
.B1(n_414),
.B2(n_367),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_512),
.B(n_290),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_447),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_462),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_525),
.A2(n_297),
.B1(n_306),
.B2(n_376),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_517),
.B(n_338),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_538),
.B(n_338),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_508),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_468),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_468),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_460),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_460),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_482),
.B(n_357),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_486),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_467),
.B(n_351),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_464),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_486),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_464),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_487),
.B(n_351),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_464),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_487),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_464),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_488),
.B(n_358),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_488),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_497),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_497),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_447),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_506),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_506),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_511),
.B(n_360),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_525),
.B(n_401),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_704),
.A2(n_473),
.B1(n_470),
.B2(n_509),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_600),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_637),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_309),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_547),
.A2(n_511),
.B1(n_523),
.B2(n_515),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_600),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_704),
.A2(n_509),
.B1(n_432),
.B2(n_364),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_658),
.B(n_401),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_602),
.B(n_330),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_602),
.B(n_381),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_628),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_560),
.B(n_495),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_604),
.A2(n_463),
.B1(n_498),
.B2(n_526),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_643),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_675),
.B(n_403),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_588),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_554),
.B(n_476),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_547),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_547),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_563),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_634),
.B(n_410),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_642),
.A2(n_485),
.B(n_451),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_612),
.B(n_413),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_563),
.A2(n_515),
.B1(n_513),
.B2(n_523),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_563),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_553),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_574),
.A2(n_424),
.B1(n_384),
.B2(n_426),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_603),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_476),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_651),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_545),
.B(n_476),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_643),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_545),
.B(n_413),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_568),
.B(n_416),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_568),
.B(n_421),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_679),
.B(n_421),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_680),
.B(n_269),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_570),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_643),
.A2(n_406),
.B1(n_402),
.B2(n_437),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_573),
.A2(n_379),
.B1(n_386),
.B2(n_388),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_543),
.B(n_272),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_665),
.B(n_678),
.C(n_692),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_676),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_664),
.B(n_421),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_674),
.B(n_648),
.C(n_555),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_550),
.B(n_688),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_625),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_665),
.A2(n_389),
.B1(n_390),
.B2(n_415),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_653),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_646),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_555),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_546),
.A2(n_451),
.B1(n_485),
.B2(n_522),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_589),
.B(n_299),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_590),
.B(n_301),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_591),
.A2(n_425),
.B1(n_427),
.B2(n_429),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_552),
.A2(n_522),
.B1(n_451),
.B2(n_485),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_644),
.B(n_42),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_626),
.B(n_522),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_595),
.B(n_436),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_592),
.B(n_302),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_646),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_643),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_596),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_641),
.B(n_276),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_646),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_605),
.B(n_308),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_639),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_647),
.B(n_43),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_676),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_596),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_676),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_608),
.B(n_312),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_595),
.B(n_369),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_623),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_614),
.B(n_316),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_615),
.B(n_320),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_613),
.B(n_382),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_660),
.B(n_397),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_619),
.B(n_321),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_621),
.B(n_629),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_613),
.B(n_324),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_620),
.B(n_328),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_633),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_558),
.A2(n_510),
.B1(n_479),
.B2(n_443),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_682),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_618),
.B(n_329),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_561),
.A2(n_567),
.B1(n_571),
.B2(n_565),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_581),
.A2(n_510),
.B1(n_479),
.B2(n_439),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_618),
.B(n_335),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_583),
.B(n_339),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_682),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_639),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_599),
.B(n_341),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_607),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_636),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_640),
.B(n_353),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_622),
.A2(n_377),
.B1(n_359),
.B2(n_430),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_659),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_586),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_577),
.B(n_544),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_616),
.B(n_362),
.Y(n_807)
);

AND2x6_ASAP7_75t_SL g808 ( 
.A(n_645),
.B(n_422),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_624),
.B(n_366),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_578),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_548),
.B(n_371),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_579),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_579),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_580),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_548),
.B(n_374),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_549),
.B(n_380),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_662),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_549),
.B(n_692),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_657),
.A2(n_395),
.B(n_391),
.C(n_385),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_652),
.A2(n_510),
.B(n_479),
.C(n_45),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_652),
.B(n_43),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_616),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_690),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_671),
.B(n_44),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_557),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_593),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_556),
.B(n_694),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_700),
.B(n_105),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_671),
.B(n_45),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_551),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_668),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_698),
.B(n_46),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_655),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_673),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_562),
.B(n_53),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_572),
.B(n_107),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_655),
.B(n_54),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_657),
.B(n_56),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_661),
.B(n_109),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_677),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_580),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_686),
.B(n_56),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_661),
.B(n_111),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_654),
.B(n_57),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_683),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_686),
.B(n_58),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_638),
.B(n_58),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_638),
.B(n_113),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_687),
.B(n_59),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_697),
.B(n_116),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_632),
.B(n_59),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_699),
.B(n_701),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_670),
.B(n_127),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_587),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_670),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_702),
.B(n_129),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_696),
.B(n_130),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_649),
.B(n_60),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_703),
.B(n_60),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_61),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_601),
.B(n_61),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_735),
.B(n_632),
.Y(n_863)
);

AOI21xp33_ASAP7_75t_L g864 ( 
.A1(n_791),
.A2(n_601),
.B(n_632),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_792),
.A2(n_747),
.B1(n_788),
.B2(n_718),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_726),
.A2(n_584),
.B(n_569),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_708),
.B(n_609),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_707),
.B(n_681),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_750),
.A2(n_631),
.B(n_609),
.C(n_630),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_751),
.B(n_630),
.Y(n_870)
);

AO22x1_ASAP7_75t_L g871 ( 
.A1(n_826),
.A2(n_650),
.B1(n_63),
.B2(n_65),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_792),
.A2(n_767),
.B1(n_737),
.B2(n_756),
.Y(n_872)
);

OAI321xp33_ASAP7_75t_L g873 ( 
.A1(n_744),
.A2(n_606),
.A3(n_631),
.B1(n_582),
.B2(n_584),
.C(n_576),
.Y(n_873)
);

NOR2x1_ASAP7_75t_L g874 ( 
.A(n_752),
.B(n_576),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_763),
.B(n_656),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_713),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_762),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_728),
.A2(n_594),
.B(n_606),
.Y(n_878)
);

AO22x1_ASAP7_75t_L g879 ( 
.A1(n_720),
.A2(n_852),
.B1(n_733),
.B2(n_783),
.Y(n_879)
);

OR2x6_ASAP7_75t_SL g880 ( 
.A(n_845),
.B(n_62),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_716),
.B(n_663),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_728),
.A2(n_667),
.B(n_672),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_731),
.A2(n_667),
.B(n_672),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_757),
.A2(n_559),
.B(n_575),
.Y(n_884)
);

INVx11_ASAP7_75t_L g885 ( 
.A(n_773),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_787),
.B(n_63),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_828),
.A2(n_597),
.B(n_598),
.Y(n_887)
);

OAI321xp33_ASAP7_75t_L g888 ( 
.A1(n_744),
.A2(n_835),
.A3(n_830),
.B1(n_833),
.B2(n_705),
.C(n_821),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_722),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_734),
.B(n_66),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_785),
.A2(n_695),
.B(n_693),
.C(n_691),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_772),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_714),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_825),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_748),
.A2(n_776),
.B(n_774),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_721),
.B(n_71),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_740),
.B(n_72),
.Y(n_897)
);

OAI22x1_ASAP7_75t_L g898 ( 
.A1(n_803),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_898)
);

BUFx12f_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_712),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_757),
.A2(n_611),
.B(n_617),
.Y(n_901)
);

CKINVDCx10_ASAP7_75t_R g902 ( 
.A(n_717),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_723),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_761),
.A2(n_610),
.B(n_627),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_825),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_724),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_797),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_801),
.B(n_741),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_721),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_736),
.A2(n_689),
.B(n_685),
.C(n_684),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_805),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_75),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_730),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

INVx4_ASAP7_75t_R g915 ( 
.A(n_779),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_755),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_709),
.A2(n_635),
.B(n_585),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_800),
.A2(n_585),
.B(n_76),
.C(n_77),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_806),
.A2(n_213),
.B(n_257),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_741),
.B(n_77),
.Y(n_920)
);

BUFx12f_ASAP7_75t_L g921 ( 
.A(n_808),
.Y(n_921)
);

AO21x1_ASAP7_75t_L g922 ( 
.A1(n_851),
.A2(n_857),
.B(n_837),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_818),
.A2(n_133),
.B(n_135),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_745),
.B(n_136),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_761),
.A2(n_141),
.B(n_146),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_769),
.A2(n_154),
.B(n_159),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_769),
.A2(n_160),
.B(n_172),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_732),
.B(n_173),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_775),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_794),
.B(n_738),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_725),
.A2(n_177),
.B(n_180),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_743),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_853),
.A2(n_181),
.B1(n_183),
.B2(n_191),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_829),
.A2(n_192),
.B1(n_197),
.B2(n_200),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_794),
.B(n_201),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_719),
.A2(n_216),
.B(n_218),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_717),
.B(n_220),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_739),
.B(n_221),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_727),
.A2(n_222),
.B(n_226),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_859),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_711),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_758),
.A2(n_235),
.B(n_236),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_759),
.A2(n_237),
.B(n_238),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_856),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_753),
.B(n_804),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_729),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_862),
.B(n_251),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_754),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_729),
.A2(n_253),
.B1(n_835),
.B2(n_834),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_824),
.A2(n_717),
.B1(n_843),
.B2(n_847),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_765),
.A2(n_781),
.B(n_771),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_817),
.B(n_831),
.Y(n_952)
);

CKINVDCx6p67_ASAP7_75t_R g953 ( 
.A(n_838),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_777),
.A2(n_780),
.B(n_784),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_749),
.B(n_764),
.C(n_782),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_L g956 ( 
.A(n_742),
.B(n_749),
.C(n_798),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_816),
.B(n_807),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_820),
.B(n_789),
.C(n_793),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_841),
.A2(n_846),
.B(n_849),
.C(n_854),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_809),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_815),
.B(n_715),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_766),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_746),
.A2(n_815),
.B(n_795),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_760),
.A2(n_820),
.B(n_848),
.C(n_839),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_706),
.A2(n_710),
.B1(n_764),
.B2(n_861),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_819),
.A2(n_827),
.B(n_858),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_778),
.B(n_782),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_832),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_840),
.B(n_844),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_797),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_854),
.A2(n_858),
.B(n_849),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_850),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_860),
.A2(n_836),
.B1(n_790),
.B2(n_802),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_796),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_778),
.B(n_786),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_770),
.B(n_822),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_789),
.B(n_793),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_855),
.B(n_842),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_810),
.B(n_842),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_812),
.A2(n_813),
.B(n_814),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_708),
.B(n_666),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_750),
.A2(n_551),
.B(n_666),
.C(n_751),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_708),
.B(n_666),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_735),
.B(n_707),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_718),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_735),
.B(n_574),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_792),
.A2(n_666),
.B1(n_590),
.B2(n_591),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_726),
.A2(n_642),
.B(n_728),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_708),
.B(n_666),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_726),
.A2(n_642),
.B(n_728),
.Y(n_990)
);

AND2x6_ASAP7_75t_L g991 ( 
.A(n_763),
.B(n_639),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_708),
.B(n_666),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_708),
.B(n_666),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_772),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_890),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_982),
.B(n_930),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_866),
.A2(n_925),
.B(n_971),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_964),
.A2(n_951),
.B(n_954),
.C(n_869),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_981),
.B(n_983),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_887),
.A2(n_904),
.B(n_901),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_870),
.A2(n_958),
.B(n_884),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_958),
.A2(n_878),
.B(n_957),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_984),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_986),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_908),
.B(n_868),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_989),
.B(n_992),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_882),
.A2(n_883),
.B(n_949),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_921),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_922),
.A2(n_910),
.A3(n_865),
.B(n_918),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_950),
.A2(n_937),
.B1(n_952),
.B2(n_934),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_993),
.B(n_945),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_985),
.B(n_894),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_894),
.B(n_905),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_890),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_980),
.A2(n_987),
.B(n_969),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_950),
.B(n_956),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_864),
.B(n_920),
.C(n_897),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

CKINVDCx12_ASAP7_75t_R g1019 ( 
.A(n_937),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_985),
.B(n_900),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_893),
.B(n_886),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_905),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_915),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_960),
.B(n_967),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_941),
.B(n_940),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_863),
.B(n_896),
.Y(n_1026)
);

OAI22x1_ASAP7_75t_L g1027 ( 
.A1(n_912),
.A2(n_896),
.B1(n_880),
.B2(n_937),
.Y(n_1027)
);

NAND3x1_ASAP7_75t_L g1028 ( 
.A(n_902),
.B(n_975),
.C(n_871),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_963),
.A2(n_961),
.B(n_966),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_912),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_909),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_867),
.B(n_955),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_972),
.A2(n_938),
.B(n_935),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_946),
.A2(n_933),
.A3(n_965),
.B(n_931),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_909),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_899),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_SL g1037 ( 
.A1(n_924),
.A2(n_928),
.B(n_872),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_877),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_944),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_914),
.B(n_929),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_881),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_874),
.B(n_968),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_932),
.B(n_879),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_936),
.A2(n_939),
.A3(n_919),
.B(n_942),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_888),
.A2(n_973),
.B(n_891),
.C(n_947),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_953),
.B(n_903),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_973),
.A2(n_913),
.B(n_906),
.C(n_943),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_923),
.A2(n_898),
.A3(n_926),
.B(n_927),
.Y(n_1048)
);

AOI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_917),
.A2(n_977),
.B(n_976),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_911),
.B(n_916),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_873),
.A2(n_974),
.B(n_948),
.C(n_889),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_962),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_L g1053 ( 
.A1(n_902),
.A2(n_885),
.B1(n_979),
.B2(n_978),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_892),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_907),
.A2(n_970),
.B(n_892),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_875),
.A2(n_991),
.B1(n_994),
.B2(n_970),
.Y(n_1056)
);

AOI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_875),
.A2(n_949),
.B(n_964),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_991),
.A2(n_642),
.B(n_726),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_950),
.A2(n_937),
.B1(n_952),
.B2(n_934),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_958),
.B(n_864),
.C(n_920),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_984),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_890),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_890),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_930),
.A2(n_964),
.B(n_951),
.C(n_954),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_922),
.A2(n_959),
.A3(n_990),
.B(n_988),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_988),
.A2(n_642),
.B(n_726),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_922),
.A2(n_959),
.A3(n_990),
.B(n_988),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_908),
.B(n_574),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_982),
.B(n_930),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_921),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_984),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_890),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_982),
.B(n_930),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_890),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_950),
.A2(n_937),
.B1(n_952),
.B2(n_934),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_984),
.B(n_735),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_950),
.A2(n_937),
.B1(n_952),
.B2(n_934),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_908),
.A2(n_588),
.B(n_574),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_950),
.A2(n_937),
.B1(n_952),
.B2(n_934),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_981),
.B(n_983),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_981),
.B(n_983),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_894),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_984),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_L g1086 ( 
.A1(n_908),
.A2(n_588),
.B(n_574),
.Y(n_1086)
);

INVx3_ASAP7_75t_SL g1087 ( 
.A(n_984),
.Y(n_1087)
);

OA22x2_ASAP7_75t_L g1088 ( 
.A1(n_937),
.A2(n_950),
.B1(n_640),
.B2(n_620),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_930),
.A2(n_964),
.B(n_951),
.C(n_954),
.Y(n_1089)
);

CKINVDCx14_ASAP7_75t_R g1090 ( 
.A(n_984),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_988),
.A2(n_990),
.B(n_895),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_984),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_981),
.B(n_983),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_922),
.A2(n_959),
.A3(n_990),
.B(n_988),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_L g1096 ( 
.A(n_984),
.B(n_937),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_890),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_890),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_890),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_SL g1101 ( 
.A(n_984),
.B(n_566),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_890),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_984),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_908),
.B(n_574),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_L g1105 ( 
.A(n_864),
.B(n_879),
.C(n_908),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_981),
.B(n_983),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_958),
.B(n_864),
.C(n_920),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_930),
.A2(n_964),
.B(n_951),
.C(n_954),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_982),
.B(n_930),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_982),
.B(n_930),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_981),
.B(n_983),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_981),
.B(n_983),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_894),
.B(n_985),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_981),
.B(n_983),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_937),
.B(n_604),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_988),
.A2(n_990),
.B(n_959),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_984),
.B(n_735),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_890),
.Y(n_1119)
);

CKINVDCx6p67_ASAP7_75t_R g1120 ( 
.A(n_1036),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_999),
.B(n_1006),
.Y(n_1121)
);

CKINVDCx6p67_ASAP7_75t_R g1122 ( 
.A(n_1087),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1073),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1017),
.A2(n_1045),
.B(n_1011),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1096),
.B(n_1084),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1114),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1018),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_SL g1128 ( 
.A1(n_1010),
.A2(n_1077),
.B(n_1059),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1105),
.B(n_1005),
.C(n_1060),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_1111),
.B(n_1110),
.C(n_1071),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1103),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1078),
.B(n_1118),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1080),
.B(n_1086),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1088),
.A2(n_1116),
.B1(n_1016),
.B2(n_1059),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1091),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1016),
.A2(n_1075),
.B(n_996),
.C(n_1071),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1114),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1040),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_SL g1140 ( 
.A(n_1039),
.Y(n_1140)
);

AOI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1010),
.A2(n_1079),
.B(n_1077),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1088),
.A2(n_1104),
.B1(n_1070),
.B2(n_1025),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1000),
.A2(n_1065),
.B(n_1062),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1061),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_1084),
.B(n_1022),
.Y(n_1145)
);

AO21x2_ASAP7_75t_L g1146 ( 
.A1(n_1092),
.A2(n_1107),
.B(n_1099),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1090),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_1117),
.A2(n_997),
.B(n_1002),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1094),
.B(n_1106),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1112),
.B(n_1113),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1093),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1085),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_995),
.B(n_1014),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1002),
.A2(n_997),
.B(n_1068),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1081),
.A2(n_1041),
.B1(n_1116),
.B2(n_1037),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1003),
.Y(n_1156)
);

AOI222xp33_ASAP7_75t_L g1157 ( 
.A1(n_1027),
.A2(n_1053),
.B1(n_1115),
.B2(n_1024),
.C1(n_1021),
.C2(n_1101),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1116),
.B(n_1026),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1046),
.B(n_1030),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1019),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1063),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1064),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1041),
.A2(n_1119),
.B1(n_1100),
.B2(n_1102),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1097),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1098),
.B(n_1037),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1008),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1001),
.A2(n_1015),
.B(n_998),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1033),
.A2(n_1089),
.B(n_1109),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1004),
.B(n_1035),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_1072),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1032),
.B(n_1043),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1066),
.A2(n_1047),
.A3(n_1051),
.B(n_1058),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

OAI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1108),
.A2(n_1057),
.B1(n_1028),
.B2(n_1056),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1007),
.A2(n_1029),
.B(n_1055),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1049),
.A2(n_1057),
.B(n_1001),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1004),
.A2(n_1023),
.B1(n_1031),
.B2(n_1038),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1050),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1052),
.B(n_1050),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_1020),
.B(n_1012),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1054),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1067),
.A2(n_1095),
.B(n_1069),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1034),
.A2(n_1044),
.B(n_1067),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1069),
.A2(n_1044),
.B(n_1009),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1009),
.Y(n_1186)
);

NOR2xp67_ASAP7_75t_L g1187 ( 
.A(n_1048),
.B(n_1009),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1048),
.B(n_1034),
.Y(n_1188)
);

AND2x4_ASAP7_75t_SL g1189 ( 
.A(n_1044),
.B(n_894),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_999),
.B(n_1006),
.Y(n_1190)
);

BUFx2_ASAP7_75t_R g1191 ( 
.A(n_1008),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_1010),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1093),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1090),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1008),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1078),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1078),
.B(n_1118),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1005),
.B(n_908),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1096),
.B(n_894),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1090),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1078),
.B(n_1118),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1096),
.B(n_1013),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1136),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1171),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1142),
.B(n_1198),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1192),
.A2(n_1135),
.B1(n_1141),
.B2(n_1155),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1137),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1130),
.A2(n_1129),
.B(n_1124),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1172),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1169),
.A2(n_1184),
.B(n_1187),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1150),
.B(n_1135),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1150),
.B(n_1139),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1198),
.B(n_1196),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1132),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1128),
.A2(n_1192),
.B1(n_1138),
.B2(n_1126),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1197),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1201),
.B(n_1121),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1130),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1166),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1171),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1190),
.B(n_1146),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1151),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1146),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1186),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1189),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1148),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1183),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1151),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1126),
.B(n_1138),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1185),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1168),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1193),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1193),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1168),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1133),
.A2(n_1154),
.B(n_1143),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1196),
.B(n_1158),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1195),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1228),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1225),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1226),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1232),
.B(n_1188),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1223),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1232),
.B(n_1188),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1235),
.B(n_1188),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1219),
.B(n_1177),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1207),
.B(n_1133),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1231),
.B(n_1176),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1215),
.A2(n_1157),
.B(n_1178),
.Y(n_1250)
);

INVxp67_ASAP7_75t_SL g1251 ( 
.A(n_1203),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1227),
.B(n_1173),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1224),
.B(n_1173),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1234),
.B(n_1175),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1207),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1211),
.B(n_1175),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1211),
.A2(n_1202),
.B1(n_1147),
.B2(n_1131),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1218),
.B(n_1160),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1209),
.B(n_1164),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1243),
.B(n_1236),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1243),
.B(n_1210),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1255),
.B(n_1208),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1239),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1257),
.A2(n_1205),
.B1(n_1256),
.B2(n_1206),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1242),
.B(n_1214),
.Y(n_1265)
);

AND2x4_ASAP7_75t_SL g1266 ( 
.A(n_1241),
.B(n_1229),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1255),
.B(n_1208),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1243),
.B(n_1236),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1242),
.B(n_1209),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1245),
.B(n_1210),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1244),
.B(n_1216),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1240),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1248),
.B(n_1233),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1250),
.B(n_1194),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1250),
.B(n_1200),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1258),
.B(n_1122),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1251),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1244),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1261),
.B(n_1246),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1266),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1266),
.B(n_1257),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1263),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1272),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1260),
.B(n_1253),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1260),
.B(n_1253),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1265),
.B(n_1271),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1272),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1261),
.B(n_1249),
.Y(n_1289)
);

OR2x6_ASAP7_75t_SL g1290 ( 
.A(n_1271),
.B(n_1256),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1260),
.B(n_1253),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1265),
.B(n_1247),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1268),
.B(n_1252),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1268),
.B(n_1252),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1285),
.B(n_1273),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1284),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1287),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1283),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1287),
.B(n_1273),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1284),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1285),
.B(n_1264),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1283),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1288),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1281),
.B(n_1266),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1288),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1285),
.B(n_1261),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1286),
.B(n_1291),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1282),
.A2(n_1275),
.B1(n_1274),
.B2(n_1270),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1292),
.B(n_1279),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1308),
.A2(n_1290),
.B1(n_1281),
.B2(n_1280),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1298),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1306),
.B(n_1289),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1304),
.A2(n_1277),
.B(n_1281),
.C(n_1290),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1298),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1297),
.Y(n_1315)
);

AOI32xp33_ASAP7_75t_L g1316 ( 
.A1(n_1301),
.A2(n_1280),
.A3(n_1290),
.B1(n_1289),
.B2(n_1276),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1307),
.B(n_1286),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1302),
.Y(n_1318)
);

OAI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1306),
.A2(n_1280),
.B(n_1292),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1299),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1299),
.B(n_1286),
.Y(n_1321)
);

OAI21xp33_ASAP7_75t_L g1322 ( 
.A1(n_1295),
.A2(n_1309),
.B(n_1280),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1309),
.A2(n_1278),
.B(n_1269),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1296),
.A2(n_1261),
.B1(n_1270),
.B2(n_1289),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1296),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1300),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1311),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1325),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1311),
.Y(n_1329)
);

NOR3xp33_ASAP7_75t_SL g1330 ( 
.A(n_1313),
.B(n_1238),
.C(n_1221),
.Y(n_1330)
);

AOI21xp33_ASAP7_75t_L g1331 ( 
.A1(n_1310),
.A2(n_1248),
.B(n_1258),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1313),
.A2(n_1230),
.B(n_1178),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1323),
.B(n_1291),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1320),
.B(n_1291),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1316),
.A2(n_1319),
.B1(n_1322),
.B2(n_1312),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1315),
.A2(n_1321),
.B(n_1324),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1321),
.B(n_1293),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1333),
.B(n_1317),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1330),
.A2(n_1335),
.B1(n_1332),
.B2(n_1336),
.Y(n_1339)
);

OAI211xp5_ASAP7_75t_L g1340 ( 
.A1(n_1330),
.A2(n_1147),
.B(n_1259),
.C(n_1167),
.Y(n_1340)
);

OAI211xp5_ASAP7_75t_L g1341 ( 
.A1(n_1331),
.A2(n_1259),
.B(n_1167),
.C(n_1213),
.Y(n_1341)
);

OAI211xp5_ASAP7_75t_L g1342 ( 
.A1(n_1334),
.A2(n_1258),
.B(n_1164),
.C(n_1254),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1329),
.A2(n_1312),
.B(n_1326),
.Y(n_1343)
);

NAND4xp25_ASAP7_75t_L g1344 ( 
.A(n_1337),
.B(n_1237),
.C(n_1212),
.D(n_1206),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1328),
.A2(n_1326),
.B1(n_1312),
.B2(n_1318),
.C(n_1314),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1329),
.A2(n_1280),
.B1(n_1289),
.B2(n_1314),
.Y(n_1346)
);

AOI21xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1327),
.A2(n_1230),
.B(n_1204),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1332),
.A2(n_1289),
.B1(n_1270),
.B2(n_1318),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1338),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1339),
.B(n_1204),
.Y(n_1350)
);

AND4x1_ASAP7_75t_L g1351 ( 
.A(n_1348),
.B(n_1191),
.C(n_1204),
.D(n_1140),
.Y(n_1351)
);

OAI221xp5_ASAP7_75t_L g1352 ( 
.A1(n_1341),
.A2(n_1254),
.B1(n_1267),
.B2(n_1262),
.C(n_1269),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1340),
.B(n_1144),
.C(n_1123),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1346),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1345),
.B(n_1293),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1343),
.B(n_1293),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1344),
.B(n_1300),
.Y(n_1357)
);

AOI211x1_ASAP7_75t_L g1358 ( 
.A1(n_1351),
.A2(n_1342),
.B(n_1347),
.C(n_1303),
.Y(n_1358)
);

NOR2x1_ASAP7_75t_L g1359 ( 
.A(n_1350),
.B(n_1120),
.Y(n_1359)
);

NAND4xp25_ASAP7_75t_L g1360 ( 
.A(n_1350),
.B(n_1212),
.C(n_1220),
.D(n_1217),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1354),
.B(n_1152),
.C(n_1127),
.Y(n_1361)
);

NAND4xp75_ASAP7_75t_L g1362 ( 
.A(n_1349),
.B(n_1140),
.C(n_1170),
.D(n_1195),
.Y(n_1362)
);

NAND5xp2_ASAP7_75t_L g1363 ( 
.A(n_1353),
.B(n_1230),
.C(n_1199),
.D(n_1125),
.E(n_1220),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1357),
.B(n_1303),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1355),
.B(n_1305),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1356),
.B(n_1305),
.Y(n_1366)
);

NOR2x1_ASAP7_75t_L g1367 ( 
.A(n_1359),
.B(n_1352),
.Y(n_1367)
);

NOR3xp33_ASAP7_75t_L g1368 ( 
.A(n_1361),
.B(n_1362),
.C(n_1363),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_SL g1369 ( 
.A(n_1364),
.B(n_1353),
.C(n_1199),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1360),
.B(n_1180),
.C(n_1156),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1366),
.B(n_1217),
.Y(n_1371)
);

NOR4xp75_ASAP7_75t_L g1372 ( 
.A(n_1365),
.B(n_1262),
.C(n_1267),
.D(n_1241),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_L g1373 ( 
.A(n_1358),
.B(n_1179),
.Y(n_1373)
);

NOR2x1_ASAP7_75t_L g1374 ( 
.A(n_1359),
.B(n_1179),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1359),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1371),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1375),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1294),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1377),
.B(n_1373),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1377),
.B(n_1367),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1376),
.Y(n_1381)
);

OR3x1_ASAP7_75t_L g1382 ( 
.A(n_1379),
.B(n_1368),
.C(n_1372),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1380),
.A2(n_1378),
.B(n_1374),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1382),
.B(n_1381),
.Y(n_1384)
);

OAI22x1_ASAP7_75t_L g1385 ( 
.A1(n_1383),
.A2(n_1370),
.B1(n_1159),
.B2(n_1163),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1383),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1386),
.A2(n_1181),
.B(n_1182),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1384),
.A2(n_1125),
.B(n_1174),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1385),
.A2(n_1162),
.B(n_1161),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1388),
.A2(n_1163),
.B(n_1153),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1390),
.B(n_1387),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1391),
.A2(n_1389),
.B(n_1181),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1392),
.A2(n_1145),
.B1(n_1165),
.B2(n_1181),
.Y(n_1393)
);


endmodule