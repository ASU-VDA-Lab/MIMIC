module fake_jpeg_1125_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_21),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_43),
.B1(n_46),
.B2(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_64),
.B1(n_68),
.B2(n_50),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_69),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_50),
.B1(n_33),
.B2(n_2),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_33),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_15),
.C(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_3),
.B(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_74),
.C(n_77),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_12),
.B(n_23),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_11),
.B(n_22),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_86),
.B1(n_81),
.B2(n_88),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_16),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_96),
.B(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_93),
.Y(n_98)
);

OAI31xp33_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_90),
.A3(n_92),
.B(n_17),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_87),
.B(n_10),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_9),
.B1(n_20),
.B2(n_18),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_6),
.B1(n_25),
.B2(n_5),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_4),
.Y(n_104)
);


endmodule