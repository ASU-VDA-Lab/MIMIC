module fake_jpeg_26968_n_217 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_25),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_1),
.C(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_25),
.B1(n_16),
.B2(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_16),
.B1(n_24),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_27),
.B1(n_17),
.B2(n_5),
.Y(n_48)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_31),
.Y(n_52)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_37),
.B(n_41),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_57),
.B1(n_71),
.B2(n_75),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_30),
.B(n_31),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_76),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_61),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_31),
.C(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_67),
.Y(n_101)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

CKINVDCx11_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_36),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_37),
.B1(n_50),
.B2(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_36),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_36),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_37),
.A3(n_17),
.B1(n_41),
.B2(n_12),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_99),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_3),
.B(n_4),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_118),
.B1(n_92),
.B2(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_57),
.B1(n_68),
.B2(n_64),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_108),
.B1(n_120),
.B2(n_97),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_62),
.B1(n_76),
.B2(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_63),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_53),
.B1(n_45),
.B2(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_45),
.B1(n_4),
.B2(n_6),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_125),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_94),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_122),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_92),
.B1(n_98),
.B2(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_88),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_92),
.B1(n_98),
.B2(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_143),
.B(n_115),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_144),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_91),
.B(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_91),
.C(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_103),
.C(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_3),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_160),
.C(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_163),
.B1(n_152),
.B2(n_131),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_105),
.Y(n_158)
);

OA21x2_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_132),
.B(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_114),
.C(n_108),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_137),
.B1(n_157),
.B2(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_134),
.B1(n_142),
.B2(n_141),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_156),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_133),
.B1(n_144),
.B2(n_132),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_130),
.C(n_143),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_156),
.C(n_127),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_164),
.B(n_138),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_169),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_177),
.A2(n_149),
.B1(n_154),
.B2(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_172),
.B1(n_174),
.B2(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_165),
.B(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_176),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_101),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_193),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_174),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_197),
.C(n_3),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_187),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_126),
.B1(n_101),
.B2(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_101),
.B1(n_183),
.B2(n_7),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_203),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_196),
.B1(n_194),
.B2(n_197),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_192),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_10),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_202),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_210),
.B(n_208),
.C(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_203),
.C(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_206),
.C2(n_191),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_6),
.B(n_8),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_9),
.Y(n_217)
);


endmodule