module fake_jpeg_2944_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_61),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_55),
.Y(n_101)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_17),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_2),
.B(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_6),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_76),
.Y(n_94)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_18),
.B(n_7),
.CON(n_76),
.SN(n_76)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_90),
.B1(n_97),
.B2(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_109),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_24),
.B1(n_32),
.B2(n_29),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_99),
.B1(n_95),
.B2(n_87),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_41),
.A2(n_39),
.B1(n_24),
.B2(n_19),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_95),
.B1(n_81),
.B2(n_87),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_19),
.B1(n_36),
.B2(n_23),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_31),
.B1(n_35),
.B2(n_18),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_31),
.B1(n_18),
.B2(n_10),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_69),
.B1(n_52),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_18),
.B1(n_8),
.B2(n_10),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_108),
.B1(n_103),
.B2(n_79),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_42),
.B(n_18),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_96),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_94),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_130),
.C(n_136),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_7),
.B(n_8),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_121),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_7),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_120),
.B(n_126),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_92),
.B(n_89),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_125),
.B1(n_136),
.B2(n_121),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_79),
.Y(n_129)
);

CKINVDCx10_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_88),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_102),
.B1(n_82),
.B2(n_88),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_102),
.C(n_96),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_136),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_114),
.Y(n_140)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_143),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_144),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_112),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_115),
.B(n_109),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_161),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_134),
.C(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_139),
.B1(n_145),
.B2(n_154),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_165),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_170),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_117),
.A2(n_125),
.B(n_135),
.C(n_122),
.D(n_149),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_119),
.B1(n_133),
.B2(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_124),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_134),
.B(n_141),
.C(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_181),
.C(n_184),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_154),
.B1(n_168),
.B2(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_189),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_151),
.C(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_161),
.C(n_167),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_158),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_192),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_150),
.C(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_156),
.C(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_164),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_171),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_165),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_185),
.C(n_186),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_154),
.B1(n_171),
.B2(n_170),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_201),
.B1(n_184),
.B2(n_181),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_179),
.A2(n_182),
.B1(n_177),
.B2(n_178),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_172),
.B(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_172),
.B(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_208),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_211),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_213),
.B1(n_214),
.B2(n_205),
.Y(n_218)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_193),
.C(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_193),
.C(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.C(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_200),
.B(n_201),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_209),
.B(n_208),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_219),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_202),
.B1(n_210),
.B2(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_228),
.Y(n_229)
);

OAI31xp33_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_227),
.A3(n_222),
.B(n_206),
.Y(n_230)
);

AOI31xp67_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_175),
.A3(n_194),
.B(n_213),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_211),
.CI(n_214),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_189),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_211),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_229),
.B(n_223),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_228),
.B(n_231),
.C(n_207),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_230),
.B1(n_227),
.B2(n_236),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);


endmodule