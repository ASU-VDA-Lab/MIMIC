module fake_jpeg_28965_n_461 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_461);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_461;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_72),
.Y(n_142)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_78),
.Y(n_101)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_80),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_92),
.Y(n_154)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_99),
.Y(n_137)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_11),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_109),
.B(n_131),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_47),
.B1(n_53),
.B2(n_78),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_127),
.B1(n_138),
.B2(n_149),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_119),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_66),
.B(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_36),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_51),
.A2(n_29),
.B1(n_37),
.B2(n_41),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

BUFx4f_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_141),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_54),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g169 ( 
.A(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_45),
.B1(n_43),
.B2(n_33),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_58),
.A2(n_67),
.B1(n_63),
.B2(n_90),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_37),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_162),
.B(n_163),
.Y(n_234)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_29),
.B1(n_41),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_165),
.A2(n_177),
.B1(n_187),
.B2(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_22),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_22),
.Y(n_167)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_35),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_173),
.Y(n_221)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_34),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_93),
.C(n_80),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_153),
.C(n_120),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_34),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_179),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_110),
.A2(n_41),
.B1(n_14),
.B2(n_15),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_39),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_101),
.B1(n_151),
.B2(n_140),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_197),
.Y(n_238)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_124),
.B(n_28),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_142),
.B(n_28),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_24),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_24),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_0),
.B(n_3),
.Y(n_196)
);

INVx2_ASAP7_75t_R g197 ( 
.A(n_135),
.Y(n_197)
);

CKINVDCx12_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_135),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_119),
.Y(n_229)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_115),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_216),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_158),
.B1(n_126),
.B2(n_157),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_215),
.B(n_169),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_111),
.C(n_105),
.Y(n_223)
);

OA22x2_ASAP7_75t_SL g228 ( 
.A1(n_161),
.A2(n_144),
.B1(n_152),
.B2(n_102),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_235),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_175),
.A2(n_117),
.B1(n_103),
.B2(n_150),
.Y(n_232)
);

CKINVDCx9p33_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_170),
.Y(n_247)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_241),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_210),
.B(n_196),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_269),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_177),
.B(n_165),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_259),
.B(n_260),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_257),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_217),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_210),
.B(n_228),
.C(n_234),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_169),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_264),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_168),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_262),
.A2(n_263),
.B(n_227),
.Y(n_293)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_224),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_223),
.A2(n_219),
.B(n_226),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_226),
.B(n_225),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_199),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_218),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_285),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_238),
.C(n_222),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_282),
.C(n_295),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_238),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_244),
.A2(n_228),
.B1(n_216),
.B2(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_286),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_211),
.C(n_221),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_182),
.B1(n_120),
.B2(n_122),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_258),
.A2(n_153),
.B1(n_122),
.B2(n_134),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_292),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_134),
.B1(n_174),
.B2(n_101),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_259),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_220),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_252),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_220),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_257),
.C(n_267),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

XNOR2x1_ASAP7_75t_SL g304 ( 
.A(n_271),
.B(n_253),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_305),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_271),
.A2(n_260),
.B(n_254),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_288),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_242),
.Y(n_310)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_316),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_260),
.B(n_263),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_315),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_277),
.B(n_262),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_265),
.B(n_251),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_274),
.C(n_296),
.Y(n_322)
);

INVx6_ASAP7_75t_SL g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_243),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_292),
.B1(n_278),
.B2(n_287),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_288),
.A2(n_248),
.B(n_178),
.Y(n_321)
);

AO22x1_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_306),
.B1(n_317),
.B2(n_309),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_327),
.C(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_297),
.A2(n_280),
.B1(n_279),
.B2(n_284),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_338),
.B1(n_319),
.B2(n_321),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_282),
.C(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_294),
.C(n_291),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_329),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_275),
.C(n_287),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_334),
.C(n_336),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_275),
.C(n_283),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_318),
.C(n_305),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_283),
.C(n_249),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_311),
.C(n_303),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_297),
.A2(n_286),
.B1(n_289),
.B2(n_276),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_314),
.A2(n_276),
.B1(n_290),
.B2(n_246),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_340),
.A2(n_307),
.B1(n_320),
.B2(n_321),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_310),
.Y(n_347)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_341),
.A2(n_298),
.B1(n_301),
.B2(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_348),
.A2(n_355),
.B1(n_361),
.B2(n_362),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_341),
.B1(n_338),
.B2(n_340),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_308),
.B1(n_315),
.B2(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_304),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_370),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_264),
.Y(n_354)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_332),
.C(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_299),
.B1(n_311),
.B2(n_246),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_299),
.B1(n_245),
.B2(n_233),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_328),
.B(n_248),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_367),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_346),
.A2(n_245),
.B1(n_233),
.B2(n_250),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_368),
.Y(n_371)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_369),
.B(n_335),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_248),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_351),
.C(n_353),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_375),
.A2(n_351),
.B1(n_333),
.B2(n_324),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_360),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_337),
.B1(n_331),
.B2(n_322),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_209),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_356),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_363),
.Y(n_385)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_385),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_341),
.Y(n_388)
);

OAI321xp33_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_365),
.A3(n_349),
.B1(n_355),
.B2(n_361),
.C(n_348),
.Y(n_391)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_391),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_359),
.B(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_392),
.B(n_394),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_398),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_376),
.B(n_200),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_395),
.B(n_396),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_377),
.B(n_261),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_212),
.C(n_209),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_399),
.B(n_404),
.C(n_387),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_212),
.B(n_178),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_402),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_189),
.B(n_194),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_401),
.A2(n_389),
.B1(n_383),
.B2(n_381),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_231),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_419),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_405),
.A2(n_379),
.B1(n_371),
.B2(n_374),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_410),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_194),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_381),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_373),
.B1(n_388),
.B2(n_380),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_414),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_403),
.C(n_392),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_419),
.C(n_190),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_398),
.B(n_230),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_208),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_415),
.B(n_417),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_401),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_390),
.C(n_400),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_412),
.A2(n_390),
.B(n_402),
.Y(n_421)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_205),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_427),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_423),
.B(n_426),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_418),
.A2(n_407),
.B(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_409),
.A2(n_189),
.B(n_191),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_428),
.B(n_432),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_180),
.C(n_206),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_433),
.C(n_428),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_186),
.Y(n_432)
);

XOR2x2_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_201),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_119),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_148),
.B1(n_140),
.B2(n_151),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_436),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_130),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_206),
.C(n_172),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_202),
.C(n_25),
.Y(n_450)
);

OAI221xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_15),
.B1(n_125),
.B2(n_11),
.C(n_113),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_443),
.A2(n_202),
.B(n_114),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_431),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_445),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_437),
.A2(n_427),
.B(n_11),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_446),
.A2(n_440),
.B(n_441),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_150),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_447),
.A2(n_442),
.B(n_436),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_448),
.B(n_450),
.Y(n_452)
);

AOI322xp5_ASAP7_75t_L g456 ( 
.A1(n_453),
.A2(n_454),
.A3(n_438),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_3),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_449),
.C(n_447),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_455),
.A2(n_456),
.B(n_452),
.Y(n_457)
);

AOI322xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_453),
.C2(n_454),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_8),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_460),
.Y(n_461)
);


endmodule