module fake_netlist_6_1408_n_126 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_126);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_126;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_100;
wire n_121;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_10),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_2),
.Y(n_54)
);

NAND3x1_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.C(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_1),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_3),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_8),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_4),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_4),
.Y(n_67)
);

NOR2x1p5_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_34),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_43),
.Y(n_76)
);

XNOR2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_43),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_63),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_64),
.Y(n_82)
);

AO21x2_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_47),
.B(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_61),
.B(n_64),
.C(n_63),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_67),
.B(n_56),
.C(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_42),
.B(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_45),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_56),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_73),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_36),
.Y(n_94)
);

OR2x6_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_55),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_R g98 ( 
.A(n_91),
.B(n_9),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

OAI31xp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_86),
.A3(n_84),
.B(n_91),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_92),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_95),
.B1(n_88),
.B2(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_96),
.B1(n_88),
.B2(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_101),
.B(n_83),
.Y(n_115)
);

OAI221xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_95),
.B1(n_82),
.B2(n_107),
.C(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_55),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_116),
.B1(n_95),
.B2(n_87),
.Y(n_121)
);

AOI31xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_51),
.A3(n_91),
.B(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_85),
.B1(n_81),
.B2(n_83),
.Y(n_123)
);

AOI31xp33_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_81),
.A3(n_83),
.B(n_11),
.Y(n_124)
);

XOR2x1_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_81),
.Y(n_125)
);

OAI221xp5_ASAP7_75t_R g126 ( 
.A1(n_125),
.A2(n_124),
.B1(n_123),
.B2(n_15),
.C(n_89),
.Y(n_126)
);


endmodule