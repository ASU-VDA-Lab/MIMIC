module fake_jpeg_5286_n_142 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx2_ASAP7_75t_SL g50 ( 
.A(n_33),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_6),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_43),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_10),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_31),
.B1(n_26),
.B2(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_62),
.B1(n_31),
.B2(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_51),
.B(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_69),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_43),
.C(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_58),
.B1(n_55),
.B2(n_48),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_44),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_43),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_63),
.C(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_85),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_57),
.B1(n_35),
.B2(n_13),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_60),
.C(n_67),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_69),
.B1(n_72),
.B2(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_90),
.B1(n_35),
.B2(n_15),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_12),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_65),
.B1(n_46),
.B2(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_85),
.A3(n_81),
.B1(n_65),
.B2(n_42),
.C1(n_75),
.C2(n_83),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_11),
.B1(n_33),
.B2(n_24),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_30),
.C(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_106),
.C(n_12),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_21),
.B(n_12),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_108),
.B(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_33),
.B1(n_34),
.B2(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_94),
.B(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_115),
.B1(n_34),
.B2(n_5),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_97),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_106),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_116),
.C(n_0),
.Y(n_122)
);

AOI31xp67_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_88),
.A3(n_12),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_5),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_123),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_105),
.C(n_100),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_122),
.B(n_4),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_98),
.B1(n_104),
.B2(n_20),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_124),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_34),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_109),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_111),
.B(n_112),
.C(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_7),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_123),
.A3(n_4),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_8),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_8),
.B1(n_3),
.B2(n_1),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_137),
.B(n_3),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_132),
.C(n_126),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_140),
.Y(n_142)
);


endmodule