module fake_jpeg_28954_n_31 (n_0, n_3, n_2, n_1, n_31);

input n_0;
input n_3;
input n_2;
input n_1;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_4;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g4 ( 
.A(n_3),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_1),
.Y(n_5)
);

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g9 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_10),
.Y(n_13)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_10),
.A2(n_7),
.B1(n_5),
.B2(n_4),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_13),
.B(n_4),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_9),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_19),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_15),
.B(n_11),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_10),
.B(n_8),
.Y(n_23)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_9),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_8),
.C(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_28),
.B(n_3),
.Y(n_31)
);


endmodule