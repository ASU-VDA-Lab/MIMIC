module fake_netlist_1_6347_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
BUFx3_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
AOI31xp67_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .A3(n_2), .B(n_1), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_4), .B1(n_3), .B2(n_9), .Y(n_13) );
OAI21xp33_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_11), .B(n_9), .Y(n_14) );
NAND3x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_12), .C(n_7), .Y(n_15) );
NOR2x1_ASAP7_75t_L g16 ( .A(n_14), .B(n_7), .Y(n_16) );
OR3x1_ASAP7_75t_L g17 ( .A(n_15), .B(n_2), .C(n_0), .Y(n_17) );
OAI21xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_16), .B(n_6), .Y(n_18) );
endmodule