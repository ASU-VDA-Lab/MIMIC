module fake_jpeg_31320_n_119 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_23),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_24),
.B1(n_23),
.B2(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_49),
.B1(n_36),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_17),
.B1(n_15),
.B2(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_39),
.Y(n_67)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_61),
.B1(n_43),
.B2(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_21),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_40),
.B1(n_47),
.B2(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_43),
.B1(n_38),
.B2(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_13),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_53),
.B1(n_40),
.B2(n_38),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_64),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_88),
.B(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_12),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_55),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_70),
.C(n_71),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_68),
.B(n_78),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_80),
.C(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_92),
.B1(n_97),
.B2(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_102),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_110),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_95),
.B(n_76),
.Y(n_110)
);

AOI31xp33_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_106),
.A3(n_4),
.B(n_3),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_4),
.A3(n_8),
.B1(n_9),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_72),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_113),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_116),
.Y(n_119)
);


endmodule