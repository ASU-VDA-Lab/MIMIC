module real_jpeg_12210_n_16 (n_5, n_4, n_8, n_0, n_12, n_272, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_272;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_29),
.B1(n_32),
.B2(n_45),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_71),
.B1(n_72),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_132),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_132),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_132),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_53),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_31),
.B1(n_71),
.B2(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_7),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_70),
.B(n_71),
.C(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_10),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_81),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_148),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_99),
.B1(n_100),
.B2(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_10),
.B(n_87),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_71),
.B1(n_72),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_157),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_157),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_13),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_36),
.B1(n_71),
.B2(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_71),
.B1(n_72),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_79),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_79),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_79),
.Y(n_230)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_19),
.B(n_113),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_83),
.B2(n_112),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_66),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_22),
.A2(n_23),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_26),
.A2(n_99),
.B(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_27),
.A2(n_37),
.B1(n_123),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_37),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_28),
.A2(n_37),
.B(n_125),
.Y(n_201)
);

CKINVDCx6p67_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_32),
.B(n_49),
.C(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_32),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_33),
.A2(n_100),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_50),
.B(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_42),
.A2(n_56),
.B(n_198),
.C(n_200),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_42),
.B(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_43),
.B(n_57),
.C(n_59),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_52),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_46),
.A2(n_91),
.B(n_104),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_46),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_46),
.A2(n_51),
.B1(n_205),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_51),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_46),
.A2(n_51),
.B1(n_213),
.B2(n_223),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_50),
.B(n_148),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_66),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_61),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_55),
.A2(n_152),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_60),
.B1(n_70),
.B2(n_75),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_59),
.A2(n_75),
.B(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g199 ( 
.A(n_60),
.B(n_148),
.CON(n_199),
.SN(n_199)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_62),
.A2(n_87),
.B1(n_151),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_62),
.A2(n_87),
.B1(n_186),
.B2(n_199),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_77),
.B(n_80),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_67),
.A2(n_76),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_78),
.B1(n_81),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_68),
.A2(n_81),
.B1(n_156),
.B2(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_69)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_96),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_128),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_90),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_99),
.A2(n_100),
.B1(n_228),
.B2(n_236),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_100),
.B(n_148),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_118),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_119),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_126),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_130),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_265),
.B(n_270),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_174),
.B1(n_190),
.B2(n_264),
.C(n_272),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_138),
.B(n_163),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_159),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_160),
.C(n_161),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_154),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_141),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_173),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_175),
.B(n_188),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_176),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_178),
.B(n_180),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.C(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_263),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_258),
.B(n_262),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_214),
.B(n_257),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_209),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_194),
.B(n_209),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_206),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_196),
.B(n_202),
.C(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_201),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_212),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_252),
.B(n_256),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_242),
.B(n_251),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_231),
.B(n_241),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_224),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.B(n_240),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_247),
.C(n_250),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);


endmodule