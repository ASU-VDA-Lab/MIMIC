module fake_jpeg_27854_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_32),
.B1(n_19),
.B2(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_25),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g107 ( 
.A(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_16),
.B(n_22),
.C(n_19),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_36),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_86),
.Y(n_117)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_32),
.B1(n_19),
.B2(n_20),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_32),
.B1(n_13),
.B2(n_9),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_34),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_41),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_24),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_55),
.B1(n_51),
.B2(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_16),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_34),
.CI(n_41),
.CON(n_103),
.SN(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_97),
.A2(n_99),
.B(n_104),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_105),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_31),
.Y(n_109)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_112),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_66),
.B(n_84),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_78),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_67),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_119),
.B(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_80),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_131),
.B(n_135),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_71),
.B1(n_73),
.B2(n_70),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_100),
.B1(n_97),
.B2(n_96),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_66),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_92),
.Y(n_157)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_97),
.B(n_102),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_16),
.B(n_4),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_62),
.B1(n_83),
.B2(n_72),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_112),
.B1(n_62),
.B2(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_143),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_77),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_82),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_87),
.C(n_74),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_22),
.C(n_5),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_171),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_90),
.B1(n_108),
.B2(n_104),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_162),
.B1(n_176),
.B2(n_139),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_92),
.B1(n_72),
.B2(n_85),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_121),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_131),
.B1(n_130),
.B2(n_133),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_110),
.B(n_91),
.C(n_88),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_165),
.B(n_170),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_110),
.B1(n_63),
.B2(n_56),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_63),
.B(n_59),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_153),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_77),
.B1(n_106),
.B2(n_59),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_31),
.C(n_16),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_16),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_3),
.B(n_4),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_179),
.B(n_4),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_22),
.B1(n_10),
.B2(n_11),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_141),
.B(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_188),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_204),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_125),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_195),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_126),
.C(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_202),
.C(n_201),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_158),
.B1(n_148),
.B2(n_150),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_145),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_140),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_176),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_171),
.C(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_128),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_154),
.C(n_149),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_220),
.C(n_193),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_177),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_191),
.B1(n_208),
.B2(n_204),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_148),
.C(n_153),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_175),
.B(n_165),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_230),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_152),
.B1(n_166),
.B2(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_123),
.B1(n_10),
.B2(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_183),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_249),
.Y(n_256)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_187),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_202),
.C(n_195),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_248),
.C(n_254),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_216),
.B1(n_215),
.B2(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_192),
.C(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_182),
.B1(n_194),
.B2(n_199),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_203),
.B1(n_200),
.B2(n_180),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_207),
.B(n_185),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_227),
.B(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_225),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_211),
.C(n_220),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_269),
.B(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_211),
.C(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_251),
.C(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_254),
.C(n_244),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_238),
.B(n_222),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_240),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_241),
.B(n_253),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_267),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_221),
.B(n_232),
.C(n_180),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_212),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_276),
.C(n_281),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_235),
.C(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_246),
.C(n_252),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_239),
.C(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_243),
.C(n_226),
.Y(n_279)
);

BUFx4f_ASAP7_75t_SL g280 ( 
.A(n_263),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_284),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_231),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_255),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_8),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_269),
.C(n_260),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_263),
.B1(n_269),
.B2(n_256),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_269),
.B1(n_257),
.B2(n_262),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_123),
.C(n_9),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_278),
.B(n_280),
.Y(n_298)
);

AOI31xp33_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_287),
.A3(n_15),
.B(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_303),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_292),
.B(n_297),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_8),
.B(n_12),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_306),
.B(n_13),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_12),
.B(n_13),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_307),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_308),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_15),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_15),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_309),
.C(n_313),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_315),
.A3(n_300),
.B1(n_7),
.B2(n_6),
.C(n_5),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_5),
.B(n_6),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_7),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_300),
.Y(n_321)
);


endmodule