module fake_jpeg_2518_n_408 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_52),
.B(n_57),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_85),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_33),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_80),
.Y(n_101)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_88),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_1),
.C(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_3),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_90),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_19),
.A2(n_3),
.B(n_4),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_44),
.Y(n_130)
);

INVx2_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_100),
.B(n_112),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_37),
.B1(n_34),
.B2(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_104),
.A2(n_124),
.B1(n_106),
.B2(n_105),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_87),
.B1(n_67),
.B2(n_34),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_108),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_58),
.A2(n_97),
.B1(n_94),
.B2(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_109),
.A2(n_118),
.B1(n_149),
.B2(n_111),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_42),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_28),
.B1(n_32),
.B2(n_45),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_117),
.B1(n_32),
.B2(n_96),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_32),
.B1(n_45),
.B2(n_31),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_34),
.B1(n_31),
.B2(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_37),
.B1(n_44),
.B2(n_32),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_83),
.B1(n_76),
.B2(n_73),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_21),
.B(n_39),
.C(n_38),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_127),
.B(n_128),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_21),
.B(n_39),
.C(n_38),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_22),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_50),
.B(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_51),
.B(n_36),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_154),
.Y(n_233)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_17),
.B(n_95),
.C(n_32),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_113),
.B(n_150),
.C(n_103),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_177),
.B1(n_182),
.B2(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_125),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_172),
.B1(n_180),
.B2(n_193),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_121),
.B1(n_140),
.B2(n_101),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_175),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_68),
.B1(n_65),
.B2(n_37),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_179),
.B1(n_190),
.B2(n_106),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_35),
.B1(n_29),
.B2(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_35),
.B1(n_29),
.B2(n_23),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_101),
.A2(n_22),
.B1(n_17),
.B2(n_53),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_4),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_189),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_101),
.A2(n_122),
.B1(n_137),
.B2(n_132),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_100),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_186),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_12),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_12),
.B1(n_141),
.B2(n_147),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_195),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_198),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_110),
.B(n_133),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_119),
.B(n_99),
.Y(n_218)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_110),
.B1(n_129),
.B2(n_145),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_129),
.B1(n_110),
.B2(n_124),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_206),
.B1(n_208),
.B2(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_162),
.B1(n_173),
.B2(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_105),
.B1(n_144),
.B2(n_145),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_144),
.B1(n_102),
.B2(n_119),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_223),
.B1(n_183),
.B2(n_148),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_218),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_99),
.C(n_123),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_230),
.C(n_176),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_156),
.A2(n_172),
.B1(n_170),
.B2(n_178),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_136),
.B1(n_139),
.B2(n_142),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_123),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_136),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_139),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_170),
.A2(n_103),
.B(n_148),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_158),
.B(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

BUFx4f_ASAP7_75t_SL g235 ( 
.A(n_205),
.Y(n_235)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_204),
.B(n_169),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_236),
.B(n_241),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_160),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_209),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_192),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_249),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_210),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_188),
.C(n_174),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_164),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_214),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_227),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_181),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_251),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_180),
.B1(n_191),
.B2(n_155),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_260),
.B1(n_202),
.B2(n_218),
.Y(n_265)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_223),
.A2(n_198),
.B1(n_139),
.B2(n_142),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_258),
.B1(n_207),
.B2(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_163),
.B(n_194),
.C(n_154),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_221),
.B(n_231),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_202),
.A2(n_213),
.B1(n_199),
.B2(n_215),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_171),
.B1(n_142),
.B2(n_134),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_134),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_200),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_237),
.B1(n_253),
.B2(n_259),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_225),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_268),
.B(n_274),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_273),
.A2(n_240),
.B(n_257),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_214),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_220),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_275),
.B(n_279),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_220),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_257),
.B(n_255),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_307),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_290),
.A2(n_305),
.B(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_237),
.B1(n_239),
.B2(n_253),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_253),
.B1(n_258),
.B2(n_243),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_306),
.B(n_291),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_252),
.B1(n_238),
.B2(n_236),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_280),
.C(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_301),
.C(n_302),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_213),
.B1(n_260),
.B2(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_299),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_247),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_246),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_303),
.B(n_309),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_273),
.B(n_266),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_232),
.B1(n_248),
.B2(n_234),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_272),
.A2(n_232),
.B1(n_199),
.B2(n_242),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_200),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_254),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_283),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_318),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_283),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_285),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_323),
.B(n_333),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_273),
.B(n_276),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_284),
.B(n_262),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_325),
.A2(n_326),
.B(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_232),
.B(n_265),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_277),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_300),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_331),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_286),
.B(n_277),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_286),
.B(n_277),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_263),
.C(n_235),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_292),
.C(n_293),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_338),
.C(n_342),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_293),
.C(n_289),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_318),
.C(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_296),
.C(n_295),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_298),
.B1(n_294),
.B2(n_300),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_345),
.A2(n_329),
.B1(n_321),
.B2(n_325),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_296),
.C(n_308),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_278),
.C(n_269),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.Y(n_359)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_235),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_322),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_361),
.B1(n_338),
.B2(n_337),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_326),
.C(n_312),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_354),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_343),
.A2(n_316),
.B1(n_329),
.B2(n_294),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_355),
.A2(n_360),
.B1(n_344),
.B2(n_346),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_347),
.A2(n_320),
.B(n_315),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_357),
.A2(n_287),
.B(n_272),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_316),
.B1(n_331),
.B2(n_314),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_341),
.A2(n_312),
.B1(n_332),
.B2(n_320),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_349),
.Y(n_368)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_366),
.B(n_281),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_336),
.B(n_347),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_233),
.B(n_229),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_358),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_369),
.A2(n_370),
.B1(n_377),
.B2(n_360),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_SL g371 ( 
.A1(n_356),
.A2(n_262),
.A3(n_342),
.B1(n_348),
.B2(n_281),
.C1(n_278),
.C2(n_211),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_371),
.B(n_376),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_373),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_361),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_375),
.A2(n_287),
.B1(n_262),
.B2(n_233),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_363),
.B(n_348),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_355),
.A2(n_287),
.B1(n_254),
.B2(n_199),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_364),
.C(n_359),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_380),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_359),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_381),
.A2(n_386),
.B1(n_228),
.B2(n_205),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_364),
.Y(n_382)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_362),
.C(n_365),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_228),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_387),
.A2(n_367),
.B(n_373),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_368),
.C(n_375),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_390),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_394),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_383),
.A2(n_377),
.B1(n_229),
.B2(n_222),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_230),
.Y(n_400)
);

OAI211xp5_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_385),
.B(n_379),
.C(n_386),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_399),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_393),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_389),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_391),
.C(n_388),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_403),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_401),
.A2(n_398),
.B(n_395),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_222),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_405),
.B(n_201),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_201),
.Y(n_408)
);


endmodule