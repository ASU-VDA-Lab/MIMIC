module fake_netlist_5_2126_n_1814 (n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_48, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_1814);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_1814;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_82;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_111;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_105;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_87;
wire n_150;
wire n_1728;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_51;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_101;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_94;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_59;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_72;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1561;
wire n_1267;
wire n_1165;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_114;
wire n_96;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_129;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_49;
wire n_310;
wire n_54;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_70;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_91;
wire n_1565;
wire n_1809;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_117;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1538;
wire n_272;
wire n_1162;
wire n_1199;
wire n_1779;
wire n_352;
wire n_53;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_71;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_121;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_64;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_103;
wire n_97;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_52;
wire n_784;
wire n_110;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_61;
wire n_678;
wire n_697;
wire n_127;
wire n_1222;
wire n_75;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_116;
wire n_1710;
wire n_284;
wire n_1128;
wire n_139;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_100;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_133;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_106;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_93;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_122;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_90;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_123;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_131;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_109;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_88;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_65;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_69;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_73;
wire n_309;
wire n_512;
wire n_1591;
wire n_84;
wire n_130;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_112;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_55;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_102;
wire n_77;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_83;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_58;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_128;
wire n_120;
wire n_327;
wire n_135;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_62;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_86;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_74;
wire n_1139;
wire n_515;
wire n_57;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_132;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_50;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_107;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_149;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_85;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_118;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_108;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_66;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_126;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_89;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_115;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_137;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_124;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_119;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_67;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_68;
wire n_867;
wire n_186;
wire n_134;
wire n_587;
wire n_63;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_138;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_95;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_104;
wire n_682;
wire n_1567;
wire n_56;
wire n_141;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_140;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_78;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_98;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_80;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_92;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_79;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_76;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_81;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_60;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_113;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_99;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_0),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_22),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_21),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_17),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_6),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_51),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_63),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_56),
.B1(n_62),
.B2(n_72),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_63),
.B(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_72),
.Y(n_123)
);

AOI21x1_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_64),
.B(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_108),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_54),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_54),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_71),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_114),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_52),
.B(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_58),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_55),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_109),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_107),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_121),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_58),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_110),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_R g180 ( 
.A(n_146),
.B(n_110),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

AND3x1_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_87),
.C(n_75),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_117),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_135),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_129),
.B(n_130),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_113),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_129),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_R g208 ( 
.A(n_134),
.B(n_113),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_130),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_130),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_130),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_130),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_156),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_130),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_107),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_111),
.Y(n_234)
);

NAND2x1p5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_141),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_111),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_132),
.Y(n_245)
);

NAND3x1_ASAP7_75t_L g246 ( 
.A(n_170),
.B(n_86),
.C(n_69),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_200),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_148),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_191),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_194),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_144),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_153),
.B(n_134),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_69),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

BUFx4f_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_175),
.B(n_141),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_176),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_161),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_154),
.B(n_70),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_180),
.B(n_128),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_159),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

BUFx6f_ASAP7_75t_SL g282 ( 
.A(n_177),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_166),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_202),
.B(n_204),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_166),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_162),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_209),
.B(n_128),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_205),
.B(n_177),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_164),
.B(n_70),
.Y(n_290)
);

OR2x6_ASAP7_75t_L g291 ( 
.A(n_169),
.B(n_145),
.Y(n_291)
);

INVx4_ASAP7_75t_SL g292 ( 
.A(n_177),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_181),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_168),
.B(n_80),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_174),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_174),
.A2(n_120),
.B1(n_132),
.B2(n_141),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_174),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_184),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_171),
.B(n_109),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_147),
.B(n_74),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_183),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_185),
.B(n_144),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_172),
.A2(n_67),
.B1(n_74),
.B2(n_93),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_147),
.B(n_80),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_186),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_147),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_161),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_147),
.B(n_144),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_195),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_195),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_221),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_211),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_139),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_212),
.Y(n_322)
);

AO22x2_ASAP7_75t_L g323 ( 
.A1(n_233),
.A2(n_67),
.B1(n_86),
.B2(n_84),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_219),
.A2(n_120),
.B1(n_95),
.B2(n_77),
.Y(n_324)
);

NAND2x1p5_ASAP7_75t_L g325 ( 
.A(n_244),
.B(n_128),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_251),
.B(n_56),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_212),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_215),
.A2(n_90),
.B(n_75),
.C(n_93),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_62),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_213),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_226),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_219),
.B(n_132),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_226),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_213),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_253),
.B(n_59),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_224),
.Y(n_339)
);

AO22x2_ASAP7_75t_L g340 ( 
.A1(n_233),
.A2(n_84),
.B1(n_87),
.B2(n_90),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_216),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_220),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_214),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_296),
.B(n_120),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_139),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_222),
.B(n_132),
.Y(n_348)
);

AO22x2_ASAP7_75t_L g349 ( 
.A1(n_253),
.A2(n_145),
.B1(n_120),
.B2(n_61),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_234),
.A2(n_120),
.B1(n_79),
.B2(n_132),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_247),
.B(n_139),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_217),
.A2(n_128),
.B1(n_144),
.B2(n_120),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_247),
.B(n_142),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_220),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_252),
.B(n_61),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_120),
.B1(n_132),
.B2(n_140),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_222),
.B(n_120),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_222),
.B(n_142),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_236),
.B(n_142),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_262),
.B(n_135),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_223),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_244),
.B(n_128),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_223),
.Y(n_363)
);

BUFx4f_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_228),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_249),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_244),
.B(n_128),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_275),
.B(n_71),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_228),
.Y(n_369)
);

OAI221xp5_ASAP7_75t_L g370 ( 
.A1(n_225),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_225),
.B(n_83),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_236),
.B(n_142),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_280),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_250),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_290),
.B(n_97),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_214),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_237),
.A2(n_97),
.B(n_142),
.C(n_133),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_250),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_247),
.B(n_217),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_258),
.B(n_92),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_281),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_247),
.B(n_124),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_260),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_260),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_283),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_244),
.B(n_128),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_243),
.Y(n_391)
);

NAND2x1p5_ASAP7_75t_L g392 ( 
.A(n_244),
.B(n_128),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_243),
.B(n_91),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_283),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_284),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_217),
.B(n_128),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_284),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_261),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_261),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_232),
.B(n_128),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_264),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_294),
.B(n_76),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_264),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_302),
.Y(n_405)
);

BUFx4f_ASAP7_75t_L g406 ( 
.A(n_291),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_227),
.B(n_124),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_227),
.B(n_124),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_293),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_312),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_227),
.B(n_124),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_285),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_317),
.A2(n_262),
.B(n_313),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx3_ASAP7_75t_SL g415 ( 
.A(n_341),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_317),
.A2(n_262),
.B(n_255),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_291),
.B1(n_218),
.B2(n_214),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_336),
.B(n_293),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_291),
.C(n_245),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_348),
.A2(n_255),
.B(n_232),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_336),
.B(n_301),
.Y(n_421)
);

O2A1O1Ixp5_ASAP7_75t_L g422 ( 
.A1(n_364),
.A2(n_305),
.B(n_257),
.C(n_288),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_237),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_238),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_358),
.B(n_357),
.Y(n_425)
);

O2A1O1Ixp33_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_303),
.B(n_301),
.C(n_307),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_333),
.A2(n_255),
.B(n_232),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_326),
.B(n_329),
.C(n_393),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_346),
.A2(n_242),
.B1(n_238),
.B2(n_241),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_321),
.B(n_257),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_321),
.B(n_347),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_347),
.B(n_257),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_360),
.A2(n_255),
.B(n_232),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_346),
.A2(n_242),
.B1(n_241),
.B2(n_267),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_360),
.A2(n_214),
.B(n_271),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_330),
.B(n_257),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_407),
.A2(n_271),
.B(n_268),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

AOI22x1_ASAP7_75t_L g443 ( 
.A1(n_349),
.A2(n_230),
.B1(n_231),
.B2(n_270),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_326),
.B(n_301),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_372),
.A2(n_303),
.B(n_307),
.C(n_289),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_329),
.B(n_307),
.Y(n_447)
);

O2A1O1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_372),
.A2(n_303),
.B(n_230),
.C(n_231),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_338),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_381),
.A2(n_265),
.B(n_270),
.Y(n_450)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_351),
.Y(n_451)
);

BUFx12f_ASAP7_75t_L g452 ( 
.A(n_373),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_335),
.B(n_259),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_342),
.B(n_259),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_338),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_393),
.B(n_78),
.C(n_81),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_375),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_328),
.A2(n_230),
.B(n_231),
.C(n_306),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_407),
.A2(n_268),
.B(n_256),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_402),
.B(n_304),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_344),
.B(n_259),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_351),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_366),
.B(n_248),
.Y(n_464)
);

AOI21xp33_ASAP7_75t_L g465 ( 
.A1(n_349),
.A2(n_304),
.B(n_246),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_408),
.A2(n_268),
.B(n_256),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_354),
.Y(n_467)
);

AND2x2_ASAP7_75t_SL g468 ( 
.A(n_364),
.B(n_406),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_361),
.B(n_259),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_363),
.B(n_259),
.Y(n_471)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_369),
.B(n_239),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_408),
.A2(n_268),
.B(n_256),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_334),
.B(n_248),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_368),
.B(n_304),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_411),
.A2(n_256),
.B(n_271),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_345),
.A2(n_218),
.B1(n_259),
.B2(n_282),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_411),
.A2(n_268),
.B(n_256),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_379),
.B(n_304),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_353),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_400),
.A2(n_271),
.B(n_314),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_345),
.B(n_380),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_400),
.A2(n_271),
.B(n_314),
.Y(n_485)
);

CKINVDCx10_ASAP7_75t_R g486 ( 
.A(n_318),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_380),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_406),
.A2(n_240),
.B(n_239),
.C(n_269),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_367),
.A2(n_269),
.B(n_274),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_365),
.B(n_263),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_315),
.B(n_240),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_L g492 ( 
.A1(n_328),
.A2(n_306),
.B(n_263),
.C(n_267),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_316),
.B(n_319),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_318),
.B(n_235),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_320),
.B(n_273),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_386),
.B(n_309),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_367),
.A2(n_273),
.B(n_274),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_359),
.A2(n_311),
.B(n_298),
.C(n_277),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_331),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_385),
.B(n_272),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_322),
.B(n_265),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_327),
.B(n_399),
.Y(n_502)
);

AOI21xp33_ASAP7_75t_L g503 ( 
.A1(n_349),
.A2(n_246),
.B(n_311),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_399),
.B(n_218),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

NOR2x1p5_ASAP7_75t_SL g507 ( 
.A(n_401),
.B(n_278),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_374),
.A2(n_235),
.B(n_309),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_337),
.B(n_259),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_325),
.A2(n_235),
.B(n_309),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_376),
.A2(n_282),
.B1(n_254),
.B2(n_297),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_337),
.B(n_218),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_401),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_355),
.A2(n_218),
.B1(n_282),
.B2(n_300),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_248),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_324),
.A2(n_218),
.B1(n_300),
.B2(n_272),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_325),
.A2(n_254),
.B(n_276),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_362),
.A2(n_254),
.B(n_151),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_323),
.B(n_248),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_350),
.A2(n_218),
.B1(n_300),
.B2(n_272),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_389),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_362),
.A2(n_151),
.B(n_310),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_403),
.B(n_272),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_371),
.B(n_295),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_377),
.B(n_295),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_403),
.B(n_310),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_394),
.B(n_405),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_395),
.B(n_292),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_397),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_390),
.A2(n_310),
.B(n_277),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_390),
.A2(n_392),
.B(n_352),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_522),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_429),
.A2(n_447),
.B1(n_445),
.B2(n_418),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g536 ( 
.A(n_468),
.B(n_356),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_448),
.A2(n_404),
.B(n_388),
.C(n_387),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_412),
.B(n_323),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_SL g539 ( 
.A(n_435),
.B(n_382),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_432),
.A2(n_436),
.B1(n_417),
.B2(n_423),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_423),
.B(n_323),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_484),
.B(n_340),
.Y(n_546)
);

CKINVDCx6p67_ASAP7_75t_R g547 ( 
.A(n_486),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g548 ( 
.A1(n_511),
.A2(n_378),
.B(n_376),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_484),
.B(n_340),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_476),
.B(n_340),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_480),
.B(n_376),
.Y(n_552)
);

O2A1O1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_465),
.A2(n_279),
.B(n_278),
.C(n_286),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_427),
.A2(n_392),
.B(n_396),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_310),
.Y(n_555)
);

OAI21xp33_ASAP7_75t_SL g556 ( 
.A1(n_528),
.A2(n_279),
.B(n_286),
.Y(n_556)
);

AO21x1_ASAP7_75t_L g557 ( 
.A1(n_511),
.A2(n_298),
.B(n_297),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_437),
.A2(n_396),
.B(n_119),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_SL g559 ( 
.A(n_465),
.B(n_118),
.C(n_300),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_451),
.B(n_292),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_421),
.A2(n_300),
.B1(n_292),
.B2(n_140),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_440),
.B(n_300),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_467),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_428),
.B(n_433),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_469),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_415),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_431),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_420),
.A2(n_118),
.B(n_292),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_512),
.B(n_138),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_300),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_509),
.B(n_138),
.Y(n_575)
);

O2A1O1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_426),
.A2(n_133),
.B(n_137),
.C(n_126),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_517),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_517),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_456),
.B(n_135),
.C(n_138),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_434),
.B(n_2),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g584 ( 
.A(n_494),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

O2A1O1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_446),
.A2(n_133),
.B(n_137),
.C(n_126),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_419),
.A2(n_133),
.B(n_137),
.C(n_126),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_487),
.B(n_433),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_464),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_439),
.A2(n_118),
.B(n_137),
.Y(n_592)
);

AO31x2_ASAP7_75t_L g593 ( 
.A1(n_438),
.A2(n_137),
.A3(n_126),
.B(n_135),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_499),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_594)
);

O2A1O1Ixp5_ASAP7_75t_L g595 ( 
.A1(n_422),
.A2(n_126),
.B(n_135),
.C(n_133),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_SL g596 ( 
.A(n_503),
.B(n_7),
.C(n_8),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_473),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_433),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_475),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_413),
.A2(n_138),
.B(n_133),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_416),
.A2(n_479),
.B(n_459),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_481),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_441),
.A2(n_138),
.B(n_133),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_487),
.B(n_135),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_520),
.B(n_8),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_458),
.A2(n_138),
.B(n_125),
.C(n_12),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_514),
.B(n_138),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_482),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_466),
.A2(n_138),
.B(n_135),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_515),
.B(n_9),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_424),
.B(n_430),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_516),
.B(n_138),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_501),
.B(n_9),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_474),
.A2(n_125),
.B(n_38),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_500),
.A2(n_140),
.B1(n_125),
.B2(n_15),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_451),
.B(n_140),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_463),
.B(n_10),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_477),
.A2(n_125),
.B(n_42),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_425),
.A2(n_125),
.B(n_40),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_495),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_424),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_495),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_490),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_430),
.A2(n_125),
.B1(n_16),
.B2(n_17),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_501),
.B(n_140),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_482),
.Y(n_630)
);

BUFx2_ASAP7_75t_SL g631 ( 
.A(n_463),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_490),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_SL g633 ( 
.A1(n_425),
.A2(n_140),
.B(n_36),
.C(n_34),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_503),
.A2(n_140),
.B1(n_125),
.B2(n_19),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_483),
.A2(n_125),
.B(n_33),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_485),
.A2(n_508),
.B(n_523),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_450),
.A2(n_519),
.B(n_438),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_451),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_496),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_444),
.B(n_140),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_450),
.A2(n_510),
.B(n_532),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_463),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_524),
.A2(n_140),
.B1(n_125),
.B2(n_23),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

OAI21x1_ASAP7_75t_SL g646 ( 
.A1(n_492),
.A2(n_12),
.B(n_18),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_488),
.A2(n_125),
.B(n_140),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_478),
.A2(n_125),
.B1(n_28),
.B2(n_29),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_444),
.A2(n_140),
.B1(n_31),
.B2(n_32),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_140),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_SL g651 ( 
.A(n_504),
.B(n_25),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_491),
.A2(n_32),
.B1(n_140),
.B2(n_521),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_504),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_518),
.A2(n_140),
.B(n_531),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_453),
.B(n_140),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_SL g656 ( 
.A(n_454),
.B(n_462),
.C(n_470),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_SL g657 ( 
.A(n_471),
.B(n_489),
.C(n_497),
.Y(n_657)
);

OAI22x1_ASAP7_75t_L g658 ( 
.A1(n_443),
.A2(n_472),
.B1(n_529),
.B2(n_507),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_529),
.B(n_429),
.C(n_384),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_498),
.A2(n_429),
.B1(n_435),
.B2(n_445),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_429),
.A2(n_384),
.B(n_445),
.C(n_234),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_427),
.A2(n_437),
.B(n_420),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_429),
.A2(n_384),
.B(n_445),
.C(n_447),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_560),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_624),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_541),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_569),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_560),
.Y(n_671)
);

INVx6_ASAP7_75t_L g672 ( 
.A(n_630),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_638),
.Y(n_674)
);

CKINVDCx6p67_ASAP7_75t_R g675 ( 
.A(n_547),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_544),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_549),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_641),
.B(n_637),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_630),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_549),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_630),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_566),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_632),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_572),
.B(n_575),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_662),
.A2(n_636),
.B(n_601),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_585),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_579),
.B(n_608),
.Y(n_689)
);

BUFx2_ASAP7_75t_SL g690 ( 
.A(n_567),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_597),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_656),
.B(n_654),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_618),
.Y(n_693)
);

INVx6_ASAP7_75t_SL g694 ( 
.A(n_565),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_630),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_593),
.Y(n_696)
);

CKINVDCx11_ASAP7_75t_R g697 ( 
.A(n_590),
.Y(n_697)
);

BUFx2_ASAP7_75t_SL g698 ( 
.A(n_577),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_568),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_627),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_573),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_599),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_540),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_642),
.Y(n_706)
);

NAND2x1p5_ASAP7_75t_L g707 ( 
.A(n_572),
.B(n_575),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_589),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_589),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_543),
.B(n_551),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_563),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_533),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_563),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_598),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_598),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_591),
.B(n_639),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_612),
.A2(n_536),
.B1(n_659),
.B2(n_594),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_602),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_536),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_550),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_545),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_591),
.B(n_639),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_564),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_645),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_573),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_578),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_631),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_603),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_587),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_578),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_623),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_644),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_653),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_640),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_625),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_626),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_535),
.B(n_663),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_614),
.B(n_609),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_584),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_619),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_653),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_593),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_538),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_605),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_537),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_615),
.Y(n_750)
);

BUFx4f_ASAP7_75t_SL g751 ( 
.A(n_609),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_615),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_593),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_612),
.A2(n_620),
.B1(n_606),
.B2(n_542),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_613),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_553),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_655),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_661),
.A2(n_634),
.B1(n_652),
.B2(n_552),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_574),
.Y(n_759)
);

INVx5_ASAP7_75t_L g760 ( 
.A(n_633),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_629),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_595),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_556),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_633),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_595),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_614),
.B(n_651),
.Y(n_766)
);

BUFx4_ASAP7_75t_SL g767 ( 
.A(n_581),
.Y(n_767)
);

INVx8_ASAP7_75t_L g768 ( 
.A(n_539),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_658),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_559),
.Y(n_770)
);

BUFx4f_ASAP7_75t_SL g771 ( 
.A(n_582),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_548),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_660),
.Y(n_774)
);

INVx6_ASAP7_75t_SL g775 ( 
.A(n_596),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_557),
.B(n_634),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_648),
.A2(n_628),
.B1(n_622),
.B2(n_617),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_562),
.Y(n_778)
);

BUFx2_ASAP7_75t_SL g779 ( 
.A(n_616),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_650),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_582),
.B(n_596),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_554),
.B(n_621),
.Y(n_782)
);

INVx6_ASAP7_75t_L g783 ( 
.A(n_559),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_717),
.A2(n_649),
.B1(n_643),
.B2(n_657),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_740),
.A2(n_657),
.B1(n_635),
.B2(n_592),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_754),
.A2(n_561),
.B1(n_647),
.B2(n_558),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_781),
.A2(n_607),
.B1(n_588),
.B2(n_571),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_735),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_687),
.A2(n_576),
.B(n_586),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_692),
.A2(n_600),
.B(n_611),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_773),
.A2(n_604),
.B1(n_758),
.B2(n_752),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_738),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_692),
.A2(n_762),
.B(n_765),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_664),
.A2(n_696),
.B(n_753),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_773),
.A2(n_771),
.B1(n_751),
.B2(n_750),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_736),
.Y(n_796)
);

OAI21x1_ASAP7_75t_SL g797 ( 
.A1(n_774),
.A2(n_777),
.B(n_772),
.Y(n_797)
);

NOR2x1_ASAP7_75t_R g798 ( 
.A(n_697),
.B(n_690),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_762),
.A2(n_765),
.B(n_745),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_683),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_679),
.A2(n_755),
.B(n_782),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_763),
.A2(n_745),
.B(n_753),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_668),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_664),
.A2(n_696),
.B(n_769),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_669),
.Y(n_805)
);

CKINVDCx9p33_ASAP7_75t_R g806 ( 
.A(n_738),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_670),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_769),
.A2(n_766),
.B(n_757),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_673),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_677),
.Y(n_810)
);

AOI21x1_ASAP7_75t_L g811 ( 
.A1(n_756),
.A2(n_749),
.B(n_782),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_676),
.B(n_716),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_704),
.A2(n_743),
.B1(n_742),
.B2(n_783),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_683),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_689),
.B(n_685),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_774),
.B(n_768),
.Y(n_817)
);

BUFx4_ASAP7_75t_SL g818 ( 
.A(n_742),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_783),
.A2(n_735),
.B1(n_775),
.B2(n_743),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_782),
.B(n_768),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_SL g821 ( 
.A1(n_776),
.A2(n_734),
.B(n_759),
.C(n_676),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_726),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_679),
.B(n_749),
.C(n_747),
.Y(n_823)
);

INVx6_ASAP7_75t_L g824 ( 
.A(n_680),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_671),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_757),
.A2(n_766),
.B(n_676),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_739),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_678),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_695),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_776),
.A2(n_749),
.B(n_684),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_760),
.A2(n_764),
.B(n_730),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_760),
.A2(n_764),
.B(n_691),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_775),
.A2(n_783),
.B1(n_770),
.B2(n_780),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_766),
.A2(n_757),
.B(n_707),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_700),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_695),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_739),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_686),
.A2(n_707),
.B(n_741),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_675),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_744),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_689),
.B(n_780),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_697),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_693),
.B(n_666),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_719),
.B(n_721),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_695),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_744),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_686),
.A2(n_707),
.B(n_741),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_679),
.A2(n_782),
.B(n_768),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_775),
.A2(n_770),
.B1(n_783),
.B2(n_743),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_671),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_686),
.A2(n_741),
.B(n_666),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_688),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_768),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_779),
.B(n_778),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_693),
.B(n_710),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_719),
.B(n_721),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_718),
.A2(n_701),
.B(n_682),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_701),
.A2(n_682),
.B(n_779),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_710),
.B(n_746),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_681),
.A2(n_747),
.B(n_748),
.C(n_706),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_746),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_695),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_725),
.B(n_748),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_760),
.A2(n_764),
.B(n_703),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_770),
.A2(n_725),
.B1(n_720),
.B2(n_761),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_682),
.A2(n_760),
.B(n_764),
.Y(n_867)
);

OAI221xp5_ASAP7_75t_L g868 ( 
.A1(n_690),
.A2(n_743),
.B1(n_712),
.B2(n_761),
.C(n_729),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_739),
.Y(n_869)
);

AOI222xp33_ASAP7_75t_L g870 ( 
.A1(n_770),
.A2(n_725),
.B1(n_761),
.B2(n_737),
.C1(n_739),
.C2(n_732),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_760),
.A2(n_764),
.B(n_778),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_727),
.A2(n_728),
.B(n_723),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_725),
.A2(n_720),
.B1(n_761),
.B2(n_737),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_671),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_720),
.A2(n_761),
.B1(n_737),
.B2(n_778),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_727),
.A2(n_728),
.B(n_711),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_733),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_778),
.A2(n_671),
.B(n_720),
.Y(n_878)
);

AO31x2_ASAP7_75t_L g879 ( 
.A1(n_720),
.A2(n_778),
.A3(n_767),
.B(n_733),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_SL g880 ( 
.A(n_675),
.B(n_667),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_671),
.A2(n_720),
.B(n_737),
.Y(n_881)
);

INVx6_ASAP7_75t_L g882 ( 
.A(n_680),
.Y(n_882)
);

CKINVDCx11_ASAP7_75t_R g883 ( 
.A(n_667),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_720),
.A2(n_737),
.B(n_665),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_716),
.A2(n_723),
.B(n_711),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_665),
.A2(n_731),
.B(n_680),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_712),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_726),
.B(n_716),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_804),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_802),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_807),
.B(n_702),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_838),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_804),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_802),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_885),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_794),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_794),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_790),
.A2(n_793),
.B(n_811),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_839),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_794),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_858),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_858),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_872),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_872),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_872),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_799),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_792),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_830),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_830),
.Y(n_909)
);

OAI22xp33_ASAP7_75t_L g910 ( 
.A1(n_813),
.A2(n_726),
.B1(n_732),
.B2(n_724),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_792),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_793),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_885),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_871),
.B(n_680),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_853),
.Y(n_915)
);

AOI222xp33_ASAP7_75t_L g916 ( 
.A1(n_784),
.A2(n_726),
.B1(n_722),
.B2(n_724),
.C1(n_674),
.C2(n_723),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_801),
.A2(n_713),
.B(n_731),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_798),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_803),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_862),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_859),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_820),
.A2(n_713),
.B(n_680),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_805),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_859),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_838),
.B(n_731),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_885),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_784),
.A2(n_702),
.B1(n_665),
.B2(n_722),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_851),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_823),
.A2(n_665),
.B1(n_709),
.B2(n_708),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_851),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_791),
.A2(n_665),
.B1(n_698),
.B2(n_674),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_810),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_853),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_852),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_791),
.A2(n_698),
.B1(n_709),
.B2(n_708),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_834),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_834),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_826),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_808),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_808),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_847),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_855),
.B(n_860),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_840),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

CKINVDCx12_ASAP7_75t_R g945 ( 
.A(n_818),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_846),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_886),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_878),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_833),
.A2(n_699),
.B1(n_705),
.B2(n_731),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_878),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_843),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_815),
.B(n_731),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_815),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_844),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_827),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_827),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_806),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_837),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_837),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_806),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_869),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_821),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_797),
.A2(n_673),
.B1(n_694),
.B2(n_714),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_821),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_796),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_816),
.B(n_695),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_848),
.A2(n_699),
.B(n_705),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_714),
.B1(n_715),
.B2(n_672),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_831),
.A2(n_832),
.B(n_871),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_833),
.A2(n_699),
.B1(n_705),
.B2(n_672),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_884),
.B(n_881),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_842),
.A2(n_694),
.B1(n_715),
.B2(n_672),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_884),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_831),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_832),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_881),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_865),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_857),
.B(n_715),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_854),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_979),
.B(n_812),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_945),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_931),
.A2(n_787),
.B1(n_786),
.B2(n_842),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_979),
.B(n_812),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_954),
.B(n_835),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_899),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_919),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_913),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_957),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_954),
.B(n_856),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_947),
.B(n_812),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_978),
.B(n_864),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_R g992 ( 
.A(n_957),
.B(n_865),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_965),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_978),
.B(n_942),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_864),
.Y(n_995)
);

NOR2x1p5_ASAP7_75t_L g996 ( 
.A(n_942),
.B(n_887),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_SL g997 ( 
.A(n_916),
.B(n_861),
.C(n_868),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_966),
.B(n_828),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_967),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_965),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_891),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_952),
.B(n_788),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_966),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_919),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_960),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_952),
.Y(n_1006)
);

AOI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_931),
.A2(n_849),
.B(n_819),
.C(n_880),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_920),
.B(n_877),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_895),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_R g1010 ( 
.A(n_960),
.B(n_865),
.Y(n_1010)
);

BUFx5_ASAP7_75t_L g1011 ( 
.A(n_889),
.Y(n_1011)
);

CKINVDCx16_ASAP7_75t_R g1012 ( 
.A(n_952),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_914),
.B(n_817),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_920),
.B(n_888),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_951),
.B(n_841),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_951),
.B(n_822),
.Y(n_1016)
);

NAND2x1p5_ASAP7_75t_L g1017 ( 
.A(n_922),
.B(n_853),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_968),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_923),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_967),
.B(n_839),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_947),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_961),
.B(n_809),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_914),
.B(n_817),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_943),
.B(n_876),
.Y(n_1024)
);

CKINVDCx6p67_ASAP7_75t_R g1025 ( 
.A(n_918),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_947),
.B(n_879),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_923),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_927),
.A2(n_963),
.B1(n_929),
.B2(n_968),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_943),
.B(n_875),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_953),
.B(n_854),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_953),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_935),
.A2(n_785),
.B1(n_883),
.B2(n_870),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_R g1034 ( 
.A(n_917),
.B(n_817),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_935),
.A2(n_853),
.B1(n_887),
.B2(n_824),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_956),
.B(n_809),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_SL g1037 ( 
.A(n_963),
.B(n_825),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_956),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_925),
.B(n_879),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_932),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_910),
.A2(n_970),
.B(n_972),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_916),
.A2(n_785),
.B1(n_883),
.B2(n_866),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_910),
.A2(n_866),
.B1(n_854),
.B2(n_873),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_946),
.B(n_875),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_958),
.Y(n_1046)
);

NOR2x1p5_ASAP7_75t_L g1047 ( 
.A(n_915),
.B(n_800),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_962),
.A2(n_882),
.B1(n_824),
.B2(n_825),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_958),
.B(n_873),
.Y(n_1049)
);

CKINVDCx16_ASAP7_75t_R g1050 ( 
.A(n_925),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_SL g1051 ( 
.A(n_962),
.B(n_825),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_922),
.B(n_882),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_934),
.B(n_879),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_972),
.B(n_882),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_970),
.A2(n_800),
.B1(n_814),
.B2(n_694),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_915),
.B(n_824),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_914),
.B(n_874),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_R g1058 ( 
.A(n_917),
.B(n_886),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_934),
.Y(n_1059)
);

NOR2x1p5_ASAP7_75t_L g1060 ( 
.A(n_915),
.B(n_814),
.Y(n_1060)
);

AND2x4_ASAP7_75t_SL g1061 ( 
.A(n_915),
.B(n_814),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_898),
.A2(n_867),
.B(n_790),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_955),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_925),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_SL g1065 ( 
.A(n_964),
.B(n_874),
.C(n_850),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_913),
.Y(n_1066)
);

BUFx4f_ASAP7_75t_SL g1067 ( 
.A(n_933),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_959),
.B(n_879),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_895),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_959),
.B(n_800),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_907),
.Y(n_1071)
);

AO21x2_ASAP7_75t_L g1072 ( 
.A1(n_974),
.A2(n_867),
.B(n_789),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_955),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_907),
.B(n_814),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_SL g1075 ( 
.A(n_964),
.B(n_874),
.C(n_850),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_955),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_911),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_971),
.B(n_800),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_933),
.B(n_829),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_911),
.Y(n_1080)
);

INVx8_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1012),
.B(n_971),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_1009),
.Y(n_1083)
);

OAI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_982),
.A2(n_938),
.B1(n_950),
.B2(n_908),
.C(n_909),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1009),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1050),
.B(n_926),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1064),
.B(n_971),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1030),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1077),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1078),
.B(n_895),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_994),
.B(n_926),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_991),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1039),
.B(n_950),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_982),
.A2(n_949),
.B1(n_892),
.B2(n_908),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1039),
.B(n_950),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_995),
.B(n_977),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1021),
.B(n_977),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1005),
.B(n_948),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_990),
.B(n_948),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1080),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1076),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1026),
.B(n_948),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_975),
.B(n_974),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1073),
.B(n_905),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1052),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1026),
.B(n_948),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_990),
.B(n_976),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_984),
.B(n_976),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1014),
.B(n_909),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1011),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_989),
.B(n_976),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_997),
.A2(n_949),
.B1(n_892),
.B2(n_917),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1002),
.B(n_973),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_980),
.B(n_983),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_987),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_980),
.B(n_973),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1052),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_987),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_998),
.B(n_1003),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1011),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_983),
.B(n_973),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1066),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1069),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1053),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_1066),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_903),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1081),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1011),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1017),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1017),
.A2(n_898),
.B(n_975),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1069),
.B(n_904),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1049),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1015),
.B(n_905),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1079),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1033),
.B(n_892),
.C(n_904),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_988),
.B(n_938),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_988),
.B(n_938),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_986),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1011),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1022),
.B(n_892),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1068),
.B(n_892),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1013),
.B(n_892),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1032),
.B(n_889),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1067),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1016),
.B(n_917),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1036),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1063),
.B(n_893),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1079),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1013),
.B(n_969),
.Y(n_1149)
);

INVxp67_ASAP7_75t_SL g1150 ( 
.A(n_992),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_1028),
.A2(n_917),
.B1(n_933),
.B2(n_914),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1057),
.B(n_940),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1081),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_933),
.B1(n_850),
.B2(n_940),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1013),
.B(n_969),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_L g1156 ( 
.A(n_981),
.B(n_715),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1004),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1019),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1081),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1027),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1023),
.B(n_1057),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1040),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1024),
.B(n_1008),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1044),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1059),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1011),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1023),
.B(n_939),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1071),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1023),
.B(n_969),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1038),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1011),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1031),
.B(n_893),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_993),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1000),
.B(n_944),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_999),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1029),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1047),
.B(n_939),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_999),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1070),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_999),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1046),
.B(n_1001),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_999),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1060),
.B(n_944),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1020),
.B(n_969),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_1045),
.B(n_898),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1020),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1018),
.A2(n_944),
.B1(n_941),
.B2(n_937),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1051),
.B(n_941),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1074),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1072),
.B(n_941),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1072),
.B(n_902),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1062),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1062),
.Y(n_1194)
);

AOI31xp33_ASAP7_75t_L g1195 ( 
.A1(n_1035),
.A2(n_937),
.A3(n_936),
.B(n_897),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1192),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_992),
.B1(n_1010),
.B2(n_1034),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1169),
.Y(n_1198)
);

NAND2x1_ASAP7_75t_L g1199 ( 
.A(n_1105),
.B(n_900),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1192),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1176),
.A2(n_897),
.A3(n_900),
.B(n_937),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1130),
.A2(n_896),
.B(n_936),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1087),
.B(n_996),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1087),
.B(n_1035),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1132),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1144),
.Y(n_1206)
);

OAI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1151),
.A2(n_1007),
.B1(n_1033),
.B2(n_1037),
.C(n_1042),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1182),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1135),
.A2(n_1037),
.B1(n_1042),
.B2(n_1025),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1144),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1089),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1177),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1187),
.A2(n_985),
.B1(n_1010),
.B2(n_1056),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1130),
.A2(n_896),
.B(n_936),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1169),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1135),
.A2(n_1048),
.B(n_1043),
.C(n_1055),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1191),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1129),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1150),
.A2(n_1054),
.B1(n_1056),
.B2(n_1067),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1089),
.Y(n_1220)
);

OAI211xp5_ASAP7_75t_L g1221 ( 
.A1(n_1112),
.A2(n_1084),
.B(n_1154),
.C(n_1094),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1134),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1177),
.B(n_1055),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1176),
.A2(n_1075),
.B(n_1065),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1105),
.A2(n_1043),
.B1(n_1054),
.B2(n_1075),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1182),
.B(n_1061),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1082),
.B(n_1048),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1103),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1191),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1129),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1129),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1175),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1175),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_1065),
.B(n_896),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1161),
.A2(n_1034),
.B1(n_1058),
.B2(n_924),
.Y(n_1235)
);

OAI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1188),
.A2(n_930),
.B(n_928),
.C(n_921),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1181),
.A2(n_930),
.B(n_928),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1143),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1193),
.A2(n_930),
.B(n_928),
.Y(n_1239)
);

NAND4xp25_ASAP7_75t_L g1240 ( 
.A(n_1117),
.B(n_1058),
.C(n_924),
.D(n_921),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1138),
.Y(n_1241)
);

AOI21xp33_ASAP7_75t_L g1242 ( 
.A1(n_1195),
.A2(n_1117),
.B(n_1185),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1143),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1134),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1129),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1193),
.A2(n_902),
.B(n_901),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1195),
.A2(n_829),
.B1(n_845),
.B2(n_863),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1161),
.A2(n_902),
.B1(n_901),
.B2(n_906),
.Y(n_1248)
);

AND2x6_ASAP7_75t_L g1249 ( 
.A(n_1166),
.B(n_863),
.Y(n_1249)
);

INVx4_ASAP7_75t_R g1250 ( 
.A(n_1127),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1138),
.Y(n_1251)
);

AOI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1185),
.A2(n_894),
.B1(n_890),
.B2(n_912),
.C(n_906),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1163),
.B(n_906),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1147),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1179),
.A2(n_1062),
.B(n_912),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1148),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1157),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1147),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1100),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1156),
.A2(n_894),
.B(n_890),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1144),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1082),
.B(n_1141),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1141),
.B(n_845),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1100),
.Y(n_1265)
);

OAI211xp5_ASAP7_75t_L g1266 ( 
.A1(n_1103),
.A2(n_715),
.B(n_836),
.C(n_863),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1148),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1104),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1109),
.A2(n_789),
.B(n_699),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1099),
.B(n_836),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1171),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1157),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1088),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1190),
.B(n_1180),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1166),
.B(n_836),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1099),
.B(n_836),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1129),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1179),
.A2(n_863),
.B(n_672),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1183),
.A2(n_699),
.A3(n_705),
.B(n_1110),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1158),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1145),
.A2(n_705),
.B(n_1103),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1129),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1124),
.B(n_1173),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1119),
.A2(n_1133),
.B(n_1144),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1178),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1104),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1166),
.B(n_1142),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1096),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1142),
.B1(n_1178),
.B2(n_1126),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1272),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1237),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1272),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1204),
.B(n_1093),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1250),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1280),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1244),
.B(n_1183),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1204),
.B(n_1093),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1227),
.B(n_1263),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1280),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1227),
.B(n_1095),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1208),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1245),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_1244),
.Y(n_1304)
);

OAI211xp5_ASAP7_75t_L g1305 ( 
.A1(n_1221),
.A2(n_1149),
.B(n_1170),
.C(n_1155),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1263),
.B(n_1095),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1208),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1242),
.A2(n_1194),
.B(n_1193),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1223),
.B(n_1190),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1207),
.A2(n_1086),
.B1(n_1146),
.B2(n_1178),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1290),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1213),
.B(n_1106),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1209),
.A2(n_1168),
.B1(n_1152),
.B2(n_1186),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1222),
.B(n_1106),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1290),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1168),
.B1(n_1152),
.B2(n_1186),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1197),
.A2(n_1170),
.B1(n_1155),
.B2(n_1149),
.C(n_1092),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1283),
.B(n_1268),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1283),
.B(n_1186),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1262),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1198),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1215),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1273),
.B(n_1096),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1237),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1222),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1256),
.Y(n_1326)
);

AND2x4_ASAP7_75t_SL g1327 ( 
.A(n_1203),
.B(n_1210),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1206),
.A2(n_1168),
.B1(n_1152),
.B2(n_1186),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1241),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1287),
.B(n_1256),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1237),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1251),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1212),
.B(n_1091),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1257),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1287),
.B(n_1106),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1228),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1287),
.B(n_1106),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1271),
.Y(n_1338)
);

OAI221xp5_ASAP7_75t_L g1339 ( 
.A1(n_1235),
.A2(n_1216),
.B1(n_1219),
.B2(n_1225),
.C(n_1240),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1211),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1267),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1268),
.B(n_1186),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1267),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1211),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1260),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1245),
.B(n_1183),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1285),
.B(n_1102),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1285),
.B(n_1102),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1201),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1205),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1284),
.B(n_1091),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1274),
.B(n_1108),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1220),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1288),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1271),
.B(n_1153),
.Y(n_1355)
);

NAND4xp25_ASAP7_75t_L g1356 ( 
.A(n_1289),
.B(n_1086),
.C(n_1179),
.D(n_1097),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1201),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1220),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1286),
.B(n_1173),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1203),
.B(n_1102),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1286),
.B(n_1238),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1210),
.A2(n_1178),
.B1(n_1153),
.B2(n_1127),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1206),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1259),
.Y(n_1364)
);

OR2x2_ASAP7_75t_SL g1365 ( 
.A(n_1206),
.B(n_1101),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1245),
.B(n_1199),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1226),
.B(n_1114),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1281),
.A2(n_1194),
.B(n_1128),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1201),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1259),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1206),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1264),
.B(n_1108),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_SL g1373 ( 
.A(n_1224),
.B(n_1159),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1265),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1265),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1238),
.B(n_1122),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1277),
.B(n_1102),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1210),
.A2(n_1168),
.B1(n_1152),
.B2(n_1126),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1295),
.B(n_1299),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1291),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1366),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_L g1383 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1320),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1338),
.B(n_1304),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1320),
.B(n_1114),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1293),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1330),
.B(n_1282),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1341),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1330),
.B(n_1282),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1296),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1300),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1312),
.B(n_1218),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1312),
.B(n_1218),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1326),
.B(n_1253),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1320),
.B(n_1264),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1327),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1327),
.B(n_1245),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1311),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1355),
.B(n_1245),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1294),
.B(n_1218),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1315),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1341),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1318),
.B(n_1243),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1294),
.B(n_1230),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1302),
.B(n_1097),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1340),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1307),
.B(n_1243),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

AOI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1305),
.A2(n_1252),
.B1(n_1247),
.B2(n_1236),
.C(n_1266),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1350),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1344),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1325),
.B(n_1254),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1318),
.B(n_1254),
.Y(n_1414)
);

AND2x2_ASAP7_75t_SL g1415 ( 
.A(n_1308),
.B(n_1230),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_L g1416 ( 
.A(n_1343),
.B(n_1199),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1353),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1358),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1309),
.B(n_1258),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1354),
.B(n_1258),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1298),
.B(n_1230),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1298),
.B(n_1231),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1301),
.B(n_1232),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1301),
.B(n_1231),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1360),
.B(n_1231),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1364),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1295),
.B(n_1232),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1365),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1343),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1370),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1336),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1339),
.A2(n_1269),
.B1(n_1249),
.B2(n_1224),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1360),
.B(n_1276),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1335),
.B(n_1337),
.Y(n_1434)
);

NAND4xp25_ASAP7_75t_L g1435 ( 
.A(n_1317),
.B(n_1313),
.C(n_1310),
.D(n_1356),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1374),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1323),
.B(n_1233),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1336),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1345),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1335),
.B(n_1337),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1361),
.B(n_1233),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1362),
.B(n_1276),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1306),
.B(n_1270),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1363),
.B(n_1248),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1306),
.B(n_1314),
.Y(n_1445)
);

AND2x4_ASAP7_75t_SL g1446 ( 
.A(n_1314),
.B(n_1275),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1384),
.B(n_1363),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1434),
.B(n_1371),
.Y(n_1448)
);

NAND2xp67_ASAP7_75t_L g1449 ( 
.A(n_1385),
.B(n_1345),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1408),
.B(n_1411),
.Y(n_1450)
);

NOR3xp33_ASAP7_75t_L g1451 ( 
.A(n_1384),
.B(n_1303),
.C(n_1371),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1381),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1381),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1380),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1434),
.B(n_1297),
.Y(n_1455)
);

AOI32xp33_ASAP7_75t_L g1456 ( 
.A1(n_1428),
.A2(n_1351),
.A3(n_1328),
.B1(n_1348),
.B2(n_1347),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1387),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1429),
.B(n_1321),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1440),
.B(n_1297),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1387),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1391),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1413),
.B(n_1365),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_1379),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1384),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1383),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_L g1466 ( 
.A(n_1383),
.B(n_1297),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1322),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1391),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1431),
.B(n_1329),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1392),
.Y(n_1471)
);

NAND4xp25_ASAP7_75t_L g1472 ( 
.A(n_1435),
.B(n_1316),
.C(n_1378),
.D(n_1319),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1423),
.B(n_1361),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1397),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1392),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1398),
.B(n_1303),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1386),
.B(n_1367),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1379),
.B(n_1377),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1399),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1399),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1446),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1427),
.B(n_1395),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1398),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1419),
.B(n_1333),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1398),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1402),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1438),
.B(n_1332),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1389),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1393),
.B(n_1377),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1389),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1446),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1445),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1402),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1407),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1407),
.Y(n_1495)
);

NAND4xp25_ASAP7_75t_L g1496 ( 
.A(n_1432),
.B(n_1319),
.C(n_1342),
.D(n_1346),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1437),
.B(n_1352),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1406),
.B(n_1359),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1412),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1393),
.B(n_1347),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_SL g1501 ( 
.A(n_1410),
.B(n_1366),
.C(n_1342),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1412),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1382),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1404),
.B(n_1414),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1445),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1396),
.A2(n_1308),
.B1(n_1348),
.B2(n_1334),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1417),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1403),
.B(n_1346),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1504),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1476),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1452),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1456),
.A2(n_1444),
.B1(n_1409),
.B2(n_1382),
.C(n_1442),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1453),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1463),
.B(n_1388),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1457),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1498),
.B(n_1420),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1460),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_1388),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1390),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1462),
.A2(n_1442),
.B1(n_1373),
.B2(n_1394),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1461),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1476),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1390),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1501),
.A2(n_1394),
.B1(n_1425),
.B2(n_1422),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1433),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1448),
.B(n_1433),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1455),
.B(n_1459),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1473),
.B(n_1420),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1483),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1469),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1471),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1501),
.A2(n_1425),
.B1(n_1405),
.B2(n_1421),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1403),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1467),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1475),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1466),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1447),
.B(n_1404),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1485),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1492),
.B(n_1438),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1449),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1485),
.B(n_1443),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1465),
.B(n_1416),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1479),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1480),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1486),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1474),
.B(n_1443),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1467),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1467),
.B(n_1401),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1464),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1494),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1495),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1450),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1499),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1490),
.Y(n_1559)
);

NAND4xp25_ASAP7_75t_L g1560 ( 
.A(n_1472),
.B(n_1382),
.C(n_1409),
.D(n_1416),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1503),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1503),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1481),
.B(n_1401),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1491),
.B(n_1405),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1482),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1464),
.B(n_1409),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1505),
.B(n_1439),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1502),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1507),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1451),
.B(n_1421),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1490),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1559),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1510),
.B(n_1451),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1477),
.Y(n_1574)
);

NAND2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1415),
.Y(n_1575)
);

OAI211xp5_ASAP7_75t_L g1576 ( 
.A1(n_1560),
.A2(n_1472),
.B(n_1496),
.C(n_1506),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1512),
.A2(n_1496),
.B1(n_1484),
.B2(n_1497),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1550),
.B(n_1458),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1458),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1531),
.B(n_1468),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1516),
.B(n_1422),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1513),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1551),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1540),
.B(n_1424),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1513),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1542),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1551),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_SL g1589 ( 
.A(n_1510),
.B(n_1439),
.Y(n_1589)
);

CKINVDCx16_ASAP7_75t_R g1590 ( 
.A(n_1553),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1522),
.B(n_1487),
.C(n_1470),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_SL g1592 ( 
.A(n_1526),
.B(n_1487),
.C(n_1470),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1424),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1516),
.B(n_1417),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1524),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1536),
.B(n_1414),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1548),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1557),
.B(n_1415),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1521),
.B(n_1525),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1521),
.B(n_1418),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1518),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1565),
.B(n_1415),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1514),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1525),
.B(n_1418),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1528),
.B(n_1426),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1524),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_1468),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1544),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1528),
.B(n_1527),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1563),
.B(n_1426),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1539),
.B(n_1441),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1514),
.B(n_1441),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1563),
.B(n_1436),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1529),
.B(n_1430),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1436),
.C(n_1430),
.D(n_1346),
.Y(n_1617)
);

OA211x2_ASAP7_75t_L g1618 ( 
.A1(n_1578),
.A2(n_1535),
.B(n_1534),
.C(n_1543),
.Y(n_1618)
);

AOI221x1_ASAP7_75t_L g1619 ( 
.A1(n_1599),
.A2(n_1566),
.B1(n_1571),
.B2(n_1562),
.C(n_1561),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1576),
.A2(n_1509),
.B(n_1571),
.C(n_1568),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1583),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1509),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1591),
.A2(n_1564),
.B(n_1538),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1600),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1575),
.A2(n_1518),
.B1(n_1538),
.B2(n_1530),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1602),
.A2(n_1541),
.B(n_1530),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1575),
.Y(n_1628)
);

O2A1O1Ixp5_ASAP7_75t_SL g1629 ( 
.A1(n_1599),
.A2(n_1545),
.B(n_1515),
.C(n_1517),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1630)
);

AND4x1_ASAP7_75t_L g1631 ( 
.A(n_1596),
.B(n_1564),
.C(n_1547),
.D(n_1537),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1598),
.B(n_1603),
.C(n_1577),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1600),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1610),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1592),
.A2(n_1569),
.B1(n_1511),
.B2(n_1549),
.C(n_1555),
.Y(n_1635)
);

NAND3x2_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1541),
.C(n_1566),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1610),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1575),
.A2(n_1373),
.B1(n_1515),
.B2(n_1517),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1587),
.A2(n_1519),
.B(n_1533),
.C(n_1532),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1572),
.A2(n_1544),
.B(n_1519),
.C(n_1523),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1594),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1594),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1613),
.A2(n_1308),
.B1(n_1567),
.B2(n_1561),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1581),
.A2(n_1562),
.B1(n_1567),
.B2(n_1558),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1567),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1597),
.B(n_1523),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1601),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1593),
.A2(n_1558),
.B(n_1556),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1574),
.A2(n_1556),
.B(n_1546),
.C(n_1545),
.Y(n_1649)
);

AOI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1588),
.A2(n_1533),
.B(n_1532),
.C(n_1546),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1584),
.B(n_1375),
.Y(n_1651)
);

OAI21xp33_ASAP7_75t_L g1652 ( 
.A1(n_1585),
.A2(n_1376),
.B(n_1359),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1372),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1579),
.B(n_1376),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1270),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1621),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1645),
.B(n_1573),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1622),
.B(n_1572),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1623),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1629),
.B(n_1573),
.C(n_1580),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1573),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1633),
.B(n_1589),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1606),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1637),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1630),
.B(n_1582),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1619),
.B(n_1609),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1626),
.B(n_1606),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1641),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1642),
.B(n_1647),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1624),
.B(n_1601),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1595),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1656),
.B(n_1605),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1582),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1646),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1639),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1651),
.B(n_1605),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1639),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1640),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1655),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1654),
.B(n_1589),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1632),
.B(n_1607),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1648),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1650),
.B(n_1607),
.Y(n_1688)
);

NAND2x1_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1586),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1635),
.B(n_1586),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1662),
.B(n_1620),
.C(n_1635),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1663),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1604),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1659),
.B(n_1612),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1604),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1580),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1674),
.B(n_1608),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1676),
.B(n_1615),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1673),
.B(n_1614),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1614),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1668),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_L g1704 ( 
.A(n_1660),
.B(n_1620),
.C(n_1649),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1617),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1690),
.B(n_1649),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1638),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1680),
.B(n_1618),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1669),
.B(n_1368),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1677),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1685),
.B(n_1665),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1680),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1664),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1677),
.Y(n_1716)
);

OAI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1686),
.A2(n_1687),
.B(n_1682),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1684),
.B(n_1196),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_SL g1719 ( 
.A(n_1703),
.B(n_1678),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1705),
.B(n_1658),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1691),
.A2(n_1679),
.B1(n_1681),
.B2(n_1688),
.C(n_1689),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1701),
.B(n_1675),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1703),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1701),
.A2(n_1661),
.B(n_1672),
.C(n_1657),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1692),
.B(n_1661),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1693),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1707),
.A2(n_1683),
.B(n_1666),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1671),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1694),
.B(n_1683),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1704),
.A2(n_1261),
.B(n_1179),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1693),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1200),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1695),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1714),
.B(n_1368),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1710),
.B(n_1368),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1699),
.Y(n_1736)
);

OAI211xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1712),
.A2(n_1292),
.B(n_1324),
.C(n_1331),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1717),
.C(n_1716),
.Y(n_1738)
);

OAI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1722),
.A2(n_1708),
.B1(n_1709),
.B2(n_1696),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1721),
.A2(n_1708),
.B1(n_1709),
.B2(n_1706),
.C(n_1715),
.Y(n_1740)
);

AND4x1_ASAP7_75t_L g1741 ( 
.A(n_1738),
.B(n_1702),
.C(n_1711),
.D(n_1713),
.Y(n_1741)
);

AOI211xp5_ASAP7_75t_L g1742 ( 
.A1(n_1723),
.A2(n_1718),
.B(n_1331),
.C(n_1324),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1727),
.A2(n_1292),
.B1(n_1357),
.B2(n_1349),
.C(n_1369),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1728),
.B(n_1217),
.C(n_1196),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1729),
.A2(n_1275),
.B(n_1217),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1719),
.B(n_1229),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1736),
.A2(n_1224),
.B1(n_1249),
.B2(n_1369),
.Y(n_1747)
);

OAI21xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1726),
.A2(n_1357),
.B(n_1349),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1724),
.A2(n_1229),
.B1(n_1200),
.B2(n_1234),
.C(n_1125),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1725),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1720),
.A2(n_1278),
.B(n_1275),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1730),
.A2(n_1153),
.B1(n_1159),
.B2(n_1127),
.C(n_1122),
.Y(n_1752)
);

NAND4xp25_ASAP7_75t_L g1753 ( 
.A(n_1733),
.B(n_1159),
.C(n_1098),
.D(n_1137),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1732),
.A2(n_1730),
.B1(n_1731),
.B2(n_1735),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1234),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1740),
.A2(n_1737),
.B1(n_1118),
.B2(n_1115),
.Y(n_1756)
);

AOI21xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1739),
.A2(n_1234),
.B(n_1115),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1752),
.A2(n_1118),
.B1(n_1136),
.B2(n_1137),
.C(n_1098),
.Y(n_1758)
);

O2A1O1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1746),
.A2(n_1083),
.B(n_1085),
.C(n_1123),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1754),
.A2(n_1136),
.B(n_1085),
.C(n_1083),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1741),
.B(n_1189),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1750),
.A2(n_1083),
.B1(n_1085),
.B2(n_1123),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1742),
.A2(n_1083),
.B(n_1085),
.C(n_1123),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1745),
.A2(n_1278),
.B(n_1123),
.C(n_1255),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1751),
.A2(n_1189),
.B(n_1184),
.C(n_1131),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1753),
.A2(n_1189),
.B(n_1184),
.C(n_1131),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1744),
.A2(n_1194),
.B(n_1172),
.C(n_1110),
.Y(n_1767)
);

OAI211xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1749),
.A2(n_1164),
.B(n_1160),
.C(n_1162),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1748),
.A2(n_1139),
.B(n_1172),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1761),
.A2(n_1743),
.B1(n_1747),
.B2(n_1755),
.C(n_1167),
.Y(n_1770)
);

NAND4xp75_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1172),
.C(n_1128),
.D(n_1110),
.Y(n_1771)
);

NOR2x1_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1189),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1279),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1768),
.B(n_1249),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1757),
.A2(n_1164),
.B1(n_1160),
.B2(n_1162),
.C(n_1165),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1255),
.C(n_1140),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1765),
.B(n_1279),
.Y(n_1777)
);

NOR3xp33_ASAP7_75t_L g1778 ( 
.A(n_1759),
.B(n_1140),
.C(n_1128),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1764),
.B(n_1167),
.C(n_1139),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1762),
.A2(n_1167),
.B(n_1139),
.C(n_1120),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_L g1781 ( 
.A(n_1770),
.B(n_1767),
.C(n_1766),
.Y(n_1781)
);

NAND4xp75_ASAP7_75t_L g1782 ( 
.A(n_1772),
.B(n_1769),
.C(n_1120),
.D(n_1239),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1773),
.A2(n_1120),
.B(n_1214),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_L g1784 ( 
.A(n_1776),
.B(n_1184),
.C(n_1214),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1774),
.A2(n_1165),
.B1(n_1184),
.B2(n_1174),
.C(n_1090),
.Y(n_1785)
);

NAND2xp33_ASAP7_75t_L g1786 ( 
.A(n_1781),
.B(n_1771),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1784),
.B(n_1778),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1782),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1785),
.Y(n_1789)
);

AOI222xp33_ASAP7_75t_L g1790 ( 
.A1(n_1783),
.A2(n_1775),
.B1(n_1777),
.B2(n_1779),
.C1(n_1780),
.C2(n_1249),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1783),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1788),
.B(n_1239),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1787),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1786),
.Y(n_1794)
);

AO22x2_ASAP7_75t_L g1795 ( 
.A1(n_1791),
.A2(n_1090),
.B1(n_1111),
.B2(n_1107),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1792),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1793),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_L g1798 ( 
.A(n_1794),
.B(n_1789),
.C(n_1790),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1795),
.B(n_1279),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1796),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1797),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1798),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1799),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1797),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1800),
.B(n_1279),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1802),
.A2(n_1249),
.B1(n_1111),
.B2(n_1107),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1801),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1807),
.B(n_1804),
.Y(n_1808)
);

OR2x6_ASAP7_75t_L g1809 ( 
.A(n_1808),
.B(n_1803),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1805),
.B1(n_1806),
.B2(n_1249),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1239),
.B1(n_1246),
.B2(n_1174),
.Y(n_1811)
);

AO21x2_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1202),
.B(n_1113),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1812),
.A2(n_1202),
.B(n_1246),
.Y(n_1813)
);

AOI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1116),
.B(n_1121),
.C(n_1113),
.Y(n_1814)
);


endmodule