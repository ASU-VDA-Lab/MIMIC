module real_aes_8737_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_1), .A2(n_151), .B(n_154), .C(n_157), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_2), .A2(n_177), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g537 ( .A(n_3), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_4), .B(n_200), .Y(n_223) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_5), .A2(n_177), .B(n_465), .Y(n_464) );
AND2x6_ASAP7_75t_L g151 ( .A(n_6), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g184 ( .A(n_7), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_41), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_41), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_9), .A2(n_231), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_10), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g469 ( .A(n_11), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_12), .B(n_206), .Y(n_508) );
INVx1_ASAP7_75t_L g143 ( .A(n_13), .Y(n_143) );
INVx1_ASAP7_75t_L g520 ( .A(n_14), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_15), .A2(n_185), .B(n_195), .C(n_198), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_16), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_17), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_18), .B(n_476), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_19), .B(n_177), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_20), .B(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_21), .A2(n_206), .B(n_207), .C(n_209), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_22), .B(n_200), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_23), .B(n_163), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_24), .A2(n_197), .B(n_198), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_25), .B(n_163), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_26), .Y(n_259) );
INVx1_ASAP7_75t_L g249 ( .A(n_27), .Y(n_249) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_28), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_29), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_30), .B(n_163), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_31), .A2(n_65), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_31), .Y(n_128) );
INVx1_ASAP7_75t_L g236 ( .A(n_32), .Y(n_236) );
INVx1_ASAP7_75t_L g458 ( .A(n_33), .Y(n_458) );
INVx2_ASAP7_75t_L g149 ( .A(n_34), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_35), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_36), .A2(n_206), .B(n_219), .C(n_221), .Y(n_218) );
INVxp67_ASAP7_75t_L g238 ( .A(n_37), .Y(n_238) );
CKINVDCx14_ASAP7_75t_R g217 ( .A(n_38), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_39), .A2(n_154), .B(n_248), .C(n_252), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_40), .A2(n_151), .B(n_154), .C(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g457 ( .A(n_42), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_43), .A2(n_165), .B(n_182), .C(n_183), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_44), .B(n_163), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_45), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_46), .Y(n_233) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_47), .A2(n_446), .B1(n_721), .B2(n_724), .C1(n_725), .C2(n_727), .Y(n_445) );
INVx1_ASAP7_75t_L g204 ( .A(n_48), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_49), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_50), .B(n_177), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_51), .A2(n_154), .B1(n_209), .B2(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_52), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_53), .Y(n_534) );
CKINVDCx14_ASAP7_75t_R g179 ( .A(n_54), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_55), .A2(n_182), .B(n_221), .C(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_56), .Y(n_500) );
INVx1_ASAP7_75t_L g466 ( .A(n_57), .Y(n_466) );
INVx1_ASAP7_75t_L g152 ( .A(n_58), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_59), .A2(n_78), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_59), .Y(n_723) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
INVx1_ASAP7_75t_SL g220 ( .A(n_61), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_62), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_63), .B(n_200), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_64), .A2(n_102), .B1(n_111), .B2(n_731), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_65), .Y(n_127) );
INVx1_ASAP7_75t_L g262 ( .A(n_66), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_SL g475 ( .A1(n_67), .A2(n_221), .B(n_476), .C(n_477), .Y(n_475) );
INVxp67_ASAP7_75t_L g478 ( .A(n_68), .Y(n_478) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_70), .A2(n_177), .B(n_178), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_71), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_72), .A2(n_177), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_73), .Y(n_461) );
INVx1_ASAP7_75t_L g494 ( .A(n_74), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_75), .A2(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g193 ( .A(n_76), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_77), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_78), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_79), .A2(n_151), .B(n_154), .C(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_80), .A2(n_177), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g196 ( .A(n_81), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_82), .B(n_237), .Y(n_488) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
INVx1_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_85), .B(n_476), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_86), .A2(n_151), .B(n_154), .C(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g119 ( .A(n_87), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g720 ( .A(n_87), .B(n_121), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_88), .A2(n_154), .B(n_261), .C(n_264), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_89), .B(n_139), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_90), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_91), .A2(n_151), .B(n_154), .C(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_92), .Y(n_512) );
INVx1_ASAP7_75t_L g474 ( .A(n_93), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_94), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_95), .B(n_237), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_96), .B(n_170), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_97), .B(n_170), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g208 ( .A(n_99), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_100), .A2(n_177), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g731 ( .A(n_104), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g717 ( .A(n_107), .B(n_121), .Y(n_717) );
NOR2x2_ASAP7_75t_L g729 ( .A(n_107), .B(n_120), .Y(n_729) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_444), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g730 ( .A(n_116), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_441), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_119), .Y(n_443) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_129), .A2(n_447), .B1(n_715), .B2(n_718), .Y(n_446) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_130), .A2(n_715), .B1(n_720), .B2(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_396), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_308), .C(n_346), .D(n_367), .E(n_384), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_280), .C(n_301), .Y(n_132) );
OAI221xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_212), .B1(n_243), .B2(n_267), .C(n_271), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_172), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_136), .B(n_269), .Y(n_288) );
OR2x2_ASAP7_75t_L g315 ( .A(n_136), .B(n_189), .Y(n_315) );
AND2x2_ASAP7_75t_L g329 ( .A(n_136), .B(n_189), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_136), .B(n_175), .Y(n_343) );
AND2x2_ASAP7_75t_L g381 ( .A(n_136), .B(n_345), .Y(n_381) );
AND2x2_ASAP7_75t_L g410 ( .A(n_136), .B(n_320), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_136), .B(n_292), .Y(n_427) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g307 ( .A(n_137), .B(n_188), .Y(n_307) );
BUFx3_ASAP7_75t_L g332 ( .A(n_137), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_137), .B(n_189), .Y(n_361) );
AND3x2_ASAP7_75t_L g374 ( .A(n_137), .B(n_375), .C(n_376), .Y(n_374) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_167), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_138), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_138), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_138), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_139), .A2(n_176), .B(n_187), .Y(n_175) );
INVx2_ASAP7_75t_L g242 ( .A(n_139), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_139), .A2(n_146), .B(n_246), .C(n_247), .Y(n_245) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_139), .A2(n_515), .B(n_521), .Y(n_514) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g171 ( .A(n_140), .B(n_141), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_153), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_146), .A2(n_259), .B(n_260), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_146), .A2(n_186), .B1(n_455), .B2(n_459), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_146), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_146), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AND2x4_ASAP7_75t_L g177 ( .A(n_147), .B(n_151), .Y(n_177) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
INVx3_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
INVx1_ASAP7_75t_L g476 ( .A(n_150), .Y(n_476) );
INVx4_ASAP7_75t_SL g186 ( .A(n_151), .Y(n_186) );
BUFx3_ASAP7_75t_L g252 ( .A(n_151), .Y(n_252) );
INVx5_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
O2A1O1Ixp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_162), .C(n_164), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_159), .A2(n_164), .B(n_262), .C(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_160), .A2(n_161), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
INVx2_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
INVx4_ASAP7_75t_L g206 ( .A(n_163), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_164), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_164), .A2(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx3_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_169), .B(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_169), .A2(n_258), .B(n_265), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g490 ( .A(n_169), .B(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_170), .Y(n_190) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_170), .A2(n_472), .B(n_479), .Y(n_471) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
INVx1_ASAP7_75t_L g297 ( .A(n_172), .Y(n_297) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_188), .Y(n_172) );
AOI32xp33_ASAP7_75t_L g352 ( .A1(n_173), .A2(n_304), .A3(n_353), .B1(n_356), .B2(n_357), .Y(n_352) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g279 ( .A(n_174), .B(n_188), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_174), .B(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_174), .B(n_329), .Y(n_357) );
OR2x2_ASAP7_75t_L g363 ( .A(n_174), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_174), .B(n_318), .Y(n_388) );
OR2x2_ASAP7_75t_L g406 ( .A(n_174), .B(n_225), .Y(n_406) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g270 ( .A(n_175), .B(n_201), .Y(n_270) );
INVx2_ASAP7_75t_L g292 ( .A(n_175), .Y(n_292) );
OR2x2_ASAP7_75t_L g314 ( .A(n_175), .B(n_201), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_175), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_175), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_175), .B(n_269), .Y(n_375) );
BUFx2_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B(n_181), .C(n_186), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_180), .A2(n_186), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_180), .A2(n_186), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_180), .A2(n_186), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_180), .A2(n_186), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_180), .A2(n_186), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_180), .A2(n_186), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_180), .A2(n_186), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
INVx5_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_185), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_185), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
INVx1_ASAP7_75t_SL g426 ( .A(n_188), .Y(n_426) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_201), .Y(n_188) );
INVx1_ASAP7_75t_SL g269 ( .A(n_189), .Y(n_269) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_189), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_189), .B(n_355), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_189), .B(n_292), .C(n_410), .Y(n_421) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_199), .Y(n_189) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_190), .A2(n_202), .B(n_211), .Y(n_201) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_190), .A2(n_215), .B(n_223), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_197), .B(n_208), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_197), .B(n_520), .Y(n_519) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_200), .A2(n_464), .B(n_470), .Y(n_463) );
INVx2_ASAP7_75t_L g320 ( .A(n_201), .Y(n_320) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_201), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_206), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g539 ( .A(n_209), .Y(n_539) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_224), .Y(n_212) );
INVx1_ASAP7_75t_L g356 ( .A(n_213), .Y(n_356) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_256), .Y(n_274) );
INVx2_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
AND2x2_ASAP7_75t_L g296 ( .A(n_214), .B(n_257), .Y(n_296) );
AND2x2_ASAP7_75t_L g311 ( .A(n_214), .B(n_244), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_214), .B(n_295), .Y(n_323) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_222), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_224), .B(n_339), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_224), .B(n_296), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_224), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_224), .B(n_290), .Y(n_418) );
BUFx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g255 ( .A(n_225), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_225), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g300 ( .A(n_225), .B(n_244), .Y(n_300) );
AND2x2_ASAP7_75t_L g326 ( .A(n_225), .B(n_256), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_225), .B(n_366), .Y(n_365) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_230), .B(n_240), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_227), .A2(n_285), .B(n_286), .Y(n_284) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_227), .A2(n_493), .B(n_499), .Y(n_492) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_SL g484 ( .A1(n_228), .A2(n_485), .B(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_229), .A2(n_454), .B(n_460), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_229), .B(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_229), .A2(n_533), .B(n_540), .Y(n_532) );
INVx1_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_235), .B(n_239), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_237), .A2(n_249), .B(n_250), .C(n_251), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_237), .A2(n_537), .B(n_538), .C(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g251 ( .A(n_239), .Y(n_251) );
INVx1_ASAP7_75t_L g286 ( .A(n_240), .Y(n_286) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_242), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_242), .A2(n_504), .B(n_511), .Y(n_503) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_255), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_244), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g290 ( .A(n_244), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_SL g295 ( .A(n_244), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_244), .B(n_282), .Y(n_348) );
OR2x2_ASAP7_75t_L g358 ( .A(n_244), .B(n_284), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_244), .B(n_326), .Y(n_386) );
OR2x2_ASAP7_75t_L g416 ( .A(n_244), .B(n_256), .Y(n_416) );
AND2x2_ASAP7_75t_L g420 ( .A(n_244), .B(n_257), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_244), .B(n_296), .Y(n_433) );
AND2x2_ASAP7_75t_L g440 ( .A(n_244), .B(n_322), .Y(n_440) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_253), .Y(n_244) );
INVx1_ASAP7_75t_SL g383 ( .A(n_255), .Y(n_383) );
AND2x2_ASAP7_75t_L g322 ( .A(n_256), .B(n_284), .Y(n_322) );
AND2x2_ASAP7_75t_L g336 ( .A(n_256), .B(n_291), .Y(n_336) );
AND2x2_ASAP7_75t_L g339 ( .A(n_256), .B(n_295), .Y(n_339) );
INVx1_ASAP7_75t_L g366 ( .A(n_256), .Y(n_366) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_268), .A2(n_314), .B(n_438), .C(n_439), .Y(n_437) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g344 ( .A(n_269), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_270), .B(n_287), .Y(n_302) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_329), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_275), .B(n_279), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_273), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g299 ( .A(n_274), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_274), .B(n_295), .Y(n_340) );
AND2x2_ASAP7_75t_L g431 ( .A(n_274), .B(n_282), .Y(n_431) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_291), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_289), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_288), .A3(n_289), .B1(n_292), .B2(n_293), .C1(n_297), .C2(n_298), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_287), .Y(n_281) );
AND2x2_ASAP7_75t_L g392 ( .A(n_282), .B(n_304), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_282), .B(n_356), .Y(n_438) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g401 ( .A(n_288), .B(n_314), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_289), .B(n_383), .Y(n_382) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_290), .B(n_322), .Y(n_379) );
AND2x2_ASAP7_75t_L g325 ( .A(n_291), .B(n_295), .Y(n_325) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_334), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_292), .A2(n_371), .B(n_431), .C(n_432), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_293), .A2(n_306), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_295), .B(n_322), .Y(n_362) );
AND2x2_ASAP7_75t_L g368 ( .A(n_295), .B(n_336), .Y(n_368) );
AND2x2_ASAP7_75t_L g402 ( .A(n_295), .B(n_304), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_296), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g412 ( .A(n_296), .Y(n_412) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_328), .B1(n_330), .B2(n_335), .Y(n_327) );
OAI22xp5_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_303), .B1(n_305), .B2(n_306), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_338), .B1(n_340), .B2(n_341), .Y(n_337) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_307), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_417), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_312), .B(n_316), .C(n_337), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OR2x2_ASAP7_75t_L g378 ( .A(n_314), .B(n_331), .Y(n_378) );
INVx1_ASAP7_75t_L g429 ( .A(n_314), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_315), .A2(n_317), .B1(n_321), .B2(n_324), .C(n_327), .Y(n_316) );
INVx2_ASAP7_75t_SL g371 ( .A(n_315), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g436 ( .A(n_318), .Y(n_436) );
AND2x2_ASAP7_75t_L g360 ( .A(n_319), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g407 ( .A(n_323), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_331), .B(n_433), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_335), .A2(n_347), .B(n_349), .C(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g424 ( .A(n_338), .Y(n_424) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_342), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g355 ( .A(n_345), .Y(n_355) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI222xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_358), .B1(n_359), .B2(n_362), .C1(n_363), .C2(n_365), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g391 ( .A(n_355), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_358), .B(n_412), .Y(n_411) );
NAND2xp33_ASAP7_75t_SL g389 ( .A(n_359), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g364 ( .A(n_361), .Y(n_364) );
AND2x2_ASAP7_75t_L g428 ( .A(n_361), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g394 ( .A(n_364), .B(n_391), .Y(n_394) );
INVx1_ASAP7_75t_L g423 ( .A(n_365), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_372), .C(n_377), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_371), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g422 ( .A1(n_374), .A2(n_402), .A3(n_407), .B1(n_423), .B2(n_424), .C1(n_425), .C2(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g409 ( .A(n_375), .B(n_410), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_380), .B2(n_382), .Y(n_377) );
INVxp33_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_389), .B2(n_392), .C(n_393), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NAND5xp2_ASAP7_75t_L g396 ( .A(n_397), .B(n_408), .C(n_422), .D(n_430), .E(n_434), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_402), .B(n_403), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp33_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_435), .B(n_436), .C(n_437), .Y(n_434) );
AOI31xp33_ASAP7_75t_L g417 ( .A1(n_412), .A2(n_418), .A3(n_419), .B(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g435 ( .A(n_433), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_441), .B(n_445), .C(n_730), .Y(n_444) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g726 ( .A(n_447), .Y(n_726) );
AND3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_640), .C(n_689), .Y(n_447) );
NOR3xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_547), .C(n_585), .Y(n_448) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_480), .B1(n_522), .B2(n_528), .C1(n_542), .C2(n_545), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_462), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_451), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_451), .B(n_590), .Y(n_681) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g558 ( .A(n_452), .B(n_471), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_452), .B(n_463), .Y(n_566) );
AND2x2_ASAP7_75t_L g601 ( .A(n_452), .B(n_578), .Y(n_601) );
OR2x2_ASAP7_75t_L g625 ( .A(n_452), .B(n_463), .Y(n_625) );
OR2x2_ASAP7_75t_L g633 ( .A(n_452), .B(n_532), .Y(n_633) );
AND2x2_ASAP7_75t_L g636 ( .A(n_452), .B(n_471), .Y(n_636) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g530 ( .A(n_453), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g544 ( .A(n_453), .B(n_471), .Y(n_544) );
AND2x2_ASAP7_75t_L g594 ( .A(n_453), .B(n_532), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_453), .B(n_463), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_453), .B(n_693), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_462), .A2(n_633), .B(n_634), .C(n_637), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_462), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_462), .B(n_577), .Y(n_699) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .Y(n_462) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_463), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g557 ( .A(n_463), .Y(n_557) );
AND2x2_ASAP7_75t_L g584 ( .A(n_463), .B(n_578), .Y(n_584) );
INVx1_ASAP7_75t_SL g592 ( .A(n_463), .Y(n_592) );
AND2x2_ASAP7_75t_L g615 ( .A(n_463), .B(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g693 ( .A(n_463), .Y(n_693) );
BUFx2_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
INVx1_ASAP7_75t_L g591 ( .A(n_471), .Y(n_591) );
INVx3_ASAP7_75t_L g616 ( .A(n_471), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_480), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_501), .Y(n_480) );
INVx1_ASAP7_75t_L g612 ( .A(n_481), .Y(n_612) );
OAI32xp33_ASAP7_75t_L g618 ( .A1(n_481), .A2(n_557), .A3(n_619), .B1(n_620), .B2(n_621), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_481), .A2(n_623), .B1(n_626), .B2(n_631), .Y(n_622) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g560 ( .A(n_482), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g638 ( .A(n_482), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g708 ( .A(n_482), .B(n_654), .Y(n_708) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
AND2x2_ASAP7_75t_L g523 ( .A(n_483), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g553 ( .A(n_483), .Y(n_553) );
INVx1_ASAP7_75t_L g572 ( .A(n_483), .Y(n_572) );
OR2x2_ASAP7_75t_L g580 ( .A(n_483), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g587 ( .A(n_483), .B(n_561), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_483), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g608 ( .A(n_483), .B(n_526), .Y(n_608) );
INVx3_ASAP7_75t_L g630 ( .A(n_483), .Y(n_630) );
AND2x2_ASAP7_75t_L g655 ( .A(n_483), .B(n_527), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_483), .B(n_620), .Y(n_703) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_490), .Y(n_483) );
INVx2_ASAP7_75t_L g527 ( .A(n_492), .Y(n_527) );
AND2x2_ASAP7_75t_L g659 ( .A(n_492), .B(n_502), .Y(n_659) );
INVx2_ASAP7_75t_L g701 ( .A(n_501), .Y(n_701) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
INVx1_ASAP7_75t_L g546 ( .A(n_502), .Y(n_546) );
AND2x2_ASAP7_75t_L g573 ( .A(n_502), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_502), .B(n_527), .Y(n_581) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_562), .Y(n_639) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g525 ( .A(n_503), .Y(n_525) );
AND2x2_ASAP7_75t_L g552 ( .A(n_503), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_503), .B(n_527), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_513), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_513), .B(n_527), .Y(n_620) );
AND2x2_ASAP7_75t_L g629 ( .A(n_513), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g654 ( .A(n_513), .Y(n_654) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g526 ( .A(n_514), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g562 ( .A(n_514), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_522), .A2(n_532), .B1(n_691), .B2(n_694), .Y(n_690) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g713 ( .A1(n_524), .A2(n_635), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_525), .B(n_630), .Y(n_647) );
INVx1_ASAP7_75t_L g672 ( .A(n_525), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_526), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_552), .Y(n_599) );
INVx2_ASAP7_75t_L g555 ( .A(n_527), .Y(n_555) );
INVx1_ASAP7_75t_L g605 ( .A(n_527), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_528), .A2(n_680), .B1(n_697), .B2(n_700), .C(n_702), .Y(n_696) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_529), .B(n_578), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_530), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g621 ( .A(n_530), .B(n_567), .Y(n_621) );
INVx3_ASAP7_75t_SL g662 ( .A(n_530), .Y(n_662) );
AND2x2_ASAP7_75t_L g606 ( .A(n_531), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g635 ( .A(n_531), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_531), .B(n_544), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_531), .B(n_590), .Y(n_676) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_532), .A2(n_604), .A3(n_626), .B1(n_674), .B2(n_676), .C1(n_677), .C2(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_543), .A2(n_546), .B(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_SL g623 ( .A(n_544), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g645 ( .A(n_544), .B(n_557), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_544), .B(n_584), .Y(n_660) );
INVxp67_ASAP7_75t_L g611 ( .A(n_546), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_546), .A2(n_618), .B(n_622), .C(n_632), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_556), .B1(n_559), .B2(n_563), .C(n_568), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g571 ( .A(n_555), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g688 ( .A(n_555), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_556), .A2(n_705), .B1(n_710), .B2(n_711), .C(n_713), .Y(n_704) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_557), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g604 ( .A(n_557), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_557), .B(n_635), .Y(n_642) );
AND2x2_ASAP7_75t_L g684 ( .A(n_557), .B(n_662), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_558), .B(n_583), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_558), .A2(n_570), .B1(n_680), .B2(n_681), .Y(n_679) );
OR2x2_ASAP7_75t_L g710 ( .A(n_558), .B(n_578), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g687 ( .A(n_561), .Y(n_687) );
AND2x2_ASAP7_75t_L g712 ( .A(n_561), .B(n_655), .Y(n_712) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g576 ( .A(n_566), .B(n_577), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_575), .B1(n_579), .B2(n_582), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g643 ( .A(n_571), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_571), .B(n_611), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g602 ( .A1(n_573), .A2(n_603), .A3(n_605), .B1(n_606), .B2(n_608), .C1(n_609), .C2(n_613), .Y(n_602) );
INVxp67_ASAP7_75t_L g596 ( .A(n_574), .Y(n_596) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_576), .A2(n_581), .B1(n_598), .B2(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_577), .B(n_590), .Y(n_677) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_578), .B(n_616), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_578), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g674 ( .A(n_580), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NAND3xp33_ASAP7_75t_SL g585 ( .A(n_586), .B(n_602), .C(n_617), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_593), .B2(n_595), .C(n_597), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_589), .B(n_594), .Y(n_593) );
INVx3_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g603 ( .A(n_594), .B(n_604), .Y(n_603) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_596), .Y(n_675) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_601), .B(n_615), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_604), .B(n_662), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_605), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g680 ( .A(n_608), .Y(n_680) );
AND2x2_ASAP7_75t_L g695 ( .A(n_608), .B(n_672), .Y(n_695) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_619), .A2(n_690), .B(n_696), .C(n_704), .Y(n_689) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g658 ( .A(n_629), .B(n_659), .Y(n_658) );
NAND2x1_ASAP7_75t_SL g700 ( .A(n_630), .B(n_701), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g670 ( .A(n_633), .Y(n_670) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g665 ( .A(n_639), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_639), .B(n_655), .Y(n_669) );
NOR5xp2_ASAP7_75t_L g640 ( .A(n_641), .B(n_656), .C(n_673), .D(n_679), .E(n_682), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_641) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_645), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g671 ( .A(n_655), .B(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_660), .B1(n_661), .B2(n_663), .C(n_666), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g709 ( .A(n_669), .Y(n_709) );
AOI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_687), .C(n_688), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx14_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx14_ASAP7_75t_R g724 ( .A(n_721), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx3_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
endmodule