module fake_jpeg_3442_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_51),
.B1(n_41),
.B2(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_66),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_40),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_42),
.C(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_51),
.B1(n_41),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_45),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_44),
.B1(n_39),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_44),
.B1(n_50),
.B2(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_8),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_6),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_0),
.B(n_2),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_100),
.B(n_7),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_98),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_3),
.B(n_4),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_73),
.C(n_16),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_112),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_109),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_17),
.B(n_34),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_100),
.B(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_73),
.B1(n_15),
.B2(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_6),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_121),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_112),
.C(n_101),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.C(n_26),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_96),
.C(n_93),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_129),
.B(n_24),
.Y(n_134)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_105),
.B1(n_99),
.B2(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_131),
.B1(n_125),
.B2(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_27),
.B(n_30),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_117),
.B1(n_124),
.B2(n_12),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_133),
.B(n_122),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_120),
.B(n_136),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_138),
.B(n_117),
.Y(n_148)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_22),
.A3(n_29),
.B1(n_28),
.B2(n_33),
.C1(n_13),
.C2(n_12),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_11),
.Y(n_150)
);


endmodule