module real_aes_7185_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_0), .A2(n_177), .B(n_178), .C(n_182), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_1), .B(n_171), .Y(n_184) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_92), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_3), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_165), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_5), .A2(n_145), .B(n_162), .C(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_6), .A2(n_165), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_7), .B(n_171), .Y(n_483) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_8), .A2(n_137), .B(n_259), .Y(n_258) );
AND2x6_ASAP7_75t_L g162 ( .A(n_9), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_10), .A2(n_145), .B(n_162), .C(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g574 ( .A(n_11), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_12), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_12), .B(n_40), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_13), .B(n_181), .Y(n_523) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_15), .A2(n_104), .B1(n_112), .B2(n_729), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_16), .B(n_156), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_17), .A2(n_157), .B(n_532), .C(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_18), .B(n_171), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_19), .B(n_199), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_20), .A2(n_145), .B(n_191), .C(n_198), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_180), .B(n_233), .C(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_22), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_23), .B(n_181), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_24), .B(n_181), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_25), .Y(n_501) );
INVx1_ASAP7_75t_L g471 ( .A(n_26), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_27), .A2(n_145), .B(n_198), .C(n_262), .Y(n_261) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_29), .Y(n_519) );
INVx1_ASAP7_75t_L g495 ( .A(n_30), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_31), .A2(n_165), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g147 ( .A(n_32), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_33), .A2(n_160), .B(n_214), .C(n_215), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_34), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_35), .A2(n_180), .B(n_480), .C(n_482), .Y(n_479) );
INVxp67_ASAP7_75t_L g496 ( .A(n_36), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_37), .B(n_264), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_38), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_39), .A2(n_145), .B(n_198), .C(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_41), .A2(n_182), .B(n_572), .C(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_42), .B(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_43), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_44), .B(n_156), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_45), .B(n_165), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_46), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_47), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_48), .A2(n_160), .B(n_214), .C(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g179 ( .A(n_49), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_50), .A2(n_126), .B1(n_440), .B2(n_441), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_50), .Y(n_440) );
INVx1_ASAP7_75t_L g243 ( .A(n_51), .Y(n_243) );
INVx1_ASAP7_75t_L g539 ( .A(n_52), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_53), .B(n_165), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_54), .A2(n_72), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_54), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_55), .Y(n_203) );
AOI222xp33_ASAP7_75t_SL g446 ( .A1(n_56), .A2(n_447), .B1(n_453), .B2(n_723), .C1(n_724), .C2(n_725), .Y(n_446) );
CKINVDCx14_ASAP7_75t_R g570 ( .A(n_57), .Y(n_570) );
INVx1_ASAP7_75t_L g163 ( .A(n_58), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_59), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_60), .B(n_171), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_61), .A2(n_152), .B(n_197), .C(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_62), .A2(n_71), .B1(n_451), .B2(n_452), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_62), .Y(n_451) );
INVx1_ASAP7_75t_L g141 ( .A(n_63), .Y(n_141) );
INVx1_ASAP7_75t_SL g481 ( .A(n_64), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_66), .B(n_156), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_67), .B(n_171), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_68), .B(n_157), .Y(n_230) );
INVx1_ASAP7_75t_L g504 ( .A(n_69), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_70), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_71), .Y(n_452) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_73), .B(n_193), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_74), .A2(n_145), .B(n_150), .C(n_160), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_75), .Y(n_252) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_77), .A2(n_165), .B(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_78), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_79), .A2(n_165), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_80), .A2(n_189), .B(n_491), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_81), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_82), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_82), .Y(n_448) );
INVx1_ASAP7_75t_L g530 ( .A(n_83), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_84), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_85), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_86), .A2(n_165), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g533 ( .A(n_87), .Y(n_533) );
INVx2_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVx1_ASAP7_75t_L g522 ( .A(n_89), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_90), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_91), .B(n_181), .Y(n_231) );
OR2x2_ASAP7_75t_L g120 ( .A(n_92), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g457 ( .A(n_92), .B(n_122), .Y(n_457) );
INVx2_ASAP7_75t_L g722 ( .A(n_92), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_93), .A2(n_145), .B(n_160), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_94), .B(n_165), .Y(n_212) );
INVx1_ASAP7_75t_L g216 ( .A(n_95), .Y(n_216) );
INVxp67_ASAP7_75t_L g255 ( .A(n_96), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_97), .B(n_137), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_98), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g151 ( .A(n_99), .Y(n_151) );
INVx1_ASAP7_75t_L g226 ( .A(n_100), .Y(n_226) );
INVx2_ASAP7_75t_L g542 ( .A(n_101), .Y(n_542) );
AND2x2_ASAP7_75t_L g245 ( .A(n_102), .B(n_201), .Y(n_245) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g730 ( .A(n_105), .Y(n_730) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_445), .Y(n_112) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_114), .B(n_442), .C(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_125), .B(n_442), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_120), .Y(n_444) );
NOR2x2_ASAP7_75t_L g723 ( .A(n_121), .B(n_722), .Y(n_723) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g721 ( .A(n_122), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g441 ( .A(n_126), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_130), .Y(n_126) );
INVx1_ASAP7_75t_L g454 ( .A(n_130), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_130), .A2(n_459), .B1(n_726), .B2(n_727), .Y(n_725) );
OR3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_348), .C(n_397), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_282), .C(n_311), .D(n_319), .E(n_334), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_205), .B(n_221), .C(n_266), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_185), .Y(n_133) );
AND2x2_ASAP7_75t_L g277 ( .A(n_134), .B(n_274), .Y(n_277) );
AND2x2_ASAP7_75t_L g310 ( .A(n_134), .B(n_186), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_134), .B(n_209), .Y(n_403) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_170), .Y(n_134) );
INVx2_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
BUFx2_ASAP7_75t_L g377 ( .A(n_135), .Y(n_377) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_168), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_136), .B(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_136), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_136), .A2(n_225), .B(n_235), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_136), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_136), .A2(n_500), .B(n_507), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_136), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_137), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_137), .A2(n_260), .B(n_261), .Y(n_259) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g237 ( .A(n_138), .Y(n_237) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_139), .B(n_140), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_164), .Y(n_143) );
INVx5_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
BUFx3_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx1_ASAP7_75t_L g234 ( .A(n_147), .Y(n_234) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
AND2x2_ASAP7_75t_L g166 ( .A(n_149), .B(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
INVx1_ASAP7_75t_L g264 ( .A(n_149), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .C(n_158), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_153), .A2(n_156), .B1(n_495), .B2(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_153), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_153), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g193 ( .A(n_154), .Y(n_193) );
INVx2_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_156), .B(n_255), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_156), .A2(n_196), .B(n_471), .C(n_472), .Y(n_470) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_157), .B(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g482 ( .A(n_159), .Y(n_482) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_161), .A2(n_174), .B(n_175), .C(n_176), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_161), .A2(n_175), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_161), .A2(n_175), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_161), .A2(n_175), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_161), .A2(n_175), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g538 ( .A1(n_161), .A2(n_175), .B(n_539), .C(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_SL g569 ( .A1(n_161), .A2(n_175), .B(n_570), .C(n_571), .Y(n_569) );
INVx4_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g165 ( .A(n_162), .B(n_166), .Y(n_165) );
BUFx3_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_162), .B(n_166), .Y(n_227) );
BUFx2_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
INVx1_ASAP7_75t_L g197 ( .A(n_167), .Y(n_197) );
AND2x2_ASAP7_75t_L g185 ( .A(n_170), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g275 ( .A(n_170), .Y(n_275) );
AND2x2_ASAP7_75t_L g361 ( .A(n_170), .B(n_274), .Y(n_361) );
AND2x2_ASAP7_75t_L g416 ( .A(n_170), .B(n_208), .Y(n_416) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_184), .Y(n_170) );
INVx2_ASAP7_75t_L g214 ( .A(n_175), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_180), .B(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g572 ( .A(n_181), .Y(n_572) );
INVx2_ASAP7_75t_L g506 ( .A(n_182), .Y(n_506) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
INVx1_ASAP7_75t_L g534 ( .A(n_183), .Y(n_534) );
INVx1_ASAP7_75t_L g333 ( .A(n_185), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_185), .B(n_209), .Y(n_380) );
INVx5_ASAP7_75t_L g274 ( .A(n_186), .Y(n_274) );
AND2x4_ASAP7_75t_L g295 ( .A(n_186), .B(n_275), .Y(n_295) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_186), .Y(n_317) );
AND2x2_ASAP7_75t_L g392 ( .A(n_186), .B(n_377), .Y(n_392) );
AND2x2_ASAP7_75t_L g395 ( .A(n_186), .B(n_210), .Y(n_395) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_202), .Y(n_186) );
AOI21xp5_ASAP7_75t_SL g187 ( .A1(n_188), .A2(n_190), .B(n_199), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_196), .Y(n_191) );
INVx2_ASAP7_75t_L g195 ( .A(n_193), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_195), .A2(n_216), .B(n_217), .C(n_218), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_195), .A2(n_218), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_195), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_L g521 ( .A1(n_195), .A2(n_506), .B(n_522), .C(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_197), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_200), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g204 ( .A(n_201), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_201), .A2(n_240), .B(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_201), .A2(n_227), .B(n_468), .C(n_469), .Y(n_467) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_201), .A2(n_568), .B(n_575), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_204), .A2(n_518), .B(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_205), .B(n_275), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_205), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_209), .Y(n_206) );
AND2x2_ASAP7_75t_L g300 ( .A(n_207), .B(n_275), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_207), .B(n_210), .Y(n_318) );
INVx1_ASAP7_75t_L g338 ( .A(n_207), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_207), .B(n_274), .Y(n_383) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_207), .Y(n_425) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_208), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_209), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_209), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_209), .A2(n_270), .B(n_331), .C(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g337 ( .A(n_209), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g346 ( .A(n_209), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g350 ( .A(n_209), .B(n_274), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_209), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g365 ( .A(n_209), .B(n_275), .Y(n_365) );
AND2x2_ASAP7_75t_L g415 ( .A(n_209), .B(n_416), .Y(n_415) );
INVx5_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
AND2x2_ASAP7_75t_L g320 ( .A(n_210), .B(n_273), .Y(n_320) );
AND2x2_ASAP7_75t_L g332 ( .A(n_210), .B(n_307), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_210), .B(n_361), .Y(n_379) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_219), .Y(n_210) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_246), .Y(n_221) );
INVx1_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_238), .Y(n_222) );
OR2x2_ASAP7_75t_L g270 ( .A(n_223), .B(n_238), .Y(n_270) );
NAND3xp33_ASAP7_75t_L g276 ( .A(n_223), .B(n_277), .C(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_223), .B(n_248), .Y(n_287) );
OR2x2_ASAP7_75t_L g302 ( .A(n_223), .B(n_290), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_223), .B(n_257), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_223), .B(n_439), .Y(n_438) );
INVx5_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_224), .B(n_248), .Y(n_305) );
AND2x2_ASAP7_75t_L g344 ( .A(n_224), .B(n_258), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_224), .B(n_257), .Y(n_372) );
OR2x2_ASAP7_75t_L g375 ( .A(n_224), .B(n_257), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_227), .A2(n_501), .B(n_502), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_227), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_232), .A2(n_263), .B(n_265), .Y(n_262) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g489 ( .A(n_237), .Y(n_489) );
INVx5_ASAP7_75t_SL g290 ( .A(n_238), .Y(n_290) );
OR2x2_ASAP7_75t_L g296 ( .A(n_238), .B(n_247), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_238), .B(n_313), .Y(n_312) );
AOI321xp33_ASAP7_75t_L g319 ( .A1(n_238), .A2(n_320), .A3(n_321), .B1(n_322), .B2(n_328), .C(n_330), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_238), .B(n_246), .Y(n_329) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_238), .Y(n_342) );
OR2x2_ASAP7_75t_L g389 ( .A(n_238), .B(n_287), .Y(n_389) );
AND2x2_ASAP7_75t_L g411 ( .A(n_238), .B(n_308), .Y(n_411) );
AND2x2_ASAP7_75t_L g430 ( .A(n_238), .B(n_248), .Y(n_430) );
OR2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_257), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_248), .B(n_257), .Y(n_271) );
AND2x2_ASAP7_75t_L g280 ( .A(n_248), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
AND2x2_ASAP7_75t_L g313 ( .A(n_248), .B(n_308), .Y(n_313) );
INVxp67_ASAP7_75t_L g343 ( .A(n_248), .Y(n_343) );
OR2x2_ASAP7_75t_L g385 ( .A(n_248), .B(n_290), .Y(n_385) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_256), .Y(n_248) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_249), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_249), .A2(n_528), .B(n_535), .Y(n_527) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_249), .A2(n_537), .B(n_543), .Y(n_536) );
OR2x2_ASAP7_75t_L g267 ( .A(n_257), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g281 ( .A(n_257), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_257), .B(n_270), .Y(n_314) );
AND2x2_ASAP7_75t_L g363 ( .A(n_257), .B(n_307), .Y(n_363) );
AND2x2_ASAP7_75t_L g401 ( .A(n_257), .B(n_290), .Y(n_401) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_258), .B(n_290), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .B(n_272), .C(n_276), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_267), .A2(n_269), .B1(n_394), .B2(n_396), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_269), .A2(n_292), .B1(n_347), .B2(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_SL g421 ( .A(n_270), .Y(n_421) );
INVx1_ASAP7_75t_SL g321 ( .A(n_271), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_273), .B(n_293), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_314), .B1(n_321), .B2(n_335), .C1(n_339), .C2(n_345), .Y(n_334) );
AND2x2_ASAP7_75t_L g424 ( .A(n_273), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_274), .B(n_294), .Y(n_369) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_274), .Y(n_406) );
AND2x2_ASAP7_75t_L g409 ( .A(n_274), .B(n_318), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_274), .B(n_425), .Y(n_435) );
INVx1_ASAP7_75t_L g326 ( .A(n_275), .Y(n_326) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_275), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g417 ( .A1(n_277), .A2(n_418), .B(n_419), .C(n_422), .Y(n_417) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_279), .B(n_341), .C(n_344), .Y(n_340) );
OR2x2_ASAP7_75t_L g368 ( .A(n_279), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_279), .B(n_295), .Y(n_396) );
OR2x2_ASAP7_75t_L g301 ( .A(n_281), .B(n_302), .Y(n_301) );
AOI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B(n_291), .C(n_303), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_284), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g390 ( .A(n_285), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_286), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g304 ( .A(n_289), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_290), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g358 ( .A(n_290), .B(n_308), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_290), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_290), .B(n_307), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_296), .B1(n_297), .B2(n_301), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_293), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_296), .A2(n_360), .B1(n_362), .B2(n_364), .C(n_366), .Y(n_359) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g414 ( .A(n_299), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g427 ( .A(n_299), .B(n_416), .Y(n_427) );
INVx1_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
INVx1_ASAP7_75t_L g418 ( .A(n_301), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_302), .A2(n_385), .B(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .B(n_309), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI21xp5_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_314), .B(n_315), .Y(n_311) );
INVx1_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_313), .A2(n_399), .B1(n_402), .B2(n_404), .C(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_321), .A2(n_411), .B1(n_412), .B2(n_414), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g387 ( .A(n_323), .Y(n_387) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp67_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g391 ( .A(n_327), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g356 ( .A(n_332), .Y(n_356) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_337), .B(n_361), .Y(n_413) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_343), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g429 ( .A(n_344), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g436 ( .A(n_344), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI211xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_351), .B(n_352), .C(n_386), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_359), .C(n_378), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g439 ( .A(n_363), .Y(n_439) );
AND2x2_ASAP7_75t_L g376 ( .A(n_365), .B(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_374), .B2(n_376), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OR2x2_ASAP7_75t_L g384 ( .A(n_372), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g437 ( .A(n_373), .Y(n_437) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI31xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .A3(n_381), .B(n_384), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .C(n_393), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_395), .Y(n_394) );
NAND5xp2_ASAP7_75t_L g397 ( .A(n_398), .B(n_410), .C(n_417), .D(n_431), .E(n_434), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_409), .A2(n_435), .B1(n_436), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_SL g433 ( .A(n_411), .Y(n_433) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B(n_428), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g724 ( .A(n_447), .Y(n_724) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_455), .B1(n_458), .B2(n_721), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g726 ( .A(n_456), .Y(n_726) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR3x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_632), .C(n_679), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_578), .C(n_603), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_516), .B1(n_544), .B2(n_547), .C(n_555), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_484), .B(n_509), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_464), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_464), .B(n_560), .Y(n_676) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AND2x2_ASAP7_75t_L g546 ( .A(n_465), .B(n_515), .Y(n_546) );
AND2x2_ASAP7_75t_L g596 ( .A(n_465), .B(n_514), .Y(n_596) );
AND2x2_ASAP7_75t_L g617 ( .A(n_465), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g622 ( .A(n_465), .B(n_589), .Y(n_622) );
OR2x2_ASAP7_75t_L g630 ( .A(n_465), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g702 ( .A(n_465), .B(n_498), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_465), .B(n_651), .Y(n_716) );
INVx3_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g561 ( .A(n_466), .B(n_475), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_466), .B(n_498), .Y(n_562) );
AND2x4_ASAP7_75t_L g584 ( .A(n_466), .B(n_515), .Y(n_584) );
AND2x2_ASAP7_75t_L g614 ( .A(n_466), .B(n_486), .Y(n_614) );
AND2x2_ASAP7_75t_L g623 ( .A(n_466), .B(n_613), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_466), .B(n_499), .Y(n_639) );
OR2x2_ASAP7_75t_L g648 ( .A(n_466), .B(n_631), .Y(n_648) );
AND2x2_ASAP7_75t_L g654 ( .A(n_466), .B(n_589), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_466), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g668 ( .A(n_466), .B(n_511), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_466), .B(n_557), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_466), .B(n_618), .Y(n_707) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx2_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
AND2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_498), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_499), .Y(n_618) );
INVx1_ASAP7_75t_L g674 ( .A(n_475), .Y(n_674) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g583 ( .A(n_485), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_486), .B(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
OR2x2_ASAP7_75t_L g631 ( .A(n_486), .B(n_498), .Y(n_631) );
OR2x2_ASAP7_75t_L g692 ( .A(n_486), .B(n_599), .Y(n_692) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .B(n_497), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_488), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g512 ( .A(n_490), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_497), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_498), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g651 ( .A(n_498), .B(n_511), .Y(n_651) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_510), .A2(n_696), .B1(n_700), .B2(n_703), .C(n_704), .Y(n_695) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_SL g558 ( .A(n_511), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_511), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g690 ( .A(n_511), .B(n_546), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_514), .B(n_560), .Y(n_682) );
AND2x2_ASAP7_75t_L g589 ( .A(n_515), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g593 ( .A(n_516), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_516), .B(n_599), .Y(n_629) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
AND2x2_ASAP7_75t_L g554 ( .A(n_517), .B(n_527), .Y(n_554) );
INVx4_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
BUFx3_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
AND3x2_ASAP7_75t_L g624 ( .A(n_517), .B(n_625), .C(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g706 ( .A(n_526), .B(n_620), .Y(n_706) );
AND2x2_ASAP7_75t_L g714 ( .A(n_526), .B(n_599), .Y(n_714) );
INVx1_ASAP7_75t_SL g719 ( .A(n_526), .Y(n_719) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
INVx1_ASAP7_75t_SL g577 ( .A(n_527), .Y(n_577) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_566), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_527), .B(n_550), .Y(n_602) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_527), .Y(n_642) );
OR2x2_ASAP7_75t_L g647 ( .A(n_527), .B(n_566), .Y(n_647) );
INVx2_ASAP7_75t_L g552 ( .A(n_536), .Y(n_552) );
AND2x2_ASAP7_75t_L g587 ( .A(n_536), .B(n_567), .Y(n_587) );
OR2x2_ASAP7_75t_L g607 ( .A(n_536), .B(n_567), .Y(n_607) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_536), .Y(n_627) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_545), .A2(n_586), .B(n_678), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_547), .A2(n_557), .A3(n_584), .B1(n_714), .B2(n_715), .C1(n_717), .C2(n_720), .Y(n_713) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_549), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g644 ( .A(n_552), .B(n_566), .Y(n_644) );
AND2x2_ASAP7_75t_L g711 ( .A(n_552), .B(n_567), .Y(n_711) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g652 ( .A(n_554), .B(n_606), .Y(n_652) );
AOI31xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .A3(n_562), .B(n_563), .Y(n_555) );
AND2x2_ASAP7_75t_L g611 ( .A(n_557), .B(n_589), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_557), .B(n_581), .Y(n_693) );
AND2x2_ASAP7_75t_L g712 ( .A(n_557), .B(n_617), .Y(n_712) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_560), .B(n_589), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_560), .B(n_618), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_560), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_560), .B(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_561), .B(n_618), .Y(n_650) );
INVx1_ASAP7_75t_L g694 ( .A(n_561), .Y(n_694) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_576), .Y(n_564) );
INVxp67_ASAP7_75t_L g646 ( .A(n_565), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_566), .B(n_577), .Y(n_582) );
INVx1_ASAP7_75t_L g688 ( .A(n_566), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_566), .B(n_665), .Y(n_699) );
BUFx3_ASAP7_75t_L g599 ( .A(n_567), .Y(n_599) );
AND2x2_ASAP7_75t_L g625 ( .A(n_567), .B(n_577), .Y(n_625) );
INVx2_ASAP7_75t_L g665 ( .A(n_567), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_576), .B(n_698), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_585), .C(n_594), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_580), .A2(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_581), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_581), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g661 ( .A(n_582), .B(n_607), .Y(n_661) );
INVx3_ASAP7_75t_L g592 ( .A(n_584), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_588), .B1(n_591), .B2(n_593), .Y(n_585) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_587), .A2(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g636 ( .A(n_587), .B(n_600), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_587), .B(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g591 ( .A(n_590), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g660 ( .A(n_590), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_591), .A2(n_605), .B(n_610), .Y(n_604) );
OAI22xp33_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_597), .B1(n_601), .B2(n_602), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_596), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_615), .C(n_628), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g670 ( .A1(n_605), .A2(n_671), .B1(n_675), .B2(n_676), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g675 ( .A(n_607), .B(n_608), .Y(n_675) );
AND2x2_ASAP7_75t_L g683 ( .A(n_608), .B(n_664), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_SL g691 ( .A1(n_609), .A2(n_692), .B(n_693), .C(n_694), .Y(n_691) );
OR2x2_ASAP7_75t_L g718 ( .A(n_609), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_621), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_617), .A2(n_654), .B(n_655), .C(n_658), .Y(n_653) );
OAI21xp33_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g686 ( .A(n_625), .B(n_644), .Y(n_686) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_627), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_629), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_633), .B(n_653), .C(n_666), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_637), .C(n_645), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g663 ( .A(n_642), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_642), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_648), .C(n_649), .Y(n_645) );
INVx2_ASAP7_75t_SL g657 ( .A(n_647), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_648), .A2(n_659), .B1(n_661), .B2(n_662), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_670), .C(n_677), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g720 ( .A(n_674), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_695), .C(n_708), .D(n_713), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B(n_684), .C(n_691), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_689), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_685), .A2(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_692), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g728 ( .A(n_721), .Y(n_728) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
endmodule