module fake_jpeg_14157_n_138 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_29),
.A2(n_35),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_30),
.B(n_32),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_6),
.B1(n_8),
.B2(n_14),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_23),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_20),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_37),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_74),
.B(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_11),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_11),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_72),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_31),
.A2(n_28),
.B1(n_20),
.B2(n_15),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_42),
.B(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_38),
.B(n_24),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_86),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_74),
.B1(n_69),
.B2(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_84),
.B1(n_87),
.B2(n_70),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_31),
.B(n_52),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_45),
.C(n_34),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_22),
.B1(n_49),
.B2(n_12),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_12),
.B(n_6),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_12),
.B1(n_63),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_93),
.B1(n_81),
.B2(n_70),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_12),
.B1(n_58),
.B2(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_58),
.C(n_77),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_101),
.B1(n_84),
.B2(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_95),
.B1(n_80),
.B2(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_61),
.C(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_59),
.C(n_88),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_79),
.C(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_114),
.C(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_86),
.C(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_55),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_106),
.C(n_98),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_125),
.C(n_96),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_107),
.A3(n_102),
.B1(n_97),
.B2(n_108),
.C1(n_90),
.C2(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_107),
.C(n_108),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_124),
.B1(n_119),
.B2(n_65),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_128),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_77),
.C(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_65),
.B1(n_64),
.B2(n_68),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_65),
.B(n_131),
.Y(n_135)
);

AOI21x1_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_127),
.B(n_68),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_134),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_135),
.B(n_133),
.Y(n_138)
);


endmodule