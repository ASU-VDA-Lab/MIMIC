module real_jpeg_18445_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_487),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_0),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_1),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_1),
.B(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_1),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_2),
.Y(n_488)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_3),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_3),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_4),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_4),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_5),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_5),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_63),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_5),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_6),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_6),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_6),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_6),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_6),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_6),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_6),
.B(n_455),
.Y(n_454)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_7),
.Y(n_215)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_7),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g458 ( 
.A(n_7),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_8),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_8),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_9),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_173),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_9),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_9),
.B(n_432),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g440 ( 
.A(n_9),
.B(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_10),
.Y(n_447)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_11),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_12),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_12),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_12),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_12),
.B(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_12),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_12),
.B(n_213),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_14),
.B(n_85),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_14),
.B(n_139),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_14),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_14),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_14),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_14),
.B(n_407),
.Y(n_406)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_15),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_63),
.Y(n_62)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_16),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_16),
.B(n_172),
.Y(n_171)
);

NAND2x2_ASAP7_75t_SL g222 ( 
.A(n_16),
.B(n_223),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_17),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_178),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_R g20 ( 
.A(n_21),
.B(n_177),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_153),
.Y(n_22)
);

NOR2x1_ASAP7_75t_SL g177 ( 
.A(n_23),
.B(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_113),
.C(n_128),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_24),
.A2(n_25),
.B1(n_113),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_75),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_26),
.B(n_77),
.C(n_95),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.C(n_59),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_27),
.B(n_44),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

INVxp33_ASAP7_75t_SL g127 ( 
.A(n_28),
.Y(n_127)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_39),
.B(n_43),
.C(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_39),
.B(n_171),
.C(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_39),
.A2(n_42),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_41),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.C(n_55),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_45),
.A2(n_46),
.B1(n_55),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_49),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_50),
.B(n_120),
.Y(n_279)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_131),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_51),
.B(n_121),
.C(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_57),
.Y(n_258)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2x2_ASAP7_75t_SL g187 ( 
.A(n_59),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_67),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_65),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_61),
.B(n_66),
.C(n_67),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_61),
.B(n_115),
.C(n_121),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_61),
.B(n_255),
.C(n_257),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_61),
.A2(n_65),
.B1(n_255),
.B2(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_66),
.B1(n_80),
.B2(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_62),
.B(n_212),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_64),
.Y(n_401)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_64),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_80),
.C(n_84),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_73),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_73),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_95),
.B2(n_96),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.C(n_90),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_145),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_80),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_80),
.A2(n_135),
.B1(n_143),
.B2(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_80),
.B(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_86),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_148),
.C(n_151),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_90),
.A2(n_91),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_90),
.A2(n_91),
.B1(n_151),
.B2(n_152),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_94),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_94),
.Y(n_284)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_110),
.C(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_105),
.B(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_108),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_149),
.C(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_110),
.A2(n_111),
.B1(n_150),
.B2(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_125),
.C(n_126),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_121),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_122),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_144),
.C(n_147),
.Y(n_128)
);

XOR2x1_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_141),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_130),
.B(n_133),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_135),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_135),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_135),
.A2(n_193),
.B1(n_247),
.B2(n_248),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_140),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_140),
.A2(n_290),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_141),
.B(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_143),
.B(n_406),
.Y(n_413)
);

XNOR2x1_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_147),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_171),
.A2(n_175),
.B1(n_195),
.B2(n_196),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_225),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_185),
.B(n_187),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_189),
.B(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_203),
.C(n_206),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_190),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_200),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_191),
.B(n_194),
.Y(n_309)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g308 ( 
.A(n_200),
.B(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_355)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.C(n_222),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_208),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_216),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_209),
.B(n_212),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_214),
.Y(n_403)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_216),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_218),
.A2(n_222),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_218),
.Y(n_315)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_220),
.Y(n_441)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_222),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_371),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_348),
.B(n_362),
.C(n_363),
.D(n_370),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_320),
.B(n_347),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_305),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_231),
.B(n_305),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_277),
.C(n_298),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_232),
.B(n_322),
.Y(n_321)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_259),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_260),
.C(n_263),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_245),
.C(n_254),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_234),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJx3_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_238),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_242),
.B(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_245),
.A2(n_246),
.B1(n_254),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_257),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_269),
.C(n_274),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_298),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_289),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_280),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_285),
.B(n_288),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_474),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_291),
.Y(n_474)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_302),
.C(n_304),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_308),
.C(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_311),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_318),
.C(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_323),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.C(n_331),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_324),
.A2(n_325),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_327),
.A2(n_328),
.B1(n_331),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_331),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.C(n_336),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_332),
.B(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_335),
.B(n_336),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.C(n_346),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_337),
.A2(n_338),
.B1(n_346),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2x2_ASAP7_75t_L g424 ( 
.A(n_342),
.B(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_346),
.Y(n_426)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_349),
.B(n_364),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_360),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_360),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_356),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_366),
.C(n_367),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_368),
.Y(n_370)
);

NAND4xp25_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.D(n_375),
.Y(n_371)
);

OAI21x1_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_480),
.B(n_486),
.Y(n_375)
);

AOI21x1_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_468),
.B(n_479),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_427),
.B(n_467),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_411),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_379),
.B(n_411),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_397),
.C(n_404),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_380),
.B(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_381),
.B(n_393),
.C(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_393),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_397),
.A2(n_404),
.B1(n_405),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_402),
.Y(n_437)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_421),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_422),
.C(n_424),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_413),
.B(n_416),
.C(n_419),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_419),
.B2(n_420),
.Y(n_414)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_461),
.B(n_466),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_448),
.B(n_460),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_436),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_430),
.B(n_436),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_435),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_440),
.C(n_442),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_442),
.B2(n_443),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_453),
.B(n_459),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_452),
.Y(n_459)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx6_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_463),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_478),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g479 ( 
.A(n_469),
.B(n_478),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_476),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_475),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_475),
.C(n_476),
.Y(n_481)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);


endmodule