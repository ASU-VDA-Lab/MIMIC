module fake_netlist_6_3880_n_134 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_134);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_134;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_20),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_6),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_11),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_23),
.B(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_32),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_13),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_10),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_19),
.B(n_9),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_35),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_44),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_39),
.B(n_43),
.C(n_47),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_38),
.C(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_35),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_45),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_40),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_35),
.B(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AO21x2_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_55),
.B(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_65),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_67),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_75),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_94),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_88),
.Y(n_105)
);

OAI211xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_37),
.B(n_43),
.C(n_101),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_91),
.B1(n_89),
.B2(n_43),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_40),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

AOI222xp33_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_49),
.B1(n_64),
.B2(n_71),
.C1(n_69),
.C2(n_73),
.Y(n_123)
);

NOR4xp25_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_71),
.C(n_73),
.D(n_63),
.Y(n_124)
);

OAI211xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_70),
.B(n_73),
.C(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_63),
.C(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_119),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_116),
.B(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_118),
.Y(n_133)
);

OAI221xp5_ASAP7_75t_R g134 ( 
.A1(n_133),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.C(n_128),
.Y(n_134)
);


endmodule