module fake_jpeg_11223_n_476 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_4),
.B(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_50),
.Y(n_99)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_51),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_2),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_1),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_72),
.Y(n_127)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_77),
.Y(n_121)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_43),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_95),
.B(n_101),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_29),
.B1(n_33),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_98),
.A2(n_113),
.B1(n_129),
.B2(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_103),
.B(n_110),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_50),
.A2(n_29),
.B1(n_43),
.B2(n_23),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_107),
.A2(n_143),
.B(n_92),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_24),
.B1(n_39),
.B2(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_116),
.B(n_124),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_31),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_31),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_18),
.B1(n_20),
.B2(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_48),
.B(n_41),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_145),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_38),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_8),
.C(n_11),
.Y(n_184)
);

OR2x4_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_35),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_12),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_59),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_63),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_7),
.Y(n_177)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_153),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_93),
.A2(n_75),
.B1(n_74),
.B2(n_68),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_151),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_36),
.B(n_35),
.C(n_23),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_152),
.A2(n_158),
.B(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_35),
.B1(n_23),
.B2(n_22),
.Y(n_154)
);

AOI22x1_ASAP7_75t_L g242 ( 
.A1(n_154),
.A2(n_193),
.B1(n_199),
.B2(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_22),
.B(n_20),
.C(n_18),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_159),
.A2(n_165),
.B1(n_167),
.B2(n_174),
.Y(n_228)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_161),
.A2(n_168),
.B1(n_199),
.B2(n_186),
.Y(n_253)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_15),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_180),
.Y(n_209)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_90),
.Y(n_171)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_115),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_172),
.A2(n_104),
.B1(n_109),
.B2(n_187),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_151),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_97),
.B(n_15),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_184),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_177),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_195),
.B(n_127),
.Y(n_212)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_185),
.Y(n_213)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_89),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_196),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_106),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_12),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_100),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_13),
.B1(n_15),
.B2(n_136),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_112),
.A2(n_108),
.B1(n_142),
.B2(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_197),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_114),
.A2(n_102),
.B1(n_142),
.B2(n_91),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_96),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_122),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_117),
.A2(n_120),
.B1(n_139),
.B2(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_141),
.B(n_99),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_127),
.Y(n_223)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_217),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_208),
.A2(n_235),
.B1(n_253),
.B2(n_219),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_139),
.B1(n_133),
.B2(n_118),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_218),
.B1(n_237),
.B2(n_244),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_212),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_118),
.B1(n_141),
.B2(n_122),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_148),
.A2(n_96),
.B(n_130),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_219),
.A2(n_229),
.B(n_210),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_104),
.B(n_114),
.C(n_132),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_221),
.B(n_223),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_148),
.A2(n_132),
.B(n_104),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_135),
.C(n_102),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_193),
.C(n_198),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_188),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_238),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_166),
.B1(n_196),
.B2(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_181),
.B(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_156),
.B(n_164),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_245),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_240),
.B1(n_221),
.B2(n_251),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_184),
.B1(n_154),
.B2(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_175),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_160),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_154),
.A2(n_193),
.B1(n_180),
.B2(n_171),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_218),
.B1(n_211),
.B2(n_244),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_162),
.B(n_182),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_250),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_169),
.B(n_185),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_149),
.B(n_157),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_248),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_260),
.C(n_264),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_258),
.B(n_268),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_208),
.A2(n_176),
.B1(n_158),
.B2(n_152),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_263),
.B1(n_266),
.B2(n_274),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_190),
.C(n_226),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_262),
.A2(n_267),
.B1(n_277),
.B2(n_288),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_208),
.A2(n_240),
.B1(n_226),
.B2(n_242),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_236),
.C(n_205),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_242),
.B1(n_214),
.B2(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_224),
.B1(n_242),
.B2(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_205),
.B(n_224),
.C(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_276),
.C(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_205),
.B(n_224),
.C(n_207),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_221),
.B1(n_214),
.B2(n_207),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_235),
.A2(n_212),
.B1(n_223),
.B2(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_222),
.A2(n_239),
.B1(n_229),
.B2(n_228),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_225),
.Y(n_285)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_241),
.B1(n_206),
.B2(n_215),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_205),
.B(n_233),
.C(n_209),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_233),
.A2(n_249),
.B1(n_215),
.B2(n_225),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_233),
.A2(n_209),
.B1(n_220),
.B2(n_234),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_296),
.Y(n_318)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_227),
.A2(n_213),
.A3(n_250),
.B1(n_230),
.B2(n_233),
.Y(n_292)
);

AOI32xp33_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_291),
.A3(n_282),
.B1(n_289),
.B2(n_271),
.Y(n_315)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_213),
.Y(n_294)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_230),
.C(n_220),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_282),
.C(n_279),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_216),
.B(n_210),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_216),
.B(n_251),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_156),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_269),
.B(n_267),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_307),
.B(n_314),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_262),
.A2(n_255),
.B1(n_263),
.B2(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_306),
.A2(n_326),
.B1(n_323),
.B2(n_302),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_254),
.B(n_257),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_264),
.B(n_270),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_300),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_280),
.B(n_284),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_308),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_259),
.A2(n_273),
.B(n_255),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_265),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_320),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_276),
.A2(n_260),
.B(n_287),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_273),
.A2(n_299),
.B1(n_272),
.B2(n_271),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_289),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_333),
.B(n_336),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_303),
.C(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_256),
.A2(n_295),
.B(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_SL g335 ( 
.A(n_286),
.B(n_261),
.C(n_293),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_SL g349 ( 
.A(n_335),
.B(n_337),
.C(n_309),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_286),
.A2(n_275),
.B(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_322),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_318),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_343),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_328),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_310),
.Y(n_347)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_300),
.A2(n_330),
.B1(n_301),
.B2(n_309),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_306),
.B1(n_323),
.B2(n_305),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_349),
.A2(n_362),
.B1(n_364),
.B2(n_352),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_303),
.C(n_325),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_353),
.C(n_359),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_331),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_352),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_304),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_329),
.B(n_320),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_357),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_314),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_356),
.A2(n_347),
.B(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_310),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_307),
.C(n_321),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_338),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_371),
.C(n_359),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_360),
.Y(n_394)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_308),
.B(n_312),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_365),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_312),
.B(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_330),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_369),
.A2(n_305),
.B1(n_335),
.B2(n_304),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_302),
.B(n_336),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_370),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_376),
.B1(n_387),
.B2(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_316),
.B(n_327),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_383),
.B(n_388),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_348),
.A2(n_316),
.B1(n_322),
.B2(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_381),
.B(n_394),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_349),
.A2(n_339),
.B(n_364),
.C(n_370),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_398),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_350),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_369),
.Y(n_388)
);

OA21x2_ASAP7_75t_SL g391 ( 
.A1(n_344),
.A2(n_371),
.B(n_368),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_358),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_396),
.B(n_341),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_366),
.A2(n_340),
.B(n_361),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_340),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_392),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_410),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_353),
.C(n_345),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_417),
.C(n_398),
.Y(n_431)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_381),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_408),
.Y(n_421)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_411),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_345),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_413),
.Y(n_430)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_416),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_420),
.Y(n_422)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_367),
.C(n_358),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_419),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_362),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_391),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_377),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_428),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_386),
.B1(n_372),
.B2(n_399),
.Y(n_427)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_377),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_373),
.B1(n_372),
.B2(n_382),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_431),
.B(n_435),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_376),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_417),
.C(n_415),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_375),
.C(n_395),
.Y(n_435)
);

AO22x1_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_383),
.B1(n_374),
.B2(n_387),
.Y(n_437)
);

FAx1_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_383),
.CI(n_388),
.CON(n_447),
.SN(n_447)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_418),
.A2(n_388),
.B1(n_378),
.B2(n_383),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_438),
.A2(n_405),
.B1(n_408),
.B2(n_424),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_421),
.B(n_404),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_448),
.C(n_451),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_426),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_445),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_434),
.B1(n_437),
.B2(n_378),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_404),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_436),
.B1(n_384),
.B2(n_433),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_447),
.A2(n_383),
.B(n_422),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_403),
.C(n_407),
.Y(n_448)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_407),
.C(n_416),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_438),
.B1(n_424),
.B2(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g461 ( 
.A(n_454),
.B(n_455),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_460),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_421),
.C(n_425),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_459),
.A2(n_442),
.B(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_462),
.A2(n_463),
.B(n_453),
.Y(n_468)
);

NOR4xp25_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_428),
.C(n_449),
.D(n_440),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_451),
.C(n_439),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_453),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_469),
.C(n_464),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_468),
.A2(n_470),
.B(n_461),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_439),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_460),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_471),
.A2(n_472),
.B(n_458),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_458),
.B(n_455),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_474),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_469),
.Y(n_476)
);


endmodule