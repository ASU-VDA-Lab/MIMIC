module fake_netlist_1_3599_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
BUFx8_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_0), .B(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_15), .B(n_0), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
OA21x2_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_12), .B(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_19), .B(n_11), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_21), .B(n_20), .Y(n_24) );
OAI32xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .A3(n_20), .B1(n_17), .B2(n_4), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI221xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_13), .B1(n_17), .B2(n_11), .C(n_20), .Y(n_27) );
BUFx8_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
AND4x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .C(n_2), .D(n_3), .Y(n_29) );
NOR3xp33_ASAP7_75t_L g30 ( .A(n_28), .B(n_20), .C(n_2), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_20), .B1(n_13), .B2(n_3), .Y(n_33) );
AOI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_31), .B1(n_1), .B2(n_6), .Y(n_34) );
endmodule