module real_aes_1464_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_0), .A2(n_14), .B(n_15), .Y(n_13) );
AOI21xp33_ASAP7_75t_SL g17 ( .A1(n_0), .A2(n_1), .B(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g24 ( .A(n_1), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_2), .B(n_12), .Y(n_16) );
O2A1O1Ixp33_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_7), .B(n_17), .C(n_18), .Y(n_6) );
NOR2xp33_ASAP7_75t_SL g23 ( .A(n_3), .B(n_24), .Y(n_23) );
AND3x1_ASAP7_75t_L g26 ( .A(n_4), .B(n_5), .C(n_15), .Y(n_26) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_12), .B(n_13), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_SL g18 ( .A(n_19), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_21), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_22), .B(n_25), .Y(n_21) );
CKINVDCx16_ASAP7_75t_R g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
endmodule