module fake_jpeg_8002_n_308 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_52),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_65),
.B1(n_23),
.B2(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_20),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_13),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_35),
.B1(n_28),
.B2(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_36),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_65)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_74),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_83),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_75),
.Y(n_111)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_21),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_30),
.B(n_21),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_0),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_0),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_24),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_12),
.C(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_24),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_79),
.B1(n_95),
.B2(n_71),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_33),
.B1(n_31),
.B2(n_36),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_57),
.B1(n_55),
.B2(n_36),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_124),
.B1(n_45),
.B2(n_101),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_45),
.B1(n_66),
.B2(n_34),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_77),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_80),
.C(n_69),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_130),
.C(n_92),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_21),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_98),
.B1(n_86),
.B2(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_144),
.B1(n_155),
.B2(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_138),
.Y(n_167)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_83),
.B(n_92),
.C(n_77),
.D(n_70),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_104),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_72),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_89),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_75),
.B1(n_85),
.B2(n_68),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_67),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_152),
.B1(n_153),
.B2(n_108),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_115),
.C(n_113),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_74),
.B1(n_94),
.B2(n_81),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_73),
.B1(n_31),
.B2(n_33),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_91),
.B(n_64),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_33),
.B1(n_36),
.B2(n_42),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_0),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_110),
.B(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_91),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_106),
.A2(n_114),
.B(n_111),
.C(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_114),
.A3(n_109),
.B1(n_151),
.B2(n_135),
.C1(n_138),
.C2(n_163),
.Y(n_166)
);

OA21x2_ASAP7_75t_SL g213 ( 
.A1(n_166),
.A2(n_173),
.B(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_114),
.B(n_109),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_180),
.B(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

OA21x2_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_107),
.B(n_105),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_7),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_91),
.B(n_116),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_146),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_192),
.C(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_119),
.B(n_87),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_194),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_119),
.B(n_87),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_5),
.B(n_7),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_117),
.B1(n_2),
.B2(n_3),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_140),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_137),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_133),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_165),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_211),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_219),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_180),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_10),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_177),
.CI(n_171),
.CON(n_221),
.SN(n_221)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_235),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_205),
.B(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_217),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_183),
.B(n_189),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_216),
.B(n_207),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_169),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_218),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_256),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_251),
.B(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_173),
.B1(n_220),
.B2(n_185),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_254),
.B1(n_191),
.B2(n_219),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_206),
.C(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_257),
.C(n_259),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_212),
.B1(n_182),
.B2(n_191),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_166),
.B1(n_194),
.B2(n_186),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_197),
.B1(n_210),
.B2(n_190),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_164),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_231),
.B(n_178),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_197),
.C(n_164),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_261),
.B(n_268),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_223),
.B(n_239),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_271),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_209),
.B1(n_240),
.B2(n_237),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_249),
.B1(n_242),
.B2(n_241),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_215),
.B(n_196),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_250),
.C(n_259),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_225),
.C(n_187),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_266),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_182),
.B1(n_165),
.B2(n_193),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_257),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_284),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_187),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_282),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_268),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_283),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_271),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_267),
.B1(n_272),
.B2(n_265),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_291),
.B1(n_11),
.B2(n_15),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_178),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_292),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_269),
.B1(n_221),
.B2(n_225),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_15),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_16),
.C(n_285),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_16),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_293),
.Y(n_301)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_302),
.B(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_303),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_296),
.B1(n_304),
.B2(n_285),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_307),
.Y(n_308)
);


endmodule