module fake_jpeg_9813_n_208 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_23),
.B1(n_35),
.B2(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_24),
.B1(n_31),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_17),
.B2(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_18),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_23),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_19),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_71),
.B(n_18),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_35),
.B1(n_29),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_84),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_89),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_33),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_46),
.B(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_42),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_46),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_59),
.B1(n_74),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_80),
.B1(n_79),
.B2(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_107),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_46),
.B(n_42),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_117),
.C(n_4),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_84),
.B1(n_81),
.B2(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_111),
.B1(n_90),
.B2(n_3),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_59),
.B1(n_74),
.B2(n_44),
.Y(n_111)
);

NOR2x1p5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_48),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_95),
.B(n_94),
.C(n_75),
.D(n_93),
.Y(n_125)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_1),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_5),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_48),
.B(n_3),
.C(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_2),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_99),
.B1(n_124),
.B2(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_127),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_133),
.B1(n_144),
.B2(n_114),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_83),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_104),
.C(n_116),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_75),
.B1(n_80),
.B2(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_103),
.B1(n_120),
.B2(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_132),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_136),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_9),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_4),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_5),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_123),
.B(n_122),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_108),
.B(n_119),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_158),
.B(n_142),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_136),
.B1(n_125),
.B2(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_159),
.C(n_144),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_104),
.C(n_111),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_117),
.B1(n_10),
.B2(n_6),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_149),
.B1(n_152),
.B2(n_150),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_171),
.B1(n_161),
.B2(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_142),
.B1(n_148),
.B2(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_168),
.B1(n_162),
.B2(n_171),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.C(n_146),
.Y(n_174)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_161),
.A3(n_147),
.B1(n_152),
.B2(n_154),
.C(n_159),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_180),
.B(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_164),
.B1(n_167),
.B2(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_174),
.C(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_183),
.B1(n_182),
.B2(n_165),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_196),
.Y(n_199)
);

NAND4xp25_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_181),
.C(n_173),
.D(n_156),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_197),
.B(n_183),
.Y(n_200)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_187),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_194),
.B(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_196),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_165),
.B1(n_186),
.B2(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_192),
.C(n_199),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_199),
.B(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_207),
.A2(n_203),
.B(n_193),
.Y(n_208)
);


endmodule