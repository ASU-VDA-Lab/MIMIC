module fake_jpeg_16057_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_65),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_42),
.B1(n_57),
.B2(n_52),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_73),
.B1(n_55),
.B2(n_44),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_38),
.B1(n_56),
.B2(n_47),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_51),
.B1(n_54),
.B2(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_103),
.Y(n_120)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_100),
.Y(n_124)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_43),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_112),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_3),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_114),
.B(n_4),
.Y(n_122)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_113),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_41),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_90),
.Y(n_132)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_111),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_116),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_120),
.B1(n_93),
.B2(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_150),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_106),
.B1(n_126),
.B2(n_97),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_109),
.B(n_129),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_127),
.B1(n_106),
.B2(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_149),
.B(n_41),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_151),
.B1(n_154),
.B2(n_60),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_25),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_27),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_23),
.C(n_37),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_21),
.B(n_36),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_20),
.B1(n_35),
.B2(n_8),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_28),
.B(n_31),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_91),
.C(n_17),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_15),
.C(n_29),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_14),
.Y(n_169)
);


endmodule