module fake_netlist_6_657_n_1825 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1825);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1825;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_86),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_40),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_118),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_28),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_69),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_83),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_58),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_57),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_44),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_5),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_139),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_44),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_40),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_94),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_109),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_48),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_33),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_9),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_63),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_80),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_29),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_141),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_21),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_45),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_70),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_102),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_68),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_91),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_93),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_19),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_98),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_42),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_90),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_140),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_1),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_136),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_43),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_31),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_159),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_25),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_96),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_9),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_81),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_51),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_60),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_129),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_36),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_134),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_59),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_74),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_71),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_99),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_53),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_158),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_106),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_100),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_145),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_103),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_41),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_22),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_161),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_18),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_1),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_61),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_25),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_7),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_115),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_58),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_88),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_41),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_116),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_35),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_95),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_53),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_17),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_11),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_19),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_105),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_62),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_49),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_37),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_51),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_89),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_65),
.Y(n_320)
);

CKINVDCx6p67_ASAP7_75t_R g321 ( 
.A(n_124),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_13),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_54),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_128),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_133),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_117),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_84),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_47),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_193),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_193),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_272),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_175),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_172),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_175),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_176),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_173),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_202),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_221),
.B(n_169),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_176),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_177),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_221),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_319),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_182),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_185),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_191),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_210),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_191),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_187),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_190),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_198),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_196),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_200),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_208),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_197),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_178),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_201),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_201),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_172),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_229),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_220),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_229),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_238),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_273),
.B(n_0),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_238),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_224),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_225),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_244),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_271),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_170),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_244),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_252),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_252),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_260),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_260),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_228),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_267),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_267),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_286),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_232),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_292),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_246),
.B(n_2),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_181),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_292),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_297),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_234),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_297),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_271),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_298),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_298),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_235),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_236),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_301),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_301),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_203),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_203),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_248),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_248),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_348),
.B(n_275),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_340),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_275),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_374),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_340),
.B(n_279),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_339),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_333),
.A2(n_281),
.B1(n_330),
.B2(n_258),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

AND3x2_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_264),
.C(n_216),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_335),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_343),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_375),
.B(n_296),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_338),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_356),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_338),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_349),
.B(n_296),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_361),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_366),
.B(n_279),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_367),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_371),
.Y(n_470)
);

BUFx8_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_351),
.B(n_179),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_398),
.B(n_281),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_379),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_382),
.B(n_170),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_435),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_337),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_458),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_425),
.B(n_179),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_424),
.B(n_342),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_435),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_344),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_425),
.B(n_350),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_353),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_479),
.B(n_354),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_425),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_458),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_479),
.B(n_359),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_413),
.B(n_386),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_413),
.B(n_386),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_456),
.B(n_360),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_448),
.B(n_362),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_448),
.B(n_364),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_458),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_457),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_473),
.A2(n_312),
.B1(n_316),
.B2(n_318),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_456),
.A2(n_365),
.B1(n_369),
.B2(n_380),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_415),
.B(n_180),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_413),
.B(n_415),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_387),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_450),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_457),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_436),
.A2(n_226),
.B1(n_219),
.B2(n_206),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_430),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_439),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_415),
.B(n_381),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_180),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_429),
.B(n_186),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_390),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_471),
.B(n_395),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_464),
.B(n_387),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_415),
.B(n_401),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_415),
.B(n_407),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_422),
.B(n_408),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

AO22x1_ASAP7_75t_L g550 ( 
.A1(n_464),
.A2(n_316),
.B1(n_318),
.B2(n_323),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_422),
.B(n_211),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_440),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_433),
.A2(n_195),
.B1(n_306),
.B2(n_247),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_422),
.B(n_170),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_422),
.B(n_240),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_471),
.B(n_174),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_422),
.B(n_250),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g563 ( 
.A(n_474),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_474),
.B(n_388),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_471),
.A2(n_268),
.B1(n_263),
.B2(n_289),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_189),
.C(n_186),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_421),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_462),
.Y(n_568)
);

INVx4_ASAP7_75t_SL g569 ( 
.A(n_484),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_434),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_439),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_431),
.B(n_251),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_464),
.B(n_254),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_419),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_442),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_450),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_434),
.B(n_345),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_471),
.B(n_174),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_451),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_451),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_454),
.B(n_434),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

AND2x2_ASAP7_75t_SL g589 ( 
.A(n_464),
.B(n_216),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_464),
.B(n_388),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_471),
.B(n_174),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_436),
.B(n_174),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_467),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_484),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_454),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_454),
.B(n_257),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_454),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_414),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_454),
.B(n_347),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_467),
.B(n_241),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_467),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_467),
.B(n_241),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_419),
.B(n_461),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_463),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_463),
.B(n_269),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_467),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_418),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_468),
.B(n_170),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_465),
.B(n_389),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_468),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_466),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_466),
.A2(n_242),
.B1(n_266),
.B2(n_239),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_468),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_472),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_418),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_418),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_472),
.A2(n_323),
.B1(n_324),
.B2(n_290),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_475),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_468),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_475),
.B(n_389),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_477),
.B(n_352),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_426),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_476),
.B(n_241),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_477),
.B(n_183),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_478),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_426),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_478),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_487),
.B(n_480),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_496),
.B(n_261),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_589),
.B(n_170),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_589),
.B(n_523),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_589),
.B(n_476),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_495),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_597),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_503),
.B(n_476),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_503),
.B(n_476),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_597),
.B(n_480),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_498),
.B(n_188),
.C(n_184),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_503),
.B(n_476),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_634),
.B(n_476),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_634),
.B(n_476),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_507),
.B(n_508),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_507),
.B(n_482),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_628),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_531),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_508),
.B(n_482),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_525),
.B(n_482),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_535),
.A2(n_328),
.B1(n_305),
.B2(n_302),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_510),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_603),
.B(n_482),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_525),
.B(n_482),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_521),
.B(n_482),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_628),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_521),
.B(n_486),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_532),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_533),
.B(n_189),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_510),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_601),
.A2(n_287),
.B1(n_270),
.B2(n_276),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_499),
.B(n_511),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_521),
.B(n_486),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_490),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_563),
.B(n_194),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_486),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_537),
.B(n_486),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_538),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_516),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_537),
.B(n_544),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_564),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_544),
.B(n_486),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_546),
.B(n_486),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_518),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_481),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_546),
.B(n_486),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_549),
.B(n_486),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_490),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_549),
.B(n_446),
.Y(n_695)
);

AO221x1_ASAP7_75t_L g696 ( 
.A1(n_555),
.A2(n_324),
.B1(n_207),
.B2(n_214),
.C(n_199),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_521),
.B(n_264),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_533),
.A2(n_284),
.B1(n_277),
.B2(n_280),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_548),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_552),
.B(n_446),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_535),
.A2(n_302),
.B1(n_290),
.B2(n_305),
.Y(n_701)
);

AND2x6_ASAP7_75t_SL g702 ( 
.A(n_582),
.B(n_391),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_550),
.B(n_192),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_554),
.B(n_446),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_520),
.B(n_204),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_446),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_529),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_548),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_493),
.B(n_328),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_561),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_630),
.B(n_481),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_535),
.A2(n_586),
.B1(n_543),
.B2(n_545),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_490),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_561),
.B(n_446),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_550),
.B(n_192),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_534),
.B(n_209),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_572),
.B(n_459),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_547),
.B(n_500),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_578),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_578),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_535),
.A2(n_299),
.B1(n_303),
.B2(n_308),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_579),
.B(n_459),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_579),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_580),
.B(n_459),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_580),
.B(n_584),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_584),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_586),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_585),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_502),
.B(n_213),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_585),
.B(n_460),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_493),
.B(n_314),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_501),
.B(n_294),
.C(n_223),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_493),
.B(n_327),
.Y(n_736)
);

AND2x6_ASAP7_75t_SL g737 ( 
.A(n_535),
.B(n_391),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_526),
.B(n_581),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_612),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_490),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_587),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_542),
.B(n_590),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_493),
.B(n_329),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_551),
.A2(n_505),
.B1(n_575),
.B2(n_598),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_596),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_596),
.B(n_460),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_576),
.A2(n_515),
.B1(n_512),
.B2(n_558),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_460),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_519),
.B(n_259),
.C(n_256),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_567),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_483),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_536),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_542),
.B(n_483),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_607),
.B(n_469),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_557),
.B(n_484),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_614),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_562),
.A2(n_199),
.B1(n_205),
.B2(n_207),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_614),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_619),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_619),
.B(n_469),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_622),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_557),
.B(n_484),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

AND2x6_ASAP7_75t_SL g766 ( 
.A(n_536),
.B(n_392),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_626),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_620),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_493),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_636),
.B(n_469),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_636),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_606),
.B(n_452),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_590),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_494),
.B(n_470),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_560),
.A2(n_426),
.B(n_485),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_494),
.B(n_470),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_494),
.B(n_470),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_494),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_514),
.B(n_452),
.Y(n_779)
);

O2A1O1Ixp5_ASAP7_75t_L g780 ( 
.A1(n_514),
.A2(n_233),
.B(n_326),
.C(n_320),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_514),
.B(n_485),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_536),
.A2(n_233),
.B1(n_205),
.B2(n_214),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_514),
.Y(n_783)
);

AND2x6_ASAP7_75t_SL g784 ( 
.A(n_536),
.B(n_392),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_571),
.B(n_215),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_536),
.B(n_485),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_497),
.Y(n_787)
);

AOI221xp5_ASAP7_75t_L g788 ( 
.A1(n_530),
.A2(n_565),
.B1(n_322),
.B2(n_317),
.C(n_313),
.Y(n_788)
);

AND3x1_ASAP7_75t_L g789 ( 
.A(n_530),
.B(n_625),
.C(n_394),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_602),
.A2(n_231),
.B(n_243),
.C(n_245),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_531),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_571),
.B(n_452),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_559),
.A2(n_591),
.B1(n_583),
.B2(n_540),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_522),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_571),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_566),
.A2(n_231),
.B1(n_243),
.B2(n_245),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_557),
.A2(n_326),
.B1(n_249),
.B2(n_255),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_489),
.B(n_452),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_489),
.A2(n_249),
.B(n_255),
.C(n_262),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_492),
.B(n_452),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_492),
.B(n_452),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_497),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_759),
.B(n_488),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_638),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_778),
.A2(n_642),
.B(n_680),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_639),
.B(n_504),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_778),
.A2(n_560),
.B(n_541),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_714),
.A2(n_560),
.B(n_541),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_682),
.B(n_571),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_685),
.B(n_570),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_638),
.B(n_557),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_719),
.B(n_712),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_685),
.B(n_570),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_793),
.A2(n_632),
.B1(n_605),
.B2(n_262),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_659),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_738),
.B(n_791),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_641),
.A2(n_541),
.B(n_491),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_699),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_713),
.B(n_745),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_641),
.A2(n_541),
.B(n_491),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_645),
.A2(n_652),
.B(n_646),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_640),
.A2(n_506),
.B(n_504),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_774),
.A2(n_777),
.B(n_776),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_638),
.B(n_644),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_706),
.A2(n_227),
.B(n_217),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_742),
.B(n_506),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_643),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_643),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_667),
.A2(n_574),
.B(n_491),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_651),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_667),
.A2(n_574),
.B(n_491),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_768),
.A2(n_283),
.B1(n_320),
.B2(n_282),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_795),
.B(n_513),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_640),
.A2(n_513),
.B(n_528),
.C(n_629),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_655),
.A2(n_557),
.B1(n_609),
.B2(n_629),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_661),
.A2(n_524),
.B(n_568),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_651),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_658),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_661),
.A2(n_524),
.B(n_568),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_669),
.A2(n_574),
.B(n_528),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_638),
.B(n_594),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_731),
.A2(n_265),
.B(n_282),
.C(n_283),
.Y(n_842)
);

BUFx8_ASAP7_75t_L g843 ( 
.A(n_709),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_649),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_659),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_754),
.B(n_517),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_R g847 ( 
.A(n_794),
.B(n_522),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_648),
.B(n_393),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_655),
.B(n_517),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_669),
.A2(n_574),
.B(n_613),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_696),
.A2(n_557),
.B1(n_265),
.B2(n_241),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_644),
.B(n_594),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_637),
.A2(n_788),
.B(n_689),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_539),
.B(n_577),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_644),
.A2(n_553),
.B1(n_627),
.B2(n_527),
.Y(n_855)
);

AOI33xp33_ASAP7_75t_L g856 ( 
.A1(n_739),
.A2(n_409),
.A3(n_393),
.B1(n_394),
.B2(n_396),
.B3(n_399),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_779),
.A2(n_577),
.B(n_527),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_649),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_729),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_729),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_666),
.A2(n_539),
.B(n_595),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_670),
.B(n_553),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_658),
.Y(n_863)
);

NOR2x1_ASAP7_75t_L g864 ( 
.A(n_734),
.B(n_556),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_677),
.B(n_556),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_717),
.A2(n_617),
.B(n_593),
.C(n_627),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_683),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_679),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_662),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_748),
.A2(n_613),
.B1(n_593),
.B2(n_621),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_704),
.B(n_595),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_604),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_664),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_647),
.B(n_594),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_676),
.A2(n_615),
.B(n_609),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_753),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_666),
.A2(n_604),
.B(n_615),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_773),
.A2(n_616),
.B(n_621),
.C(n_618),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_656),
.A2(n_616),
.B(n_618),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_664),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_721),
.B(n_617),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_647),
.B(n_594),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_781),
.A2(n_594),
.B(n_497),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_656),
.A2(n_594),
.B(n_610),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_693),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_725),
.B(n_730),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_746),
.B(n_588),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_796),
.A2(n_623),
.B(n_610),
.C(n_624),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_660),
.A2(n_623),
.B(n_610),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_757),
.B(n_588),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_660),
.A2(n_623),
.B(n_631),
.C(n_624),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_751),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_672),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_762),
.B(n_588),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_786),
.A2(n_635),
.B(n_631),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_735),
.A2(n_321),
.B1(n_237),
.B2(n_253),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_647),
.A2(n_321),
.B1(n_278),
.B2(n_285),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_657),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_672),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_795),
.B(n_230),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_668),
.A2(n_409),
.B(n_396),
.C(n_399),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_665),
.A2(n_635),
.B(n_631),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_711),
.B(n_569),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_751),
.Y(n_906)
);

INVx6_ASAP7_75t_L g907 ( 
.A(n_737),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_695),
.A2(n_635),
.B(n_631),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_785),
.B(n_400),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_711),
.B(n_569),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_794),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_752),
.A2(n_635),
.B(n_624),
.C(n_588),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_675),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_700),
.A2(n_624),
.B(n_600),
.Y(n_914)
);

AND2x2_ASAP7_75t_SL g915 ( 
.A(n_789),
.B(n_400),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_763),
.B(n_600),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_765),
.B(n_600),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_673),
.B(n_402),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_671),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_650),
.B(n_402),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_678),
.A2(n_600),
.B(n_449),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_678),
.A2(n_449),
.B(n_443),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_675),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_692),
.A2(n_449),
.B(n_443),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_750),
.A2(n_304),
.B(n_295),
.Y(n_925)
);

CKINVDCx10_ASAP7_75t_R g926 ( 
.A(n_702),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_557),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_684),
.B(n_428),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_688),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_727),
.B(n_291),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_692),
.A2(n_449),
.B(n_443),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_692),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_769),
.B(n_416),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_792),
.A2(n_611),
.B1(n_484),
.B2(n_443),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_722),
.B(n_428),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_740),
.Y(n_937)
);

BUFx4f_ASAP7_75t_L g938 ( 
.A(n_703),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_740),
.A2(n_449),
.B(n_428),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_671),
.B(n_404),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_694),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_740),
.A2(n_449),
.B(n_441),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_728),
.B(n_441),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_694),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_741),
.A2(n_760),
.B(n_767),
.C(n_744),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_741),
.B(n_405),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_772),
.A2(n_449),
.B(n_441),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_703),
.B(n_274),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_744),
.B(n_444),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_760),
.B(n_444),
.Y(n_951)
);

OA22x2_ASAP7_75t_L g952 ( 
.A1(n_703),
.A2(n_307),
.B1(n_311),
.B2(n_325),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_792),
.A2(n_416),
.B(n_423),
.C(n_420),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_705),
.A2(n_611),
.B(n_484),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_767),
.B(n_405),
.Y(n_955)
);

NOR2x1p5_ASAP7_75t_L g956 ( 
.A(n_766),
.B(n_411),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_663),
.B(n_708),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_772),
.A2(n_449),
.B(n_444),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_782),
.A2(n_406),
.B(n_410),
.Y(n_959)
);

NOR2x1_ASAP7_75t_R g960 ( 
.A(n_733),
.B(n_406),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_708),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_779),
.A2(n_445),
.B(n_417),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_703),
.B(n_410),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_653),
.A2(n_445),
.B(n_417),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_784),
.B(n_92),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_654),
.A2(n_423),
.B(n_420),
.Y(n_966)
);

NAND2x1_ASAP7_75t_L g967 ( 
.A(n_769),
.B(n_611),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_733),
.A2(n_445),
.B(n_452),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_736),
.A2(n_452),
.B(n_569),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_697),
.A2(n_411),
.B(n_315),
.C(n_274),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_736),
.A2(n_569),
.B(n_611),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_743),
.A2(n_611),
.B(n_484),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_718),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_698),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_743),
.A2(n_611),
.B(n_484),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_724),
.B(n_611),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_726),
.B(n_484),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_798),
.A2(n_484),
.B(n_137),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_732),
.B(n_315),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_800),
.A2(n_131),
.B(n_79),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_747),
.A2(n_315),
.B(n_274),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_801),
.A2(n_138),
.B(n_97),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_723),
.B(n_6),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_749),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_697),
.A2(n_142),
.B(n_111),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_769),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_769),
.B(n_315),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_707),
.B(n_274),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_828),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_812),
.A2(n_716),
.B1(n_758),
.B2(n_701),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_830),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_909),
.B(n_755),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_805),
.A2(n_823),
.B(n_819),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_869),
.B(n_761),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_819),
.A2(n_783),
.B(n_775),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_807),
.A2(n_756),
.B(n_764),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_869),
.B(n_770),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_SL g998 ( 
.A(n_825),
.B(n_790),
.C(n_799),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_931),
.B(n_715),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_815),
.B(n_799),
.C(n_710),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_843),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_931),
.B(n_802),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_827),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_983),
.A2(n_716),
.B(n_710),
.C(n_681),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_837),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_818),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_818),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_973),
.B(n_787),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_853),
.B(n_803),
.C(n_983),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_915),
.A2(n_716),
.B1(n_797),
.B2(n_691),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_844),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_804),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_816),
.B(n_690),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_843),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_838),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_863),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_956),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_984),
.B(n_687),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_915),
.B(n_686),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_986),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_957),
.A2(n_764),
.B(n_756),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_808),
.A2(n_780),
.B(n_164),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_844),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_947),
.B(n_7),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_809),
.B(n_162),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_938),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_1027)
);

OA21x2_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_157),
.B(n_155),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_809),
.B(n_10),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_867),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_817),
.A2(n_154),
.B(n_152),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_810),
.B(n_130),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_820),
.A2(n_126),
.B(n_123),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_886),
.B(n_120),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_947),
.B(n_12),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_874),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_844),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_887),
.B(n_15),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_821),
.A2(n_897),
.B(n_846),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_813),
.B(n_15),
.C(n_16),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_845),
.B(n_122),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_867),
.B(n_16),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_829),
.A2(n_119),
.B(n_64),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_831),
.A2(n_18),
.B(n_21),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_813),
.B(n_23),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_913),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_955),
.B(n_963),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_929),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_834),
.A2(n_24),
.B(n_26),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_930),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_900),
.B(n_24),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_929),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_886),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_946),
.A2(n_27),
.B(n_30),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_911),
.B(n_30),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_902),
.B(n_32),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_919),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_832),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_826),
.A2(n_39),
.B(n_46),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_928),
.A2(n_806),
.B(n_852),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_852),
.A2(n_46),
.B(n_50),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_859),
.B(n_50),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_919),
.A2(n_54),
.B(n_918),
.C(n_938),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_949),
.B(n_804),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_986),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_877),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_900),
.B(n_943),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_908),
.A2(n_914),
.B(n_811),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_860),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_842),
.A2(n_988),
.B(n_903),
.C(n_987),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_941),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_814),
.A2(n_979),
.B(n_960),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_883),
.B(n_976),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_870),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_925),
.B(n_898),
.C(n_899),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_920),
.A2(n_849),
.B(n_856),
.C(n_988),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_858),
.B(n_892),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_903),
.A2(n_987),
.B(n_940),
.C(n_877),
.Y(n_1080)
);

INVx8_ASAP7_75t_L g1081 ( 
.A(n_848),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_892),
.B(n_906),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_848),
.B(n_847),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_906),
.B(n_881),
.Y(n_1084)
);

NAND2x1p5_ASAP7_75t_L g1085 ( 
.A(n_894),
.B(n_875),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_895),
.B(n_901),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_894),
.B(n_833),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_974),
.A2(n_851),
.B1(n_933),
.B2(n_937),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_883),
.A2(n_841),
.B(n_850),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_952),
.B(n_907),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_905),
.A2(n_910),
.B(n_866),
.C(n_912),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_824),
.B(n_970),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_824),
.B(n_907),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_879),
.A2(n_854),
.B(n_876),
.C(n_835),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_907),
.B(n_967),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_952),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_893),
.A2(n_923),
.B(n_945),
.C(n_961),
.Y(n_1097)
);

INVxp67_ASAP7_75t_SL g1098 ( 
.A(n_933),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_937),
.B(n_981),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_905),
.A2(n_910),
.B(n_927),
.C(n_841),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_862),
.B(n_865),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_934),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_872),
.B(n_882),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_873),
.B(n_917),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_966),
.A2(n_871),
.B(n_855),
.C(n_822),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_888),
.B(n_891),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_857),
.A2(n_836),
.B(n_839),
.Y(n_1107)
);

OA22x2_ASAP7_75t_L g1108 ( 
.A1(n_959),
.A2(n_880),
.B1(n_861),
.B2(n_878),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_864),
.A2(n_916),
.B1(n_896),
.B2(n_977),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_936),
.A2(n_944),
.B(n_950),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_951),
.B(n_934),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_965),
.B(n_851),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_985),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_964),
.B(n_890),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_904),
.B(n_962),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_972),
.B(n_975),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_840),
.B(n_885),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_965),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_935),
.A2(n_889),
.B1(n_971),
.B2(n_954),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_SL g1120 ( 
.A1(n_884),
.A2(n_969),
.B(n_921),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_968),
.A2(n_982),
.B(n_980),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_953),
.B(n_978),
.C(n_926),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_958),
.A2(n_948),
.B(n_939),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_942),
.B(n_922),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_924),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_932),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_805),
.A2(n_778),
.B(n_642),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_827),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_818),
.Y(n_1129)
);

OAI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_812),
.A2(n_674),
.B(n_639),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_815),
.B(n_531),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_828),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_819),
.A2(n_640),
.B(n_842),
.C(n_641),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_805),
.A2(n_778),
.B(n_642),
.Y(n_1134)
);

AOI222xp33_ASAP7_75t_L g1135 ( 
.A1(n_983),
.A2(n_788),
.B1(n_592),
.B2(n_674),
.C1(n_424),
.C2(n_348),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_812),
.B(n_682),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_R g1137 ( 
.A(n_815),
.B(n_531),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_983),
.B(n_674),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_L g1139 ( 
.A(n_844),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_812),
.B(n_674),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1008),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1007),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1070),
.A2(n_1040),
.B(n_993),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1127),
.A2(n_1134),
.B(n_1062),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1133),
.A2(n_999),
.B(n_1103),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1138),
.A2(n_1130),
.B(n_1010),
.C(n_1029),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1138),
.A2(n_1135),
.B1(n_1136),
.B2(n_1140),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_SL g1148 ( 
.A(n_1135),
.B(n_1077),
.C(n_1131),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_989),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_1105),
.A2(n_1107),
.B(n_1051),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1048),
.B(n_992),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_995),
.A2(n_1119),
.B(n_1117),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1101),
.A2(n_1003),
.B(n_1104),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1121),
.A2(n_1094),
.A3(n_1119),
.B(n_1023),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1021),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_991),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1106),
.A2(n_1114),
.B(n_1115),
.Y(n_1157)
);

AO32x2_ASAP7_75t_L g1158 ( 
.A1(n_1027),
.A2(n_1088),
.A3(n_990),
.B1(n_1011),
.B2(n_1056),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_1051),
.A2(n_1056),
.B(n_1097),
.Y(n_1159)
);

NOR2xp67_ASAP7_75t_SL g1160 ( 
.A(n_1050),
.B(n_1021),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1075),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1113),
.A2(n_1124),
.B(n_1019),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1016),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1095),
.B(n_1083),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1139),
.B(n_1021),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_1109),
.A2(n_1045),
.B(n_1078),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1030),
.B(n_1069),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_994),
.B(n_997),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1017),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1005),
.A2(n_1020),
.B(n_1022),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1058),
.C(n_1080),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1002),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1110),
.A2(n_996),
.B(n_1108),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1113),
.A2(n_1108),
.B(n_1021),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1129),
.B(n_1071),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1026),
.A2(n_1065),
.B(n_1032),
.C(n_1059),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1037),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1014),
.B(n_1039),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1009),
.B(n_1112),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1031),
.A2(n_1033),
.B(n_1116),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1139),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1096),
.A2(n_1046),
.B1(n_1090),
.B2(n_1081),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1018),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1049),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1113),
.A2(n_1092),
.B(n_1091),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_1044),
.B(n_1086),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1068),
.B(n_1093),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1047),
.Y(n_1188)
);

AND2x6_ASAP7_75t_L g1189 ( 
.A(n_1034),
.B(n_1067),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1052),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1060),
.A2(n_1053),
.B(n_1064),
.C(n_1043),
.Y(n_1191)
);

AO32x2_ASAP7_75t_L g1192 ( 
.A1(n_990),
.A2(n_1011),
.A3(n_1000),
.B1(n_1092),
.B2(n_1041),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_1035),
.B1(n_1093),
.B2(n_1066),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1073),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1137),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1120),
.A2(n_998),
.B(n_1111),
.Y(n_1196)
);

INVx5_ASAP7_75t_L g1197 ( 
.A(n_1055),
.Y(n_1197)
);

AOI31xp67_ASAP7_75t_L g1198 ( 
.A1(n_1004),
.A2(n_1036),
.A3(n_1128),
.B(n_1006),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1132),
.B(n_1076),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_1061),
.A2(n_1066),
.B(n_1063),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1113),
.A2(n_1100),
.B(n_1087),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1001),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1084),
.A2(n_1079),
.A3(n_1028),
.B(n_1099),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1122),
.B(n_1057),
.C(n_1034),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1081),
.A2(n_1098),
.B(n_1013),
.C(n_1067),
.Y(n_1205)
);

OAI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1042),
.A2(n_1118),
.B(n_1095),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1118),
.B(n_1095),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1102),
.B(n_1081),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1028),
.A2(n_1126),
.A3(n_1054),
.B(n_1085),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1082),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1002),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1002),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1012),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1055),
.B(n_1012),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1055),
.B(n_1038),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1024),
.A2(n_1078),
.B(n_819),
.C(n_1026),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1015),
.A2(n_1024),
.B(n_1038),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1024),
.B(n_1038),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_SL g1219 ( 
.A(n_1050),
.B(n_738),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_989),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1138),
.A2(n_1135),
.B1(n_1010),
.B2(n_674),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1121),
.A2(n_993),
.A3(n_1094),
.B(n_1119),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1140),
.B(n_812),
.Y(n_1226)
);

BUFx4f_ASAP7_75t_SL g1227 ( 
.A(n_1050),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1135),
.A2(n_674),
.B(n_788),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1070),
.A2(n_819),
.B(n_1062),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1138),
.A2(n_1135),
.B(n_639),
.C(n_674),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1008),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1140),
.B(n_812),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1070),
.A2(n_819),
.B(n_1062),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_989),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_989),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1140),
.B(n_812),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1008),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1121),
.A2(n_993),
.A3(n_1094),
.B(n_1119),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1008),
.Y(n_1240)
);

AND2x2_ASAP7_75t_SL g1241 ( 
.A(n_1138),
.B(n_1010),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_1043),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1127),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1008),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1130),
.A2(n_639),
.B(n_674),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1140),
.B(n_487),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1129),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1078),
.A2(n_819),
.B(n_1026),
.C(n_1065),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1070),
.A2(n_819),
.B(n_1040),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1140),
.B(n_487),
.Y(n_1252)
);

AO32x2_ASAP7_75t_L g1253 ( 
.A1(n_1027),
.A2(n_832),
.A3(n_1088),
.B1(n_1119),
.B2(n_990),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1138),
.A2(n_1135),
.B1(n_1010),
.B2(n_674),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1140),
.B(n_812),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_989),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1121),
.A2(n_993),
.A3(n_1094),
.B(n_1119),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1008),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_989),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1127),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1008),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1127),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1138),
.A2(n_1135),
.B(n_639),
.C(n_674),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1005),
.A2(n_819),
.B(n_778),
.Y(n_1266)
);

NAND2x1_ASAP7_75t_L g1267 ( 
.A(n_1067),
.B(n_986),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_989),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1021),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1056),
.A2(n_1080),
.B(n_1072),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1138),
.B(n_682),
.Y(n_1271)
);

BUFx8_ASAP7_75t_SL g1272 ( 
.A(n_1001),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1105),
.A2(n_993),
.B(n_1070),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1140),
.B(n_812),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1095),
.B(n_1083),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_989),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1127),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1140),
.B(n_812),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_989),
.Y(n_1281)
);

AOI221xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1130),
.A2(n_1056),
.B1(n_832),
.B2(n_1060),
.C(n_1140),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1121),
.A2(n_993),
.A3(n_1094),
.B(n_1119),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_989),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1008),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1121),
.A2(n_993),
.A3(n_1094),
.B(n_1119),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_1049),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1140),
.B(n_812),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1140),
.A2(n_812),
.B1(n_674),
.B2(n_639),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1089),
.A2(n_1123),
.B(n_1127),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_989),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_993),
.A2(n_1040),
.B(n_819),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1198),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1241),
.A2(n_1271),
.B1(n_1247),
.B2(n_1289),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1155),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1197),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1197),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1163),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1148),
.A2(n_1254),
.B1(n_1222),
.B2(n_1147),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1204),
.A2(n_1242),
.B1(n_1270),
.B2(n_1228),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1228),
.A2(n_1254),
.B1(n_1222),
.B2(n_1147),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1204),
.A2(n_1242),
.B1(n_1230),
.B2(n_1265),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1226),
.A2(n_1236),
.B1(n_1280),
.B2(n_1255),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1155),
.Y(n_1305)
);

INVx8_ASAP7_75t_L g1306 ( 
.A(n_1189),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1232),
.A2(n_1274),
.B1(n_1288),
.B2(n_1193),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1231),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1285),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1179),
.B(n_1146),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1187),
.A2(n_1182),
.B1(n_1195),
.B2(n_1193),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1188),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1272),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1202),
.Y(n_1314)
);

AO22x1_ASAP7_75t_L g1315 ( 
.A1(n_1189),
.A2(n_1164),
.B1(n_1275),
.B2(n_1287),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1269),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1141),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1181),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1259),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1227),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1178),
.A2(n_1200),
.B1(n_1151),
.B2(n_1275),
.Y(n_1321)
);

OAI22x1_ASAP7_75t_SL g1322 ( 
.A1(n_1141),
.A2(n_1240),
.B1(n_1246),
.B2(n_1238),
.Y(n_1322)
);

INVx4_ASAP7_75t_SL g1323 ( 
.A(n_1189),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1181),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1235),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1206),
.A2(n_1189),
.B1(n_1159),
.B2(n_1168),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1181),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1263),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1142),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1183),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1191),
.A2(n_1153),
.B1(n_1171),
.B2(n_1240),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1159),
.A2(n_1219),
.B1(n_1170),
.B2(n_1167),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1249),
.Y(n_1333)
);

AOI22x1_ASAP7_75t_SL g1334 ( 
.A1(n_1210),
.A2(n_1211),
.B1(n_1213),
.B2(n_1212),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1207),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1260),
.A2(n_1184),
.B1(n_1175),
.B2(n_1217),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1185),
.A2(n_1292),
.B1(n_1221),
.B2(n_1177),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1149),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1214),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1229),
.B1(n_1233),
.B2(n_1166),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1218),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1169),
.A2(n_1190),
.B1(n_1256),
.B2(n_1194),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_1229),
.B1(n_1233),
.B2(n_1166),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1220),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_1165),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1234),
.A2(n_1284),
.B1(n_1281),
.B2(n_1261),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1268),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1278),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1282),
.B(n_1199),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1218),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1145),
.A2(n_1205),
.B1(n_1174),
.B2(n_1157),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1215),
.Y(n_1352)
);

BUFx4f_ASAP7_75t_SL g1353 ( 
.A(n_1172),
.Y(n_1353)
);

BUFx8_ASAP7_75t_SL g1354 ( 
.A(n_1172),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1269),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1282),
.A2(n_1273),
.B(n_1162),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1266),
.A2(n_1201),
.B1(n_1267),
.B2(n_1152),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1160),
.A2(n_1208),
.B1(n_1291),
.B2(n_1293),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1192),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1173),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1208),
.A2(n_1158),
.B1(n_1253),
.B2(n_1192),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1192),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1253),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1150),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1150),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1223),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1216),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1176),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1158),
.A2(n_1273),
.B1(n_1250),
.B2(n_1209),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1225),
.A2(n_1244),
.B1(n_1243),
.B2(n_1277),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1237),
.A2(n_1276),
.B1(n_1258),
.B2(n_1186),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1209),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1224),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1144),
.A2(n_1161),
.B1(n_1180),
.B2(n_1279),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1245),
.A2(n_1290),
.B1(n_1264),
.B2(n_1262),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1224),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1154),
.A2(n_1286),
.B1(n_1239),
.B2(n_1257),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1154),
.A2(n_1286),
.B1(n_1239),
.B2(n_1257),
.Y(n_1378)
);

CKINVDCx6p67_ASAP7_75t_R g1379 ( 
.A(n_1251),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1154),
.A2(n_1286),
.B1(n_1257),
.B2(n_1283),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1283),
.A2(n_1148),
.B1(n_1138),
.B2(n_1241),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1203),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1143),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1203),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1228),
.A2(n_1138),
.B1(n_1148),
.B2(n_674),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1195),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1241),
.A2(n_1138),
.B1(n_674),
.B2(n_479),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1181),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1228),
.A2(n_1138),
.B1(n_1148),
.B2(n_674),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1241),
.A2(n_1138),
.B1(n_674),
.B2(n_479),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1241),
.A2(n_1138),
.B1(n_674),
.B2(n_479),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1181),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1198),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1272),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1147),
.A2(n_1228),
.B1(n_1222),
.B2(n_1254),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1198),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1231),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1156),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1141),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1231),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1241),
.B(n_1222),
.Y(n_1407)
);

OAI22x1_ASAP7_75t_L g1408 ( 
.A1(n_1222),
.A2(n_1254),
.B1(n_1147),
.B2(n_1193),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1226),
.B(n_1140),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1202),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1248),
.B(n_1252),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1197),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1197),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1155),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1148),
.A2(n_1138),
.B1(n_1241),
.B2(n_1222),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1156),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1164),
.B(n_1275),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1231),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1195),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1226),
.B(n_1140),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1198),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1294),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1371),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1397),
.A2(n_1295),
.B1(n_1300),
.B2(n_1302),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1373),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1376),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1395),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1351),
.A2(n_1422),
.B(n_1400),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1362),
.B(n_1359),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1403),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1400),
.A2(n_1422),
.B(n_1357),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1317),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1383),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1388),
.A2(n_1392),
.B1(n_1393),
.B2(n_1398),
.Y(n_1436)
);

NAND2x1_ASAP7_75t_L g1437 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1340),
.A2(n_1343),
.B(n_1367),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1323),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1407),
.B(n_1310),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1382),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1407),
.B(n_1310),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1366),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1331),
.A2(n_1337),
.B(n_1349),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1356),
.A2(n_1391),
.B(n_1386),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1369),
.Y(n_1447)
);

AO21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1381),
.A2(n_1404),
.B(n_1399),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1338),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1408),
.A2(n_1372),
.A3(n_1342),
.B(n_1346),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1366),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1307),
.B(n_1304),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.B(n_1344),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1364),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1379),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1385),
.A2(n_1406),
.B1(n_1390),
.B2(n_1412),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1379),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1306),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1372),
.B(n_1296),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1347),
.A2(n_1348),
.B(n_1384),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1323),
.B(n_1418),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1384),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1364),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1365),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1372),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1365),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1368),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1368),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1333),
.Y(n_1470)
);

NAND4xp25_ASAP7_75t_SL g1471 ( 
.A(n_1416),
.B(n_1303),
.C(n_1301),
.D(n_1332),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1380),
.B(n_1321),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1325),
.B(n_1411),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1299),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1312),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1326),
.A2(n_1402),
.B(n_1417),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1336),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1333),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1328),
.Y(n_1479)
);

CKINVDCx8_ASAP7_75t_R g1480 ( 
.A(n_1341),
.Y(n_1480)
);

BUFx8_ASAP7_75t_L g1481 ( 
.A(n_1387),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1298),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1328),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1370),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1305),
.A2(n_1316),
.B(n_1415),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1409),
.B(n_1421),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1315),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1323),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1335),
.A2(n_1339),
.B1(n_1352),
.B2(n_1308),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1334),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1339),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1413),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1345),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1413),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1352),
.B(n_1401),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1309),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1355),
.A2(n_1350),
.B(n_1414),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1425),
.A2(n_1453),
.B(n_1471),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1453),
.A2(n_1405),
.B(n_1419),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1311),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_SL g1501 ( 
.A1(n_1437),
.A2(n_1322),
.B(n_1313),
.C(n_1396),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1329),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1465),
.B(n_1355),
.Y(n_1503)
);

NAND2x1_ASAP7_75t_L g1504 ( 
.A(n_1445),
.B(n_1414),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1471),
.A2(n_1318),
.B(n_1297),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1436),
.A2(n_1297),
.B(n_1394),
.C(n_1389),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1437),
.B(n_1318),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1424),
.A2(n_1445),
.B(n_1433),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1433),
.A2(n_1430),
.B(n_1438),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1319),
.Y(n_1510)
);

AOI211xp5_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_1394),
.B(n_1389),
.C(n_1319),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1477),
.A2(n_1313),
.B1(n_1396),
.B2(n_1320),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1420),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1432),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1455),
.B(n_1467),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_SL g1516 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1449),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1449),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1434),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_SL g1521 ( 
.A(n_1461),
.B(n_1387),
.Y(n_1521)
);

AOI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1457),
.A2(n_1320),
.B1(n_1330),
.B2(n_1354),
.C(n_1353),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1456),
.B(n_1458),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1481),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1484),
.A2(n_1350),
.B(n_1327),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_SL g1526 ( 
.A1(n_1490),
.A2(n_1314),
.B(n_1410),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1496),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1430),
.A2(n_1324),
.B(n_1330),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1448),
.A2(n_1314),
.B1(n_1410),
.B2(n_1324),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1444),
.A2(n_1452),
.B(n_1484),
.C(n_1472),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1444),
.A2(n_1452),
.B(n_1472),
.C(n_1447),
.Y(n_1533)
);

AND2x6_ASAP7_75t_L g1534 ( 
.A(n_1459),
.B(n_1488),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1443),
.B(n_1454),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1479),
.Y(n_1536)
);

NAND4xp25_ASAP7_75t_L g1537 ( 
.A(n_1473),
.B(n_1490),
.C(n_1483),
.D(n_1454),
.Y(n_1537)
);

AOI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1456),
.A2(n_1458),
.B(n_1463),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1476),
.Y(n_1540)
);

A2O1A1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1468),
.A2(n_1469),
.B(n_1487),
.C(n_1448),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1431),
.B(n_1435),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_R g1543 ( 
.A(n_1470),
.B(n_1462),
.Y(n_1543)
);

AOI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1446),
.A2(n_1489),
.B1(n_1483),
.B2(n_1478),
.C(n_1487),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1426),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1427),
.A2(n_1423),
.B(n_1428),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1460),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1450),
.B(n_1474),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1446),
.B(n_1450),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1446),
.B(n_1474),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1550),
.B(n_1461),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1542),
.B(n_1442),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1550),
.B(n_1461),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1546),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1532),
.B(n_1480),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1540),
.B(n_1549),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1545),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1532),
.B(n_1463),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1549),
.B(n_1429),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1517),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1528),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1518),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1466),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1534),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1523),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1515),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1551),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1548),
.B(n_1442),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1537),
.B(n_1493),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1539),
.B(n_1451),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1534),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1538),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1555),
.A2(n_1533),
.B(n_1541),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1563),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1568),
.Y(n_1579)
);

INVx5_ASAP7_75t_L g1580 ( 
.A(n_1575),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1552),
.B(n_1530),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1557),
.B(n_1539),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1508),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1554),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1571),
.B(n_1530),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1571),
.B(n_1531),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1556),
.A2(n_1498),
.B(n_1544),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1554),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1554),
.B(n_1531),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1563),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1508),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1556),
.A2(n_1522),
.B(n_1529),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1595)
);

OAI33xp33_ASAP7_75t_L g1596 ( 
.A1(n_1562),
.A2(n_1500),
.A3(n_1519),
.B1(n_1527),
.B2(n_1512),
.B3(n_1510),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1575),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1508),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1563),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1568),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_SL g1601 ( 
.A(n_1570),
.B(n_1499),
.C(n_1511),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1570),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1575),
.B(n_1568),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1574),
.B(n_1509),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1566),
.B(n_1509),
.Y(n_1606)
);

BUFx4f_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1595),
.B(n_1574),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1584),
.B(n_1589),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1568),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1582),
.B(n_1553),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1578),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1580),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1589),
.B(n_1567),
.Y(n_1617)
);

AND2x4_ASAP7_75t_SL g1618 ( 
.A(n_1604),
.B(n_1547),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1578),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1606),
.B(n_1567),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1588),
.B(n_1575),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1588),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1578),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1593),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1600),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1577),
.A2(n_1524),
.B1(n_1560),
.B2(n_1470),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1567),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1579),
.B(n_1569),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1600),
.B(n_1569),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1606),
.B(n_1559),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1581),
.B(n_1558),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1582),
.B(n_1553),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1591),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1591),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1593),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1583),
.B(n_1572),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1593),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1599),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1631),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1627),
.A2(n_1587),
.B1(n_1601),
.B2(n_1596),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1623),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1633),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1608),
.B(n_1603),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1612),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1612),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1603),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1643),
.B(n_1580),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1626),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1620),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1624),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1618),
.A2(n_1594),
.B(n_1601),
.C(n_1573),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1633),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1580),
.Y(n_1664)
);

OAI322xp33_ASAP7_75t_L g1665 ( 
.A1(n_1627),
.A2(n_1583),
.A3(n_1605),
.B1(n_1573),
.B2(n_1585),
.C1(n_1586),
.C2(n_1596),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1624),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1626),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1609),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1609),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1622),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1622),
.B(n_1580),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1622),
.B(n_1615),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1618),
.B(n_1577),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1635),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1637),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1622),
.B(n_1580),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1637),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1622),
.B(n_1524),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1622),
.A2(n_1594),
.B1(n_1607),
.B2(n_1575),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1638),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1615),
.A2(n_1604),
.B(n_1597),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1610),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1636),
.B(n_1481),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1639),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1619),
.B(n_1605),
.Y(n_1689)
);

INVxp33_ASAP7_75t_L g1690 ( 
.A(n_1680),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1653),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1653),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1672),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1649),
.A2(n_1628),
.B(n_1621),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1648),
.B(n_1590),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1590),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1673),
.B(n_1609),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1655),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1673),
.B(n_1610),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1685),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1651),
.B(n_1642),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1661),
.B(n_1590),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1658),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1672),
.B(n_1674),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1687),
.Y(n_1710)
);

NAND2x1_ASAP7_75t_L g1711 ( 
.A(n_1672),
.B(n_1615),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1678),
.Y(n_1712)
);

INVx3_ASAP7_75t_SL g1713 ( 
.A(n_1674),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1642),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1613),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1669),
.B(n_1629),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1657),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1656),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1647),
.B(n_1629),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1663),
.B(n_1630),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1656),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1659),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1659),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1671),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1695),
.A2(n_1665),
.B1(n_1681),
.B2(n_1683),
.C(n_1674),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1702),
.B(n_1704),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1701),
.B(n_1713),
.Y(n_1728)
);

A2O1A1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1706),
.A2(n_1675),
.B(n_1664),
.C(n_1657),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1664),
.C(n_1675),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1690),
.A2(n_1580),
.B1(n_1607),
.B2(n_1604),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1707),
.B(n_1671),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1691),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1696),
.B(n_1662),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1700),
.A2(n_1501),
.B(n_1513),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1707),
.B(n_1668),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1501),
.C(n_1506),
.D(n_1505),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1708),
.A2(n_1525),
.B(n_1618),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1718),
.B(n_1630),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1691),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1693),
.A2(n_1577),
.B1(n_1607),
.B2(n_1580),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1692),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1711),
.A2(n_1577),
.B(n_1478),
.C(n_1506),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1713),
.A2(n_1693),
.B1(n_1697),
.B2(n_1543),
.Y(n_1744)
);

OAI31xp33_ASAP7_75t_L g1745 ( 
.A1(n_1708),
.A2(n_1600),
.A3(n_1628),
.B(n_1621),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1712),
.B(n_1613),
.Y(n_1746)
);

NOR4xp25_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1676),
.C(n_1688),
.D(n_1686),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1713),
.A2(n_1526),
.B(n_1491),
.C(n_1666),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1692),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1481),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1726),
.A2(n_1701),
.B1(n_1716),
.B2(n_1698),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1735),
.A2(n_1698),
.B(n_1716),
.Y(n_1753)
);

OAI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1735),
.A2(n_1577),
.B1(n_1576),
.B2(n_1725),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1709),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1728),
.B(n_1715),
.Y(n_1756)
);

AOI322xp5_ASAP7_75t_L g1757 ( 
.A1(n_1744),
.A2(n_1617),
.A3(n_1616),
.B1(n_1614),
.B2(n_1613),
.C1(n_1628),
.C2(n_1621),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1717),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1749),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1730),
.A2(n_1720),
.B1(n_1721),
.B2(n_1577),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1745),
.B(n_1747),
.C(n_1732),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1731),
.A2(n_1736),
.B1(n_1734),
.B2(n_1746),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1748),
.B(n_1481),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1749),
.B(n_1715),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1733),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1738),
.B(n_1703),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1729),
.A2(n_1699),
.B(n_1694),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1743),
.B(n_1699),
.C(n_1694),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1740),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1742),
.B(n_1705),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1750),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1759),
.B(n_1739),
.Y(n_1772)
);

XOR2xp5_ASAP7_75t_L g1773 ( 
.A(n_1761),
.B(n_1737),
.Y(n_1773)
);

AO22x1_ASAP7_75t_L g1774 ( 
.A1(n_1767),
.A2(n_1764),
.B1(n_1763),
.B2(n_1766),
.Y(n_1774)
);

OAI322xp33_ASAP7_75t_L g1775 ( 
.A1(n_1754),
.A2(n_1722),
.A3(n_1719),
.B1(n_1723),
.B2(n_1724),
.C1(n_1703),
.C2(n_1705),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1758),
.B(n_1719),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1755),
.B(n_1743),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1765),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1756),
.Y(n_1779)
);

XNOR2xp5_ASAP7_75t_L g1780 ( 
.A(n_1752),
.B(n_1495),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1771),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1770),
.Y(n_1782)
);

AO21x1_ASAP7_75t_L g1783 ( 
.A1(n_1754),
.A2(n_1723),
.B(n_1722),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1776),
.Y(n_1784)
);

NOR3xp33_ASAP7_75t_L g1785 ( 
.A(n_1774),
.B(n_1769),
.C(n_1753),
.Y(n_1785)
);

OAI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1773),
.A2(n_1777),
.B(n_1760),
.C(n_1772),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1780),
.B(n_1779),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1777),
.B(n_1768),
.C(n_1757),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1776),
.B(n_1762),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1782),
.A2(n_1769),
.B(n_1741),
.C(n_1724),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1775),
.A2(n_1714),
.B1(n_1676),
.B2(n_1660),
.C(n_1686),
.Y(n_1791)
);

OAI321xp33_ASAP7_75t_L g1792 ( 
.A1(n_1779),
.A2(n_1714),
.A3(n_1689),
.B1(n_1507),
.B2(n_1604),
.C(n_1597),
.Y(n_1792)
);

NOR4xp25_ASAP7_75t_L g1793 ( 
.A(n_1778),
.B(n_1688),
.C(n_1660),
.D(n_1684),
.Y(n_1793)
);

AOI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1788),
.A2(n_1783),
.B(n_1781),
.C(n_1689),
.Y(n_1794)
);

AOI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1786),
.A2(n_1495),
.B(n_1597),
.C(n_1614),
.Y(n_1795)
);

NAND4xp75_ASAP7_75t_L g1796 ( 
.A(n_1784),
.B(n_1614),
.C(n_1616),
.D(n_1617),
.Y(n_1796)
);

NAND5xp2_ASAP7_75t_L g1797 ( 
.A(n_1787),
.B(n_1785),
.C(n_1789),
.D(n_1792),
.E(n_1791),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_SL g1798 ( 
.A(n_1793),
.B(n_1480),
.C(n_1504),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1794),
.A2(n_1790),
.B1(n_1679),
.B2(n_1682),
.C(n_1677),
.Y(n_1799)
);

OAI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_1580),
.B(n_1667),
.C(n_1439),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1798),
.A2(n_1607),
.B(n_1617),
.C(n_1616),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1796),
.Y(n_1802)
);

NOR3xp33_ASAP7_75t_L g1803 ( 
.A(n_1797),
.B(n_1502),
.C(n_1503),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1796),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1802),
.B(n_1646),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1803),
.B(n_1625),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1502),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1801),
.B(n_1632),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1799),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_L g1810 ( 
.A(n_1809),
.B(n_1800),
.C(n_1580),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_SL g1811 ( 
.A1(n_1807),
.A2(n_1640),
.B(n_1625),
.C(n_1644),
.Y(n_1811)
);

AOI322xp5_ASAP7_75t_L g1812 ( 
.A1(n_1805),
.A2(n_1634),
.A3(n_1592),
.B1(n_1598),
.B2(n_1632),
.C1(n_1576),
.C2(n_1644),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1812),
.A2(n_1808),
.B1(n_1806),
.B2(n_1604),
.C(n_1605),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1806),
.B1(n_1810),
.B2(n_1811),
.Y(n_1814)
);

XOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1814),
.B(n_1482),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1814),
.B(n_1625),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1815),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1640),
.B1(n_1644),
.B2(n_1636),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1817),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1820),
.A2(n_1640),
.B1(n_1634),
.B2(n_1632),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1819),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1646),
.B1(n_1645),
.B2(n_1641),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_R g1824 ( 
.A1(n_1823),
.A2(n_1607),
.B1(n_1521),
.B2(n_1516),
.C(n_1604),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1494),
.B(n_1482),
.C(n_1492),
.Y(n_1825)
);


endmodule