module real_aes_6865_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g522 ( .A1(n_0), .A2(n_169), .B(n_523), .C(n_526), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_1), .B(n_518), .Y(n_527) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g167 ( .A(n_3), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_4), .B(n_170), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_5), .A2(n_487), .B(n_562), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_6), .A2(n_771), .B1(n_774), .B2(n_775), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_6), .Y(n_775) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_7), .A2(n_177), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_8), .A2(n_38), .B1(n_157), .B2(n_205), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_9), .B(n_177), .Y(n_185) );
AND2x6_ASAP7_75t_L g172 ( .A(n_10), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_11), .A2(n_172), .B(n_492), .C(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_12), .A2(n_42), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_12), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_13), .B(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_13), .B(n_39), .Y(n_467) );
INVx1_ASAP7_75t_L g151 ( .A(n_14), .Y(n_151) );
INVx1_ASAP7_75t_L g148 ( .A(n_15), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_16), .B(n_153), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_17), .B(n_170), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_18), .B(n_144), .Y(n_251) );
AO32x2_ASAP7_75t_L g221 ( .A1(n_19), .A2(n_143), .A3(n_177), .B1(n_196), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_20), .B(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_21), .B(n_144), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_22), .A2(n_58), .B1(n_157), .B2(n_205), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_23), .A2(n_85), .B1(n_153), .B2(n_157), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_24), .B(n_157), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_25), .A2(n_196), .B(n_492), .C(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_26), .A2(n_106), .B1(n_118), .B2(n_785), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_27), .A2(n_196), .B(n_492), .C(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_28), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_29), .B(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_30), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_30), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_31), .A2(n_487), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_32), .B(n_198), .Y(n_239) );
INVx2_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_34), .A2(n_490), .B(n_494), .C(n_500), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_35), .B(n_157), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_36), .B(n_198), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_37), .B(n_216), .Y(n_545) );
INVx1_ASAP7_75t_L g117 ( .A(n_39), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_40), .B(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_41), .Y(n_539) );
INVx1_ASAP7_75t_L g773 ( .A(n_42), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_43), .B(n_170), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_44), .A2(n_455), .B1(n_458), .B2(n_459), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_44), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_45), .B(n_487), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_46), .A2(n_48), .B1(n_456), .B2(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_46), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_46), .A2(n_131), .B1(n_132), .B2(n_457), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_47), .A2(n_490), .B(n_500), .C(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_48), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_49), .B(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g524 ( .A(n_50), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_51), .A2(n_94), .B1(n_205), .B2(n_206), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_52), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_53), .B(n_157), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_54), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g555 ( .A(n_55), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_56), .B(n_487), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_57), .B(n_165), .Y(n_184) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_59), .A2(n_63), .B1(n_153), .B2(n_157), .Y(n_249) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_60), .A2(n_70), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_60), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_61), .B(n_157), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_62), .B(n_157), .Y(n_213) );
INVx1_ASAP7_75t_L g173 ( .A(n_64), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_65), .B(n_487), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_66), .B(n_518), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_67), .A2(n_159), .B(n_165), .C(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_68), .B(n_157), .Y(n_168) );
INVx1_ASAP7_75t_L g147 ( .A(n_69), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_70), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_71), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_72), .B(n_170), .Y(n_498) );
AO32x2_ASAP7_75t_L g202 ( .A1(n_73), .A2(n_177), .A3(n_196), .B1(n_203), .B2(n_208), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_74), .B(n_171), .Y(n_536) );
INVx1_ASAP7_75t_L g192 ( .A(n_75), .Y(n_192) );
INVx1_ASAP7_75t_L g234 ( .A(n_76), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_77), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_78), .B(n_497), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_79), .A2(n_492), .B(n_500), .C(n_589), .Y(n_588) );
AOI222xp33_ASAP7_75t_L g472 ( .A1(n_80), .A2(n_473), .B1(n_766), .B2(n_767), .C1(n_776), .C2(n_780), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_81), .B(n_153), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_82), .Y(n_563) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_84), .B(n_496), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_86), .B(n_205), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_87), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_88), .B(n_153), .Y(n_238) );
INVx2_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_90), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_91), .B(n_195), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_92), .B(n_153), .Y(n_181) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_93), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g464 ( .A(n_93), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g477 ( .A(n_93), .B(n_466), .Y(n_477) );
INVx2_ASAP7_75t_L g765 ( .A(n_93), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_95), .A2(n_104), .B1(n_153), .B2(n_154), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_96), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_97), .Y(n_495) );
INVxp67_ASAP7_75t_L g566 ( .A(n_98), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_99), .B(n_153), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g532 ( .A(n_101), .Y(n_532) );
INVx1_ASAP7_75t_L g590 ( .A(n_102), .Y(n_590) );
AND2x2_ASAP7_75t_L g557 ( .A(n_103), .B(n_198), .Y(n_557) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx5_ASAP7_75t_SL g785 ( .A(n_108), .Y(n_785) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_115), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g466 ( .A(n_111), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_471), .Y(n_118) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g784 ( .A(n_122), .Y(n_784) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_461), .B(n_468), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_130), .B2(n_460), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_126), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_127), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_132), .B1(n_453), .B2(n_454), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_419), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_323), .C(n_407), .Y(n_133) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_266), .C(n_288), .D(n_304), .Y(n_134) );
AOI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_199), .B1(n_225), .B2(n_244), .C(n_252), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_175), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_138), .B(n_244), .Y(n_278) );
NAND4xp25_ASAP7_75t_L g318 ( .A(n_138), .B(n_306), .C(n_319), .D(n_321), .Y(n_318) );
INVxp67_ASAP7_75t_L g435 ( .A(n_138), .Y(n_435) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g317 ( .A(n_139), .B(n_255), .Y(n_317) );
AND2x2_ASAP7_75t_L g341 ( .A(n_139), .B(n_175), .Y(n_341) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g308 ( .A(n_140), .B(n_243), .Y(n_308) );
AND2x2_ASAP7_75t_L g348 ( .A(n_140), .B(n_329), .Y(n_348) );
AND2x2_ASAP7_75t_L g365 ( .A(n_140), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_140), .B(n_176), .Y(n_389) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g242 ( .A(n_141), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g260 ( .A(n_141), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g272 ( .A(n_141), .B(n_176), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_141), .B(n_186), .Y(n_294) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_149), .B(n_174), .Y(n_141) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_142), .A2(n_187), .B(n_197), .Y(n_186) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_143), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_145), .B(n_146), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_163), .B(n_172), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_159), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_152), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_152), .A2(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
INVx1_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
INVx3_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_157), .Y(n_592) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
AND2x6_ASAP7_75t_L g492 ( .A(n_158), .B(n_493), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_159), .A2(n_590), .B(n_591), .C(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_160), .A2(n_237), .B(n_238), .Y(n_236) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g497 ( .A(n_161), .Y(n_497) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
AND2x2_ASAP7_75t_L g488 ( .A(n_162), .B(n_166), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_162), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_168), .C(n_169), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_164), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_164), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_169), .A2(n_183), .B(n_184), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_169), .A2(n_195), .B1(n_223), .B2(n_224), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_169), .A2(n_195), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_170), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_170), .A2(n_189), .B(n_190), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_SL g232 ( .A1(n_170), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_170), .B(n_566), .Y(n_565) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_171), .A2(n_195), .B1(n_204), .B2(n_207), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_179), .B(n_182), .Y(n_178) );
BUFx3_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_172), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_232), .B(n_236), .Y(n_231) );
AND2x4_ASAP7_75t_L g487 ( .A(n_172), .B(n_488), .Y(n_487) );
INVx4_ASAP7_75t_SL g501 ( .A(n_172), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_172), .B(n_488), .Y(n_533) );
AND2x2_ASAP7_75t_L g275 ( .A(n_175), .B(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_175), .A2(n_325), .B1(n_328), .B2(n_330), .C(n_334), .Y(n_324) );
AND2x2_ASAP7_75t_L g383 ( .A(n_175), .B(n_348), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_175), .B(n_365), .Y(n_417) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_186), .Y(n_175) );
INVx3_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
AND2x2_ASAP7_75t_L g292 ( .A(n_176), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g346 ( .A(n_176), .B(n_261), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_176), .B(n_405), .Y(n_404) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_185), .Y(n_176) );
INVx4_ASAP7_75t_L g246 ( .A(n_177), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_177), .A2(n_542), .B(n_543), .Y(n_541) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_177), .Y(n_560) );
AND2x2_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
INVx1_ASAP7_75t_L g316 ( .A(n_186), .Y(n_316) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_186), .Y(n_322) );
AND2x2_ASAP7_75t_L g367 ( .A(n_186), .B(n_243), .Y(n_367) );
OR2x2_ASAP7_75t_L g406 ( .A(n_186), .B(n_245), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B(n_196), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx4_ASAP7_75t_L g525 ( .A(n_195), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_196), .B(n_246), .C(n_247), .Y(n_265) );
INVx2_ASAP7_75t_L g208 ( .A(n_198), .Y(n_208) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_198), .A2(n_211), .B(n_220), .Y(n_210) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_231), .B(n_239), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_198), .A2(n_486), .B(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g515 ( .A(n_198), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_198), .A2(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_199), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
AND2x2_ASAP7_75t_L g402 ( .A(n_200), .B(n_399), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_200), .B(n_384), .Y(n_434) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g333 ( .A(n_201), .B(n_257), .Y(n_333) );
AND2x2_ASAP7_75t_L g382 ( .A(n_201), .B(n_228), .Y(n_382) );
INVx1_ASAP7_75t_L g428 ( .A(n_201), .Y(n_428) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_202), .B(n_257), .Y(n_283) );
INVx1_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_202), .B(n_221), .Y(n_306) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_206), .Y(n_499) );
INVx2_ASAP7_75t_L g526 ( .A(n_206), .Y(n_526) );
INVx1_ASAP7_75t_L g513 ( .A(n_208), .Y(n_513) );
AND2x2_ASAP7_75t_L g374 ( .A(n_209), .B(n_282), .Y(n_374) );
INVx2_ASAP7_75t_L g439 ( .A(n_209), .Y(n_439) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AND2x2_ASAP7_75t_L g256 ( .A(n_210), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g269 ( .A(n_210), .B(n_229), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_210), .B(n_228), .Y(n_297) );
INVx1_ASAP7_75t_L g303 ( .A(n_210), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_210), .Y(n_320) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_210), .Y(n_332) );
INVx2_ASAP7_75t_L g400 ( .A(n_210), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
BUFx2_ASAP7_75t_L g354 ( .A(n_221), .Y(n_354) );
AND2x2_ASAP7_75t_L g399 ( .A(n_221), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_227), .B(n_336), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_227), .A2(n_398), .B(n_412), .Y(n_422) );
AND2x2_ASAP7_75t_L g447 ( .A(n_227), .B(n_333), .Y(n_447) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g369 ( .A(n_229), .Y(n_369) );
AND2x2_ASAP7_75t_L g398 ( .A(n_229), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_230), .Y(n_282) );
INVx2_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_230), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g255 ( .A(n_241), .Y(n_255) );
OR2x2_ASAP7_75t_L g268 ( .A(n_241), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g336 ( .A(n_241), .B(n_332), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_241), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g437 ( .A(n_241), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_241), .B(n_374), .Y(n_449) );
AND2x2_ASAP7_75t_L g328 ( .A(n_242), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g351 ( .A(n_242), .B(n_244), .Y(n_351) );
INVx2_ASAP7_75t_L g263 ( .A(n_243), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_243), .B(n_264), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_243), .B(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g286 ( .A(n_244), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g433 ( .A(n_244), .Y(n_433) );
AND2x2_ASAP7_75t_L g445 ( .A(n_244), .B(n_308), .Y(n_445) );
AND2x2_ASAP7_75t_L g271 ( .A(n_245), .B(n_261), .Y(n_271) );
INVx1_ASAP7_75t_L g366 ( .A(n_245), .Y(n_366) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_250), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_246), .B(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g518 ( .A(n_246), .Y(n_518) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_246), .A2(n_531), .B(n_538), .Y(n_530) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_246), .A2(n_587), .B(n_594), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_246), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_258), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_255), .B(n_302), .Y(n_311) );
OR2x2_ASAP7_75t_L g443 ( .A(n_255), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g360 ( .A(n_256), .B(n_301), .Y(n_360) );
AND2x2_ASAP7_75t_L g368 ( .A(n_256), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_256), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g451 ( .A(n_256), .B(n_298), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_257), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g438 ( .A(n_257), .B(n_301), .Y(n_438) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g290 ( .A(n_260), .B(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_L g452 ( .A(n_260), .Y(n_452) );
NOR2x1_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
AND2x2_ASAP7_75t_L g338 ( .A(n_263), .B(n_271), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_263), .B(n_406), .Y(n_432) );
INVx2_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
INVx3_ASAP7_75t_L g329 ( .A(n_264), .Y(n_329) );
OR2x2_ASAP7_75t_L g357 ( .A(n_264), .B(n_358), .Y(n_357) );
AOI311xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .A3(n_272), .B(n_273), .C(n_284), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_267), .A2(n_305), .B(n_307), .C(n_309), .Y(n_304) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g289 ( .A(n_269), .Y(n_289) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_271), .B(n_287), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_271), .B(n_272), .Y(n_440) );
AND2x2_ASAP7_75t_L g362 ( .A(n_272), .B(n_276), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_279), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g420 ( .A(n_276), .B(n_308), .Y(n_420) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AND2x2_ASAP7_75t_L g305 ( .A(n_281), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g350 ( .A(n_283), .Y(n_350) );
AND2x4_ASAP7_75t_L g412 ( .A(n_283), .B(n_381), .Y(n_412) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_286), .A2(n_352), .B1(n_364), .B2(n_368), .C1(n_370), .C2(n_374), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_292), .C(n_295), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_289), .B(n_333), .Y(n_356) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
OR2x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_378), .Y(n_377) );
OAI21xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .B(n_302), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_296), .B(n_314), .C(n_315), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_296), .A2(n_333), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_301), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g410 ( .A(n_301), .Y(n_410) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_301), .Y(n_426) );
INVx2_ASAP7_75t_L g384 ( .A(n_302), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_313), .B2(n_317), .C(n_318), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_312), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g446 ( .A(n_312), .Y(n_446) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g327 ( .A(n_319), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_319), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g385 ( .A(n_319), .B(n_333), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_319), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g418 ( .A(n_319), .B(n_353), .Y(n_418) );
BUFx3_ASAP7_75t_L g381 ( .A(n_320), .Y(n_381) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND5xp2_ASAP7_75t_L g323 ( .A(n_324), .B(n_342), .C(n_363), .D(n_375), .E(n_390), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_327), .A2(n_354), .A3(n_370), .B1(n_416), .B2(n_418), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_329), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g339 ( .A(n_333), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_349), .B1(n_351), .B2(n_352), .C(n_355), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g414 ( .A(n_346), .B(n_365), .Y(n_414) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_351), .A2(n_412), .B1(n_430), .B2(n_435), .C(n_436), .Y(n_429) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g373 ( .A(n_365), .Y(n_373) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_383), .B2(n_384), .C1(n_385), .C2(n_386), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B(n_403), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B(n_413), .C(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_423), .C(n_448), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_420), .Y(n_424) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_429), .C(n_441), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B(n_440), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B(n_452), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_455), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_464), .Y(n_470) );
NOR2x2_ASAP7_75t_L g782 ( .A(n_465), .B(n_765), .Y(n_782) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g764 ( .A(n_466), .B(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_468), .B(n_472), .C(n_783), .Y(n_471) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_475), .B1(n_478), .B2(n_764), .Y(n_473) );
INVx1_ASAP7_75t_L g777 ( .A(n_474), .Y(n_777) );
OAI22x1_ASAP7_75t_SL g776 ( .A1(n_475), .A2(n_479), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR3x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_678), .C(n_721), .Y(n_479) );
NAND5xp2_ASAP7_75t_L g480 ( .A(n_481), .B(n_605), .C(n_635), .D(n_652), .E(n_667), .Y(n_480) );
AOI221xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_528), .B1(n_568), .B2(n_574), .C(n_578), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_504), .Y(n_482) );
OR2x2_ASAP7_75t_L g583 ( .A(n_483), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g622 ( .A(n_483), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g640 ( .A(n_483), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_483), .B(n_576), .Y(n_657) );
OR2x2_ASAP7_75t_L g669 ( .A(n_483), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_483), .B(n_628), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_483), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_483), .B(n_606), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_483), .B(n_614), .Y(n_720) );
AND2x2_ASAP7_75t_L g752 ( .A(n_483), .B(n_516), .Y(n_752) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_483), .Y(n_760) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_484), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_484), .B(n_558), .Y(n_580) );
BUFx2_ASAP7_75t_L g602 ( .A(n_484), .Y(n_602) );
AND2x2_ASAP7_75t_L g631 ( .A(n_484), .B(n_505), .Y(n_631) );
AND2x2_ASAP7_75t_L g686 ( .A(n_484), .B(n_584), .Y(n_686) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_502), .Y(n_484) );
BUFx2_ASAP7_75t_L g508 ( .A(n_487), .Y(n_508) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_491), .A2(n_501), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_491), .A2(n_501), .B(n_563), .C(n_564), .Y(n_562) );
INVx5_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_498), .C(n_499), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_496), .A2(n_499), .B(n_555), .C(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_504), .B(n_640), .Y(n_649) );
OAI32xp33_ASAP7_75t_L g663 ( .A1(n_504), .A2(n_599), .A3(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_504), .B(n_665), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_504), .B(n_583), .Y(n_706) );
INVx1_ASAP7_75t_SL g735 ( .A(n_504), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g744 ( .A(n_504), .B(n_530), .C(n_686), .D(n_745), .Y(n_744) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
INVx5_ASAP7_75t_L g577 ( .A(n_505), .Y(n_577) );
AND2x2_ASAP7_75t_L g606 ( .A(n_505), .B(n_517), .Y(n_606) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_505), .Y(n_685) );
AND2x2_ASAP7_75t_L g755 ( .A(n_505), .B(n_702), .Y(n_755) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_509), .B(n_513), .Y(n_506) );
AND2x4_ASAP7_75t_L g628 ( .A(n_516), .B(n_577), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_516), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g662 ( .A(n_516), .B(n_584), .Y(n_662) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g614 ( .A(n_517), .B(n_586), .Y(n_614) );
AND2x2_ASAP7_75t_L g623 ( .A(n_517), .B(n_585), .Y(n_623) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_527), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g691 ( .A1(n_528), .A2(n_692), .B1(n_694), .B2(n_696), .C1(n_699), .C2(n_700), .Y(n_691) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_547), .Y(n_528) );
AND2x2_ASAP7_75t_L g624 ( .A(n_529), .B(n_625), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_529), .B(n_602), .C(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
INVx5_ASAP7_75t_SL g573 ( .A(n_530), .Y(n_573) );
OAI322xp33_ASAP7_75t_L g578 ( .A1(n_530), .A2(n_579), .A3(n_581), .B1(n_582), .B2(n_596), .C1(n_599), .C2(n_601), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_530), .B(n_571), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_530), .B(n_559), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
INVx2_ASAP7_75t_L g571 ( .A(n_540), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_540), .B(n_549), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_547), .B(n_609), .Y(n_664) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g643 ( .A(n_548), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_558), .Y(n_548) );
OR2x2_ASAP7_75t_L g572 ( .A(n_549), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_549), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g611 ( .A(n_549), .B(n_559), .Y(n_611) );
AND2x2_ASAP7_75t_L g634 ( .A(n_549), .B(n_571), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_549), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g650 ( .A(n_549), .B(n_609), .Y(n_650) );
AND2x2_ASAP7_75t_L g658 ( .A(n_549), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_549), .B(n_618), .Y(n_708) );
INVx5_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g598 ( .A(n_550), .B(n_573), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_550), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g625 ( .A(n_550), .B(n_559), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_550), .B(n_672), .Y(n_713) );
OR2x2_ASAP7_75t_L g729 ( .A(n_550), .B(n_673), .Y(n_729) );
AND2x2_ASAP7_75t_SL g736 ( .A(n_550), .B(n_690), .Y(n_736) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_550), .Y(n_743) );
OR2x6_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
AND2x2_ASAP7_75t_L g597 ( .A(n_558), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g647 ( .A(n_558), .B(n_571), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_558), .B(n_573), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_558), .B(n_609), .Y(n_731) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_559), .B(n_573), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_571), .Y(n_619) );
OR2x2_ASAP7_75t_L g673 ( .A(n_559), .B(n_571), .Y(n_673) );
AND2x2_ASAP7_75t_L g690 ( .A(n_559), .B(n_570), .Y(n_690) );
INVxp67_ASAP7_75t_L g712 ( .A(n_559), .Y(n_712) );
AND2x2_ASAP7_75t_L g739 ( .A(n_559), .B(n_609), .Y(n_739) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_559), .Y(n_746) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_567), .Y(n_559) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_570), .B(n_620), .Y(n_693) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g609 ( .A(n_571), .B(n_573), .Y(n_609) );
OR2x2_ASAP7_75t_L g676 ( .A(n_571), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g620 ( .A(n_572), .Y(n_620) );
OR2x2_ASAP7_75t_L g681 ( .A(n_572), .B(n_673), .Y(n_681) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g581 ( .A(n_576), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_576), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g582 ( .A(n_577), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_577), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_577), .B(n_584), .Y(n_616) );
INVx2_ASAP7_75t_L g661 ( .A(n_577), .Y(n_661) );
AND2x2_ASAP7_75t_L g674 ( .A(n_577), .B(n_614), .Y(n_674) );
AND2x2_ASAP7_75t_L g699 ( .A(n_577), .B(n_623), .Y(n_699) );
INVx1_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
INVx2_ASAP7_75t_SL g638 ( .A(n_583), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_584), .Y(n_641) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_585), .Y(n_604) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g702 ( .A(n_586), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .Y(n_587) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g671 ( .A(n_598), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_598), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_598), .A2(n_680), .B1(n_682), .B2(n_687), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_598), .B(n_690), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_599), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g633 ( .A(n_600), .Y(n_633) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OR2x2_ASAP7_75t_L g615 ( .A(n_602), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_602), .B(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g689 ( .A(n_602), .B(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_L g665 ( .A(n_604), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_612), .C(n_626), .Y(n_605) );
INVx1_ASAP7_75t_L g629 ( .A(n_606), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g737 ( .A1(n_606), .A2(n_738), .B1(n_740), .B2(n_741), .C(n_744), .Y(n_737) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g756 ( .A(n_609), .Y(n_756) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g705 ( .A(n_611), .B(n_644), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_617), .C(n_621), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OAI32xp33_ASAP7_75t_L g730 ( .A1(n_619), .A2(n_620), .A3(n_683), .B1(n_720), .B2(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g762 ( .A(n_622), .B(n_661), .Y(n_762) );
AND2x2_ASAP7_75t_L g709 ( .A(n_623), .B(n_661), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_623), .B(n_631), .Y(n_727) );
AOI31xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_629), .A3(n_630), .B(n_632), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_628), .B(n_640), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_628), .B(n_638), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_628), .A2(n_658), .B1(n_748), .B2(n_751), .C(n_753), .Y(n_747) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g653 ( .A(n_633), .B(n_654), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_642), .B1(n_645), .B2(n_648), .C1(n_650), .C2(n_651), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g718 ( .A(n_637), .Y(n_718) );
INVx1_ASAP7_75t_L g740 ( .A(n_640), .Y(n_740) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_643), .A2(n_754), .B1(n_756), .B2(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g659 ( .A(n_644), .Y(n_659) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_658), .B2(n_660), .C(n_663), .Y(n_652) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g697 ( .A(n_655), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g749 ( .A(n_655), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g724 ( .A(n_660), .Y(n_724) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g688 ( .A(n_661), .Y(n_688) );
INVx1_ASAP7_75t_L g670 ( .A(n_662), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_665), .B(n_752), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_674), .B2(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g761 ( .A(n_674), .Y(n_761) );
INVxp33_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_676), .B(n_720), .Y(n_719) );
OAI32xp33_ASAP7_75t_L g710 ( .A1(n_677), .A2(n_711), .A3(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_691), .C(n_703), .D(n_715), .Y(n_678) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_686), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx16_ASAP7_75t_R g696 ( .A(n_697), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_700), .A2(n_716), .B1(n_733), .B2(n_736), .C(n_737), .Y(n_732) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g751 ( .A(n_702), .B(n_752), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B1(n_707), .B2(n_709), .C(n_710), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_712), .B(n_743), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_722), .B(n_732), .C(n_747), .D(n_758), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .B(n_728), .C(n_730), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g763 ( .A(n_750), .Y(n_763) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B(n_763), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g779 ( .A(n_764), .Y(n_779) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
CKINVDCx14_ASAP7_75t_R g774 ( .A(n_771), .Y(n_774) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
endmodule