module fake_jpeg_97_n_205 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_205);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_76),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_0),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_60),
.B1(n_52),
.B2(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_58),
.B1(n_66),
.B2(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_64),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_59),
.C(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_56),
.B1(n_52),
.B2(n_48),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_56),
.B1(n_66),
.B2(n_72),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_64),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_63),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_65),
.B(n_55),
.C(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_50),
.B1(n_61),
.B2(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_61),
.B1(n_50),
.B2(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_67),
.B1(n_57),
.B2(n_2),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_90),
.B1(n_82),
.B2(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_67),
.B1(n_57),
.B2(n_2),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_67),
.B(n_1),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_111),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_127),
.B1(n_98),
.B2(n_15),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_5),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_12),
.B(n_14),
.C(n_15),
.D(n_16),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_7),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_30),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_100),
.B1(n_97),
.B2(n_108),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_17),
.B(n_18),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_20),
.C(n_21),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_147),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_116),
.B1(n_37),
.B2(n_38),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_33),
.B(n_34),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_36),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_141),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_134),
.Y(n_154)
);

AOI211xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_113),
.B(n_123),
.C(n_116),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_132),
.B1(n_142),
.B2(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_169),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_148),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_160),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_39),
.C(n_41),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_158),
.C(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_154),
.B1(n_151),
.B2(n_155),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_164),
.B1(n_170),
.B2(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_191),
.C(n_172),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_152),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_180),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_185),
.B(n_189),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_175),
.B(n_172),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_196),
.B(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_163),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_199),
.B1(n_167),
.B2(n_170),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_201),
.B(n_42),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_177),
.C(n_176),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_46),
.B(n_44),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_45),
.Y(n_205)
);


endmodule