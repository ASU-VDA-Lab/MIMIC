module fake_jpeg_19992_n_143 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_17),
.B1(n_19),
.B2(n_16),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_19),
.B1(n_10),
.B2(n_9),
.Y(n_37)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_41),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_26),
.B1(n_27),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_43),
.B1(n_45),
.B2(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_38),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_28),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_36),
.C(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_25),
.B1(n_22),
.B2(n_34),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_52),
.B1(n_65),
.B2(n_29),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_57),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_50),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_40),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_15),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_63),
.B(n_42),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_24),
.B(n_29),
.C(n_36),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_11),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_12),
.C(n_13),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_72),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_50),
.B(n_47),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_73),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_42),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_40),
.B1(n_24),
.B2(n_11),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_57),
.B1(n_62),
.B2(n_29),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_55),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_12),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_70),
.B1(n_79),
.B2(n_66),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_67),
.B(n_61),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_90),
.B1(n_93),
.B2(n_0),
.Y(n_105)
);

NOR4xp25_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_62),
.C(n_20),
.D(n_12),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_5),
.C(n_7),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_7),
.B1(n_9),
.B2(n_8),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_83),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_5),
.B1(n_7),
.B2(n_2),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_100),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_74),
.B(n_72),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_90),
.B(n_92),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_82),
.B1(n_81),
.B2(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_104),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_92),
.C(n_81),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_120),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_112),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_96),
.B(n_86),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_96),
.B(n_1),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_14),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_114),
.C(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_126),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_113),
.B1(n_107),
.B2(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_133),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_117),
.B(n_111),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_123),
.B(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_132),
.C(n_14),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_134),
.C(n_13),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_3),
.A3(n_4),
.B1(n_13),
.B2(n_14),
.C1(n_135),
.C2(n_136),
.Y(n_141)
);

XNOR2x2_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_3),
.Y(n_143)
);


endmodule