module real_jpeg_1258_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_70),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_55),
.B1(n_57),
.B2(n_70),
.Y(n_209)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_4),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_44),
.B1(n_66),
.B2(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_44),
.B1(n_55),
.B2(n_57),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_6),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_7),
.B(n_66),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_7),
.B(n_169),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_7),
.A2(n_32),
.B(n_33),
.C(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_7),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_7),
.B(n_38),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_219),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_7),
.B(n_52),
.C(n_55),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_7),
.B(n_96),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_7),
.B(n_85),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_128),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_55),
.B1(n_57),
.B2(n_128),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_9),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_106),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_9),
.A2(n_55),
.B1(n_57),
.B2(n_106),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_10),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_168),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_168),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_10),
.A2(n_55),
.B1(n_57),
.B2(n_168),
.Y(n_279)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_20),
.B(n_345),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g346 ( 
.A(n_14),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_15),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_15),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_16),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_16),
.A2(n_47),
.B1(n_66),
.B2(n_67),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_16),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_340),
.B(n_343),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_332),
.B(n_336),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_319),
.B(n_331),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_144),
.B(n_316),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_131),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_107),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_26),
.B(n_107),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_88),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_62),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_28),
.A2(n_29),
.B(n_48),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_62),
.C(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_48),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_30),
.A2(n_45),
.B1(n_46),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_30),
.A2(n_43),
.B1(n_45),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_30),
.A2(n_45),
.B1(n_82),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_30),
.A2(n_185),
.B(n_187),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_30),
.A2(n_187),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_31),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_31),
.A2(n_38),
.B1(n_186),
.B2(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_31),
.A2(n_38),
.B(n_323),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B(n_37),
.C(n_38),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_34),
.B1(n_74),
.B2(n_76),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_33),
.A2(n_67),
.A3(n_74),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_34),
.B(n_76),
.Y(n_191)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_38),
.B(n_165),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_39),
.A2(n_42),
.B(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_40),
.B(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_45),
.A2(n_124),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_45),
.A2(n_164),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_49),
.A2(n_54),
.B1(n_58),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_49),
.A2(n_54),
.B1(n_212),
.B2(n_246),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_49),
.A2(n_214),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_85),
.B1(n_101),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_50),
.A2(n_85),
.B1(n_122),
.B2(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_50),
.A2(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_50),
.B(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_54),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_54),
.A2(n_235),
.B(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_55),
.B(n_275),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_79),
.B2(n_87),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_64),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_80),
.C(n_84),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_64),
.B(n_135),
.C(n_142),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_73),
.B(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_76),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_67),
.A2(n_71),
.B(n_219),
.C(n_228),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_126),
.B(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_73),
.B1(n_78),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_72),
.A2(n_127),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_72),
.A2(n_169),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_72),
.A2(n_169),
.B1(n_326),
.B2(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_72),
.A2(n_169),
.B(n_334),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_73),
.A2(n_103),
.B(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_74),
.Y(n_76)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_84),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_84),
.B(n_136),
.C(n_140),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_85),
.B(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_102),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_90),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_102),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_91),
.A2(n_92),
.B1(n_99),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_97),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_93),
.A2(n_96),
.B1(n_119),
.B2(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_93),
.A2(n_219),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_94),
.A2(n_95),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_94),
.A2(n_95),
.B1(n_194),
.B2(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_94),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_94),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_94),
.A2(n_95),
.B1(n_250),
.B2(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_95),
.A2(n_209),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_95),
.B(n_223),
.Y(n_252)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_96),
.A2(n_222),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_99),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_114),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.C(n_125),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_116),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_125),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_130),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_131),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_143),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_132),
.B(n_143),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_137),
.Y(n_325)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_141),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_170),
.B(n_315),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_146),
.B(n_149),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.C(n_166),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_157),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_158),
.B(n_160),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_196),
.B(n_314),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_172),
.B(n_174),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_181),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_175),
.B(n_179),
.Y(n_299)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_181),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_188),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_182),
.B(n_184),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_188),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI31xp33_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_296),
.A3(n_306),
.B(n_311),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_240),
.B(n_295),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_224),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_199),
.B(n_224),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.C(n_216),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_200),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_205),
.C(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_210),
.B(n_216),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_220),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_236),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_237),
.C(n_239),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_226),
.B(n_231),
.C(n_232),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_290),
.B(n_294),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_259),
.B(n_289),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_253),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_249),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_271),
.B(n_288),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_282),
.B(n_287),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_277),
.B(n_281),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_285),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_310),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_330),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_330),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_329),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_324),
.B1(n_327),
.B2(n_328),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_322),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_327),
.C(n_329),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_333),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_338),
.B(n_342),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);


endmodule