module fake_jpeg_13607_n_572 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_572);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_572;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_73),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_65),
.B(n_74),
.Y(n_176)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_0),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_12),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_89),
.Y(n_169)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_99),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_94),
.B(n_108),
.Y(n_177)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_27),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_101),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_98),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_12),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_39),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_116),
.Y(n_157)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_105),
.Y(n_183)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_106),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_39),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_11),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_118),
.B(n_52),
.Y(n_181)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_123),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_40),
.B(n_2),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_45),
.B(n_32),
.C(n_46),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_145),
.A2(n_207),
.B(n_172),
.C(n_200),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_70),
.A2(n_44),
.B1(n_57),
.B2(n_43),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_147),
.A2(n_100),
.B1(n_124),
.B2(n_121),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_68),
.A2(n_26),
.B1(n_57),
.B2(n_42),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_154),
.A2(n_158),
.B1(n_192),
.B2(n_200),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_26),
.B1(n_44),
.B2(n_43),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_66),
.B(n_55),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_170),
.B(n_178),
.Y(n_223)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_80),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_90),
.B(n_50),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_174),
.B(n_179),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_96),
.B(n_50),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_46),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_48),
.Y(n_215)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_67),
.B(n_45),
.C(n_54),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_125),
.C(n_9),
.Y(n_250)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_63),
.A2(n_26),
.B1(n_57),
.B2(n_44),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_60),
.Y(n_193)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_92),
.B(n_54),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_196),
.B(n_198),
.Y(n_283)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_197),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_92),
.B(n_52),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_61),
.A2(n_43),
.B1(n_51),
.B2(n_56),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_79),
.A2(n_51),
.B1(n_48),
.B2(n_5),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_202),
.A2(n_208),
.B1(n_85),
.B2(n_112),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_89),
.B(n_51),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_98),
.Y(n_237)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_77),
.A2(n_48),
.B1(n_51),
.B2(n_5),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_78),
.B(n_51),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_107),
.Y(n_214)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_212),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_214),
.B(n_250),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_215),
.B(n_264),
.Y(n_300)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_218),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_145),
.A2(n_2),
.B(n_3),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_220),
.A2(n_237),
.B(n_249),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_222),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_227),
.B(n_233),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_128),
.B(n_2),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_138),
.B(n_2),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_140),
.B(n_3),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_236),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_156),
.B(n_59),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_59),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_234),
.B(n_240),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_5),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_238),
.A2(n_242),
.B1(n_269),
.B2(n_279),
.Y(n_323)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_239),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_5),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_149),
.A2(n_84),
.B1(n_111),
.B2(n_102),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_251),
.Y(n_303)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_248),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_135),
.A2(n_141),
.B(n_172),
.C(n_173),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_6),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_131),
.B(n_6),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_258),
.C(n_260),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_148),
.B(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_195),
.B(n_9),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_256),
.B(n_273),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_139),
.B(n_9),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_259),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_180),
.B(n_10),
.Y(n_260)
);

OR2x2_ASAP7_75t_SL g261 ( 
.A(n_149),
.B(n_10),
.Y(n_261)
);

OR2x4_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_274),
.Y(n_299)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_262),
.Y(n_338)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_127),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_271),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_161),
.B(n_10),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_168),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_153),
.B(n_10),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_165),
.A2(n_162),
.B1(n_142),
.B2(n_199),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_147),
.A2(n_11),
.B1(n_188),
.B2(n_175),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_280),
.B1(n_162),
.B2(n_132),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_133),
.B(n_206),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_164),
.B(n_199),
.Y(n_273)
);

OR2x2_ASAP7_75t_SL g274 ( 
.A(n_207),
.B(n_202),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_164),
.B(n_184),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_276),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_183),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_192),
.A2(n_158),
.B1(n_154),
.B2(n_129),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_130),
.A2(n_132),
.B1(n_166),
.B2(n_129),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_183),
.B(n_206),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_211),
.C(n_212),
.Y(n_305)
);

OR2x2_ASAP7_75t_SL g282 ( 
.A(n_134),
.B(n_155),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_211),
.B(n_144),
.C(n_151),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_285),
.A2(n_292),
.B1(n_293),
.B2(n_304),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_263),
.B(n_229),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_289),
.B(n_308),
.Y(n_379)
);

AO21x1_ASAP7_75t_SL g349 ( 
.A1(n_291),
.A2(n_333),
.B(n_213),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_214),
.A2(n_130),
.B1(n_134),
.B2(n_152),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_152),
.B1(n_155),
.B2(n_166),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_235),
.A2(n_184),
.B1(n_203),
.B2(n_144),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_248),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_230),
.B(n_211),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_276),
.A2(n_250),
.B1(n_238),
.B2(n_236),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_309),
.A2(n_312),
.B1(n_313),
.B2(n_316),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_245),
.A2(n_256),
.B1(n_251),
.B2(n_274),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_273),
.A2(n_275),
.B1(n_231),
.B2(n_223),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_220),
.A2(n_283),
.B1(n_282),
.B2(n_228),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_257),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_317),
.B(n_318),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_261),
.B(n_249),
.CI(n_260),
.CON(n_318),
.SN(n_318)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_325),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_232),
.B(n_219),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_260),
.A2(n_252),
.B(n_258),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_258),
.B(n_265),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_264),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_330),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_281),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g333 ( 
.A1(n_262),
.A2(n_246),
.B1(n_217),
.B2(n_218),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_252),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_222),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_221),
.B(n_237),
.C(n_224),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_237),
.C(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_354),
.C(n_377),
.Y(n_412)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

AO21x2_ASAP7_75t_L g343 ( 
.A1(n_326),
.A2(n_247),
.B(n_244),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_343),
.A2(n_364),
.B1(n_368),
.B2(n_376),
.Y(n_409)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_358),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_326),
.A2(n_239),
.B(n_241),
.Y(n_347)
);

INVx3_ASAP7_75t_SL g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_300),
.B(n_319),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_335),
.Y(n_388)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_355),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_216),
.C(n_271),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_322),
.B(n_216),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_360),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_311),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_369),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_309),
.A2(n_312),
.B1(n_293),
.B2(n_304),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_323),
.A2(n_254),
.B1(n_259),
.B2(n_225),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_367),
.B1(n_372),
.B2(n_284),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_366),
.B(n_375),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_323),
.A2(n_322),
.B1(n_334),
.B2(n_286),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_286),
.A2(n_222),
.B1(n_226),
.B2(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_371),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_329),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_303),
.A2(n_226),
.B1(n_330),
.B2(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_374),
.Y(n_406)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_315),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_291),
.A2(n_292),
.B1(n_306),
.B2(n_288),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_297),
.B(n_296),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_313),
.A2(n_285),
.B1(n_303),
.B2(n_296),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_380),
.B1(n_290),
.B2(n_288),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_299),
.A2(n_305),
.B1(n_318),
.B2(n_284),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_382),
.A2(n_395),
.B1(n_398),
.B2(n_404),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_362),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_391),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_415),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_357),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_355),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_408),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_364),
.A2(n_299),
.B1(n_327),
.B2(n_308),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_396),
.A2(n_410),
.B1(n_356),
.B2(n_343),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_289),
.B(n_287),
.C(n_300),
.D(n_298),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_397),
.A2(n_405),
.B(n_371),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_361),
.A2(n_287),
.B1(n_301),
.B2(n_307),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_306),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_401),
.C(n_407),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_307),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_336),
.B1(n_294),
.B2(n_320),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_367),
.B(n_332),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_331),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_345),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_365),
.A2(n_336),
.B1(n_294),
.B2(n_320),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_332),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_340),
.C(n_354),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_416),
.Y(n_463)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_406),
.Y(n_417)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_417),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_406),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_419),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_385),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_409),
.A2(n_344),
.B1(n_341),
.B2(n_339),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_420),
.A2(n_431),
.B1(n_440),
.B2(n_446),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_385),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_426),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_405),
.A2(n_349),
.B(n_356),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_384),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_392),
.Y(n_427)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_432),
.C(n_438),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_436),
.B1(n_422),
.B2(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_383),
.A2(n_347),
.B1(n_346),
.B2(n_350),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_412),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_384),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_439),
.Y(n_455)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_396),
.A2(n_378),
.B1(n_343),
.B2(n_371),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_350),
.C(n_347),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_381),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_383),
.A2(n_343),
.B1(n_352),
.B2(n_363),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_352),
.B(n_360),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_399),
.B(n_397),
.Y(n_473)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_386),
.Y(n_445)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_445),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_353),
.B1(n_351),
.B2(n_348),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_448),
.A2(n_450),
.B1(n_453),
.B2(n_469),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_382),
.B1(n_389),
.B2(n_405),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_432),
.B(n_401),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_451),
.B(n_434),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_402),
.B1(n_403),
.B2(n_395),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_435),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_454),
.B(n_449),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_390),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_456),
.B(n_468),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_388),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_458),
.C(n_467),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_407),
.C(n_413),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_425),
.A2(n_402),
.B1(n_410),
.B2(n_393),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_465),
.A2(n_417),
.B1(n_419),
.B2(n_421),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_393),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_398),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_424),
.A2(n_402),
.B1(n_404),
.B2(n_411),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_416),
.B(n_444),
.Y(n_485)
);

XNOR2x1_ASAP7_75t_L g510 ( 
.A(n_476),
.B(n_498),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_439),
.Y(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_424),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_431),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_482),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_428),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_433),
.Y(n_483)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_418),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_463),
.B(n_470),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_489),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_447),
.B(n_445),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_494),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_420),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_420),
.C(n_437),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_493),
.C(n_451),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_411),
.C(n_446),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_441),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_497),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_496),
.B(n_453),
.Y(n_511)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_466),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_475),
.A2(n_463),
.B1(n_470),
.B2(n_465),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_499),
.A2(n_512),
.B1(n_476),
.B2(n_478),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_511),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_486),
.A2(n_485),
.B(n_489),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_477),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_475),
.A2(n_447),
.B1(n_462),
.B2(n_474),
.Y(n_512)
);

AO22x1_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_466),
.B1(n_448),
.B2(n_450),
.Y(n_514)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_514),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_460),
.C(n_474),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_460),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_477),
.C(n_492),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_518),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_487),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_519),
.A2(n_514),
.B1(n_504),
.B2(n_511),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_521),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_491),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_500),
.A2(n_498),
.B(n_484),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_510),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_479),
.C(n_496),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_526),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_484),
.C(n_494),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_527),
.A2(n_529),
.B(n_430),
.Y(n_542)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_503),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_374),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_427),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_531),
.A2(n_501),
.B1(n_499),
.B2(n_505),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_534),
.A2(n_522),
.B1(n_523),
.B2(n_530),
.Y(n_545)
);

OAI31xp67_ASAP7_75t_L g536 ( 
.A1(n_523),
.A2(n_514),
.A3(n_500),
.B(n_510),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_522),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_506),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_541),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_520),
.B(n_515),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_540),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_515),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_517),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_543),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_545),
.B(n_548),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_551),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_535),
.A2(n_525),
.B(n_472),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_550),
.A2(n_553),
.B(n_532),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_472),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_373),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_552),
.B(n_537),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_443),
.C(n_369),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_555),
.B(n_558),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_547),
.A2(n_544),
.B1(n_553),
.B2(n_536),
.Y(n_558)
);

A2O1A1O1Ixp25_ASAP7_75t_L g559 ( 
.A1(n_548),
.A2(n_543),
.B(n_541),
.C(n_443),
.D(n_359),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_559),
.B(n_560),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_370),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_546),
.C(n_358),
.Y(n_563)
);

A2O1A1O1Ixp25_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_565),
.B(n_556),
.C(n_564),
.D(n_561),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_290),
.C(n_314),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_562),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_566),
.B(n_567),
.C(n_568),
.Y(n_569)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_562),
.A2(n_337),
.B(n_314),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_320),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_570),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_337),
.Y(n_572)
);


endmodule