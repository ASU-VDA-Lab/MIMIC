module fake_jpeg_29053_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_60),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_21),
.B(n_36),
.C(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_41),
.B1(n_40),
.B2(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_5),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_66),
.B1(n_63),
.B2(n_47),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_15),
.B1(n_16),
.B2(n_22),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_18),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.C(n_29),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_65),
.C(n_68),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_6),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_32),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_93),
.C(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_30),
.B(n_31),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_34),
.B(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_89),
.B1(n_98),
.B2(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_103),
.CI(n_98),
.CON(n_108),
.SN(n_108)
);


endmodule