module fake_jpeg_12454_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_10),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_1),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_76),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_65),
.C(n_74),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_60),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_104),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_69),
.B1(n_62),
.B2(n_58),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_88),
.B1(n_86),
.B2(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_68),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_71),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_79),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_125),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_69),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_28),
.C(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_60),
.B1(n_77),
.B2(n_63),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_77),
.B1(n_52),
.B2(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_66),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_52),
.B1(n_51),
.B2(n_4),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_13),
.B(n_14),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_6),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_142),
.C(n_29),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_122),
.C(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_131),
.C(n_30),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_133),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_27),
.C(n_42),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_7),
.B(n_9),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_136),
.B(n_32),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_15),
.C(n_16),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_19),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_22),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_20),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_128),
.B(n_144),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_174),
.B(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_162),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_151),
.B1(n_153),
.B2(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_167),
.C(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_177),
.C(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_186),
.C(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_183),
.C(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_159),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_180),
.C(n_163),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_23),
.B(n_33),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_35),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_37),
.Y(n_195)
);


endmodule