module fake_jpeg_6718_n_323 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_64),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_44),
.B1(n_37),
.B2(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_32),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_44),
.B1(n_37),
.B2(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_44),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_57),
.B1(n_64),
.B2(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_70),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_19),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_25),
.B(n_28),
.C(n_31),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_35),
.B1(n_63),
.B2(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_91),
.B1(n_21),
.B2(n_34),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_94),
.B1(n_90),
.B2(n_75),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_40),
.A3(n_24),
.B1(n_21),
.B2(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_89),
.B1(n_48),
.B2(n_42),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_17),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_20),
.B(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_44),
.B1(n_37),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_35),
.B1(n_40),
.B2(n_37),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_17),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_119),
.B1(n_80),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_110),
.B1(n_116),
.B2(n_70),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_R g124 ( 
.A(n_101),
.B(n_86),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_31),
.B(n_25),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_109),
.B(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_98),
.B(n_116),
.C(n_91),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_42),
.B1(n_18),
.B2(n_20),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_46),
.B1(n_39),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_86),
.B1(n_73),
.B2(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_46),
.B1(n_34),
.B2(n_41),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_69),
.B1(n_23),
.B2(n_27),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_46),
.B1(n_41),
.B2(n_39),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_81),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_138),
.B1(n_150),
.B2(n_121),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_124),
.A2(n_25),
.B(n_31),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_89),
.C(n_67),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_126),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_139),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_89),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_89),
.B(n_87),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_143),
.B(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_67),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_141),
.B1(n_95),
.B2(n_102),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_78),
.C(n_55),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_106),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_28),
.B(n_25),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_60),
.B1(n_39),
.B2(n_41),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_151),
.B1(n_93),
.B2(n_27),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_39),
.B(n_41),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_60),
.B1(n_39),
.B2(n_69),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_55),
.A3(n_47),
.B1(n_25),
.B2(n_23),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_120),
.B(n_99),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_156),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_104),
.B(n_119),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_172),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_96),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_170),
.B1(n_182),
.B2(n_148),
.Y(n_186)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_118),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_31),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_176),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_99),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_180),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_125),
.A2(n_95),
.B(n_102),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_178),
.B1(n_138),
.B2(n_150),
.Y(n_193)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_55),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_149),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_27),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_47),
.B(n_31),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_186),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_135),
.B(n_126),
.C(n_143),
.D(n_129),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_207),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_200),
.B1(n_178),
.B2(n_161),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_135),
.C(n_145),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_202),
.C(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_149),
.B1(n_93),
.B2(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_23),
.B1(n_47),
.B2(n_22),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_206),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_0),
.C(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_0),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_237),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_214),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_157),
.C(n_156),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_224),
.C(n_230),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_188),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_184),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_154),
.C(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_154),
.B(n_183),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_189),
.B(n_2),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_155),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_182),
.B1(n_160),
.B2(n_168),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_229),
.A2(n_232),
.B1(n_231),
.B2(n_230),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_160),
.C(n_1),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_8),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_16),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_191),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_203),
.B1(n_197),
.B2(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_197),
.B1(n_211),
.B2(n_206),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_188),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_199),
.C(n_193),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_250),
.C(n_221),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_212),
.C(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_3),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_232),
.B1(n_2),
.B2(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_2),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_219),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_215),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_225),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_268),
.C(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_214),
.C(n_234),
.Y(n_268)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_243),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_272),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_265),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_284),
.B(n_6),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_256),
.B1(n_249),
.B2(n_240),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_250),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_260),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_253),
.B(n_257),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_266),
.B(n_259),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_3),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_287),
.B(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_261),
.C(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_280),
.B(n_12),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_239),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_16),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_6),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_11),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_278),
.B1(n_279),
.B2(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_291),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_309),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_290),
.B(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_300),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_313),
.B(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_316),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_292),
.B(n_298),
.Y(n_313)
);

NAND4xp25_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_311),
.A2(n_13),
.B(n_15),
.C(n_315),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_317),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_15),
.Y(n_323)
);


endmodule