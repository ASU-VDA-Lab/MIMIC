module fake_jpeg_23081_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_7),
.B1(n_11),
.B2(n_15),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_16),
.A2(n_18),
.B1(n_0),
.B2(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_21),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_14),
.B(n_0),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_35),
.C(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_23),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_3),
.C(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_17),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_28),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_22),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_26),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_41),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_44),
.B1(n_42),
.B2(n_32),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_46),
.B(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_33),
.C(n_44),
.Y(n_50)
);


endmodule