module real_jpeg_32810_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_592, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_592;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_120;
wire n_155;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_0),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_0),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_0),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_0),
.B(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_0),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_0),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_0),
.B(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_1),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_1),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_1),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_2),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_2),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_2),
.B(n_370),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_2),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_2),
.B(n_410),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g590 ( 
.A(n_4),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_5),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_5),
.B(n_178),
.Y(n_177)
);

NAND2x1_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_146),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_5),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_5),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_5),
.B(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_5),
.Y(n_352)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_5),
.B(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_6),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_7),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_49),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_7),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_7),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_7),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_7),
.B(n_263),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_9),
.Y(n_220)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_9),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_10),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_10),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_10),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_10),
.B(n_406),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_11),
.Y(n_181)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_11),
.Y(n_374)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_13),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_13),
.B(n_143),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_13),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_13),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_13),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_13),
.B(n_56),
.Y(n_504)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_14),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_16),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_16),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_16),
.B(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_16),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_16),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_16),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_70),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_17),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_17),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_17),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_17),
.B(n_511),
.Y(n_510)
);

OAI311xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_121),
.A3(n_578),
.B1(n_583),
.C1(n_589),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

AOI322xp5_ASAP7_75t_L g589 ( 
.A1(n_20),
.A2(n_578),
.A3(n_585),
.B1(n_586),
.B2(n_587),
.C1(n_588),
.C2(n_590),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_21),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_23),
.B(n_586),
.Y(n_585)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_77),
.B(n_120),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_24),
.B(n_77),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_27),
.A2(n_28),
.B1(n_111),
.B2(n_176),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_28),
.B(n_68),
.C(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_31),
.Y(n_295)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_35),
.A2(n_36),
.B1(n_471),
.B2(n_475),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_35),
.A2(n_36),
.B1(n_489),
.B2(n_490),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_35),
.B(n_490),
.C(n_493),
.Y(n_543)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_36),
.B(n_475),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_36),
.B(n_475),
.Y(n_497)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_47),
.C(n_53),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2x2_ASAP7_75t_SL g289 ( 
.A(n_41),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_41),
.B(n_296),
.C(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_45),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_47),
.B(n_298),
.C(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_48),
.B(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_51),
.Y(n_308)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_52),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_52),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_68),
.C(n_73),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_53),
.A2(n_54),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_68),
.B1(n_69),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_55),
.B(n_131),
.C(n_243),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_57),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_58),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_58),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.C(n_67),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_66),
.Y(n_512)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_68),
.A2(n_69),
.B1(n_550),
.B2(n_551),
.Y(n_549)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_69),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_69),
.B(n_213),
.C(n_217),
.Y(n_251)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_72),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22x1_ASAP7_75t_L g456 ( 
.A1(n_74),
.A2(n_75),
.B1(n_135),
.B2(n_136),
.Y(n_456)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_75),
.B(n_134),
.C(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_115),
.C(n_117),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_78),
.B(n_115),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.C(n_97),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_79),
.B(n_82),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_93),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_84),
.B(n_284),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_87),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g469 ( 
.A(n_87),
.B(n_197),
.C(n_287),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_93),
.B(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_97),
.A2(n_98),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_108),
.C(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_111),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_111),
.A2(n_176),
.B1(n_508),
.B2(n_513),
.Y(n_507)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_117),
.B(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_122),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_532),
.B(n_575),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_524),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_317),
.C(n_436),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_271),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_221),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_127),
.B(n_221),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_169),
.C(n_204),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_128),
.B(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_148),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_129),
.B(n_154),
.C(n_167),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.C(n_144),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_130),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_131),
.A2(n_242),
.B1(n_243),
.B2(n_246),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_131),
.Y(n_246)
);

AO22x1_ASAP7_75t_SL g336 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_246),
.Y(n_336)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_133),
.Y(n_288)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_133),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_134),
.A2(n_135),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_134),
.B(n_176),
.C(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_325)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_154),
.B1(n_167),
.B2(n_168),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_152),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_153),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_153),
.B(n_232),
.C(n_238),
.Y(n_302)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_165),
.C(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_161),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_161),
.B(n_441),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_161),
.B(n_443),
.C(n_494),
.Y(n_493)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_163),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_163),
.Y(n_335)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_163),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_164),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_169),
.B(n_205),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.C(n_194),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_170),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_182),
.A2(n_194),
.B1(n_195),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_182),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_191),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_183),
.B(n_191),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2x2_ASAP7_75t_SL g423 ( 
.A(n_187),
.B(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_200),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_196),
.A2(n_197),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_224),
.C(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx8_ASAP7_75t_L g492 ( 
.A(n_216),
.Y(n_492)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_220),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_220),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_247),
.Y(n_221)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_239),
.Y(n_226)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_245),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_269),
.B2(n_270),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_252),
.C(n_255),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_267),
.C(n_298),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_260),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_262),
.A2(n_268),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_265),
.Y(n_455)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_271),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_272),
.B(n_275),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.Y(n_275)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_276),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_299),
.B1(n_300),
.B2(n_313),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_297),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_283),
.B(n_289),
.C(n_316),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_328),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_286),
.A2(n_287),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_328),
.Y(n_366)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_287),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_297),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_290)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_294),
.Y(n_449)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_300),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

HB1xp67_ASAP7_75t_SL g460 ( 
.A(n_302),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_303),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_311),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_309),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_310),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_311),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_312),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_313),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_339),
.B(n_435),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_337),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_319),
.B(n_337),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.C(n_326),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_320),
.B(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_336),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_331),
.A2(n_332),
.B1(n_336),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_429),
.B(n_434),
.Y(n_339)
);

OAI21x1_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_417),
.B(n_428),
.Y(n_340)
);

AOI21x1_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_387),
.B(n_416),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_361),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_361),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_355),
.C(n_358),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_344),
.A2(n_345),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_351),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_355),
.A2(n_358),
.B1(n_359),
.B2(n_397),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_355),
.Y(n_397)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_367),
.B1(n_385),
.B2(n_386),
.Y(n_361)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_366),
.C(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_367),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_375),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_376),
.C(n_380),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_398),
.B(n_415),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_394),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_404),
.B(n_414),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_401),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_409),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx12f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_420),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_423),
.C(n_425),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_SL g434 ( 
.A(n_430),
.B(n_433),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_436),
.A2(n_525),
.B(n_528),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_480),
.B1(n_515),
.B2(n_520),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_437),
.B(n_480),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_480),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_457),
.C(n_462),
.Y(n_437)
);

XNOR2x1_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_458),
.Y(n_523)
);

XOR2x2_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_447),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_448),
.C(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

MAJx2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_458)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_462),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_462)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_477),
.C(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.C(n_467),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_469),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_473),
.Y(n_476)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_572),
.C(n_574),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_485),
.B1(n_499),
.B2(n_514),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_498),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_495),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_493),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_495),
.B(n_546),
.C(n_547),
.Y(n_545)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_498),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_499),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_507),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_505),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_501),
.Y(n_539)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_504),
.Y(n_554)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_538),
.C(n_539),
.Y(n_537)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_508),
.Y(n_513)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_521),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.C(n_519),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_521),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_566),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_533),
.A2(n_576),
.B(n_577),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_558),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_534),
.B(n_558),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_535),
.A2(n_544),
.B1(n_545),
.B2(n_556),
.Y(n_534)
);

INVxp33_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_557),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_540),
.Y(n_536)
);

MAJx2_ASAP7_75t_L g565 ( 
.A(n_537),
.B(n_541),
.C(n_543),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_548),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_545),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_545),
.Y(n_568)
);

OAI33xp33_ASAP7_75t_L g576 ( 
.A1(n_545),
.A2(n_568),
.A3(n_569),
.B1(n_570),
.B2(n_571),
.B3(n_592),
.Y(n_576)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_548),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_552),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_553),
.C(n_555),
.Y(n_561)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_555),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_557),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_559),
.B(n_565),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_562),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_565),
.C(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_562),
.Y(n_580)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_563),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_571),
.Y(n_566)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_569),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_581),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_581),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_585),
.C(n_587),
.Y(n_583)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);


endmodule