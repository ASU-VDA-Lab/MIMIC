module fake_jpeg_25966_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_6),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_39),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_32),
.C(n_30),
.Y(n_62)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_17),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_47),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_50),
.C(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_59),
.B1(n_73),
.B2(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_38),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_46),
.B1(n_11),
.B2(n_14),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_37),
.B(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_22),
.B1(n_28),
.B2(n_23),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_93),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_81),
.B(n_92),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_90),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_46),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_85),
.B1(n_52),
.B2(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_53),
.B(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_97),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_72),
.B1(n_52),
.B2(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_104),
.B1(n_109),
.B2(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_75),
.B(n_84),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_63),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_77),
.B1(n_95),
.B2(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_48),
.B1(n_89),
.B2(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_117),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_64),
.C(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_92),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_76),
.B(n_49),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_131),
.B(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_89),
.B1(n_96),
.B2(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_104),
.B1(n_113),
.B2(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_109),
.B1(n_121),
.B2(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_48),
.B(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_139),
.B1(n_143),
.B2(n_126),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_115),
.C(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_137),
.C(n_138),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_119),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_144),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_110),
.B1(n_102),
.B2(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_108),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_142),
.C(n_138),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_120),
.C(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_134),
.B(n_133),
.Y(n_153)
);

XNOR2x2_ASAP7_75t_SL g154 ( 
.A(n_145),
.B(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_140),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_126),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_162),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_166),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_164),
.B(n_161),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_150),
.B(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_161),
.Y(n_170)
);

AND3x1_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_171),
.C(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_141),
.Y(n_175)
);


endmodule