module fake_jpeg_31407_n_503 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_22),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_78),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_57),
.B(n_80),
.Y(n_157)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_39),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_2),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_3),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_29),
.B(n_13),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_97),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_46),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_117),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_50),
.C(n_51),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_126),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_145),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_93),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_49),
.B1(n_43),
.B2(n_45),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_59),
.B1(n_53),
.B2(n_61),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_51),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_154),
.B(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_159),
.B(n_161),
.Y(n_249)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_76),
.B(n_100),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_48),
.B(n_23),
.C(n_42),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_162),
.B(n_171),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_163),
.A2(n_167),
.B1(n_184),
.B2(n_185),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_107),
.B1(n_66),
.B2(n_73),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_103),
.A2(n_89),
.B1(n_96),
.B2(n_94),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_168),
.A2(n_83),
.B1(n_86),
.B2(n_95),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_118),
.B(n_68),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_170),
.B(n_209),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_24),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_48),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_200),
.Y(n_213)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_84),
.B1(n_140),
.B2(n_71),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_19),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_188),
.Y(n_220)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_104),
.B(n_19),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_157),
.B(n_40),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_197),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_19),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_124),
.B1(n_146),
.B2(n_138),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_153),
.B1(n_146),
.B2(n_138),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_19),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_42),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_121),
.B(n_40),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_101),
.A2(n_49),
.B1(n_31),
.B2(n_79),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_131),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_208),
.Y(n_215)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_145),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_137),
.A2(n_31),
.B1(n_34),
.B2(n_43),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_62),
.B1(n_63),
.B2(n_106),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_119),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_171),
.Y(n_228)
);

NAND2x1p5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_63),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_214),
.B(n_221),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_230),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_88),
.B(n_62),
.Y(n_221)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_243),
.B1(n_250),
.B2(n_169),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_239),
.Y(n_266)
);

XOR2x1_ASAP7_75t_SL g229 ( 
.A(n_162),
.B(n_131),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_229),
.A2(n_39),
.B(n_46),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_124),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_129),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_170),
.B1(n_195),
.B2(n_169),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_167),
.A2(n_129),
.B1(n_147),
.B2(n_144),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_160),
.B(n_111),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_246),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_168),
.B1(n_170),
.B2(n_173),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_188),
.A2(n_111),
.B1(n_127),
.B2(n_106),
.Y(n_251)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_263),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_258),
.A2(n_281),
.B1(n_243),
.B2(n_250),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_268),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_168),
.B1(n_147),
.B2(n_144),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_211),
.B1(n_227),
.B2(n_237),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_218),
.B(n_196),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_273),
.B1(n_240),
.B2(n_246),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_201),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_176),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_271),
.B(n_281),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_222),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_272),
.B(n_282),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_191),
.B1(n_187),
.B2(n_190),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_178),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_215),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_165),
.B1(n_172),
.B2(n_181),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_213),
.B(n_191),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_246),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_289),
.Y(n_302)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_241),
.A2(n_194),
.B(n_179),
.C(n_166),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_213),
.B(n_165),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_174),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_225),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_221),
.Y(n_305)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_219),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_288),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_249),
.C(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_297),
.B(n_298),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_249),
.C(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_252),
.C(n_214),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_300),
.B(n_310),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_312),
.B1(n_322),
.B2(n_321),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_305),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_214),
.B(n_221),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_317),
.B(n_326),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_308),
.A2(n_313),
.B1(n_315),
.B2(n_325),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_225),
.C(n_177),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_258),
.A2(n_211),
.B1(n_223),
.B2(n_212),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_264),
.A2(n_235),
.B1(n_231),
.B2(n_219),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_282),
.B1(n_278),
.B2(n_255),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_271),
.B(n_256),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_224),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_284),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_283),
.A2(n_205),
.B1(n_235),
.B2(n_231),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_255),
.A2(n_245),
.B1(n_202),
.B2(n_224),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_257),
.A2(n_286),
.B(n_256),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_280),
.A2(n_245),
.B1(n_193),
.B2(n_127),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_277),
.B1(n_272),
.B2(n_269),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_286),
.B(n_268),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_325),
.B1(n_299),
.B2(n_322),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_303),
.B(n_266),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_348),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_333),
.B(n_349),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_346),
.B1(n_347),
.B2(n_355),
.Y(n_366)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_256),
.B1(n_265),
.B2(n_261),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_341),
.A2(n_358),
.B1(n_279),
.B2(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_327),
.B(n_266),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_345),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_304),
.B(n_263),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_326),
.A2(n_261),
.B1(n_274),
.B2(n_276),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_285),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_290),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_311),
.B(n_293),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_351),
.B(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_87),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_296),
.A2(n_300),
.B1(n_316),
.B2(n_313),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_132),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_261),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_279),
.B1(n_34),
.B2(n_45),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_194),
.B(n_142),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_314),
.B(n_318),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_270),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_297),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_377),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_302),
.Y(n_364)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_310),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_340),
.Y(n_370)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_298),
.C(n_329),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_333),
.C(n_337),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_305),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_375),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_343),
.B(n_294),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_307),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_323),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_378),
.A2(n_386),
.B(n_356),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_379),
.A2(n_381),
.B1(n_334),
.B2(n_335),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_318),
.Y(n_385)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_357),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_388),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_355),
.B(n_295),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_270),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_369),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_405),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_395),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_368),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_400),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_347),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_409),
.C(n_412),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_366),
.A2(n_331),
.B1(n_341),
.B2(n_358),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_403),
.B1(n_381),
.B2(n_378),
.Y(n_436)
);

AOI21xp33_ASAP7_75t_L g400 ( 
.A1(n_384),
.A2(n_330),
.B(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_366),
.A2(n_374),
.B1(n_387),
.B2(n_383),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_330),
.B(n_352),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_347),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_410),
.A2(n_367),
.B1(n_363),
.B2(n_383),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_380),
.A2(n_356),
.B1(n_353),
.B2(n_354),
.Y(n_411)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_411),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_353),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_334),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_416),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_359),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_377),
.C(n_386),
.Y(n_419)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_378),
.B(n_390),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_395),
.B(n_412),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_398),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_399),
.B1(n_413),
.B2(n_416),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_409),
.C(n_393),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_433),
.C(n_415),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_363),
.B1(n_367),
.B2(n_376),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_429),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_390),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_390),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_397),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_385),
.C(n_378),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_382),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_436),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_439),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_438),
.Y(n_454)
);

OAI321xp33_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_435),
.A3(n_430),
.B1(n_429),
.B2(n_436),
.C(n_410),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_442),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_392),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_446),
.Y(n_464)
);

INVx11_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_420),
.B(n_394),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_450),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_392),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_419),
.B(n_382),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_418),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_391),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_433),
.A2(n_391),
.B(n_183),
.Y(n_452)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

AOI22x1_ASAP7_75t_L g453 ( 
.A1(n_427),
.A2(n_189),
.B1(n_139),
.B2(n_142),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_453),
.B(n_145),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_451),
.A2(n_426),
.B1(n_417),
.B2(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_465),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_431),
.B(n_434),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_451),
.A2(n_418),
.B1(n_423),
.B2(n_34),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_460),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_139),
.C(n_45),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_446),
.C(n_443),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_449),
.B(n_3),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_4),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_448),
.Y(n_469)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_447),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_471),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_444),
.B(n_442),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_464),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_453),
.C(n_38),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_46),
.C(n_8),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_38),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_5),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_468),
.B(n_6),
.Y(n_477)
);

AOI31xp33_ASAP7_75t_L g484 ( 
.A1(n_477),
.A2(n_456),
.A3(n_454),
.B(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_7),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_482),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_467),
.Y(n_482)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_484),
.A2(n_486),
.A3(n_480),
.B1(n_473),
.B2(n_478),
.C1(n_10),
.C2(n_11),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_485),
.Y(n_491)
);

A2O1A1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_474),
.A2(n_464),
.B(n_459),
.C(n_463),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_487),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_493),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_488),
.B(n_480),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_490),
.B(n_482),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_495),
.B1(n_481),
.B2(n_491),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_492),
.B(n_483),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_498),
.B(n_8),
.Y(n_499)
);

AOI322xp5_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_486),
.A3(n_478),
.B1(n_493),
.B2(n_12),
.C1(n_8),
.C2(n_11),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_10),
.B(n_11),
.Y(n_500)
);

A2O1A1O1Ixp25_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_10),
.B(n_11),
.C(n_12),
.D(n_46),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_25),
.B(n_430),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_25),
.C(n_121),
.Y(n_503)
);


endmodule