module fake_jpeg_7681_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_17),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_61),
.Y(n_83)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_65),
.Y(n_84)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_21),
.B1(n_17),
.B2(n_65),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_33),
.B(n_38),
.C(n_23),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_27),
.B(n_29),
.C(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_85),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_24),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_58),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_93),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_71),
.B1(n_69),
.B2(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_104),
.B(n_20),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_64),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_27),
.B(n_28),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_31),
.B1(n_15),
.B2(n_45),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_26),
.B(n_20),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_58),
.B1(n_31),
.B2(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_15),
.B1(n_69),
.B2(n_72),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_78),
.C(n_82),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.C(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_82),
.C(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_91),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_100),
.B1(n_104),
.B2(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_103),
.B1(n_99),
.B2(n_72),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_71),
.B1(n_15),
.B2(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_63),
.B1(n_59),
.B2(n_29),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_81),
.B(n_20),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_127),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_20),
.B(n_26),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_53),
.C(n_62),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_89),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_148),
.C(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_109),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_150),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_90),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_110),
.A3(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_153),
.B1(n_120),
.B2(n_121),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_35),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_89),
.B1(n_97),
.B2(n_35),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_141),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_174),
.B1(n_149),
.B2(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_160),
.B1(n_164),
.B2(n_155),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_133),
.B1(n_131),
.B2(n_112),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_129),
.C(n_123),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_173),
.C(n_152),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_128),
.B(n_126),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_135),
.B(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_131),
.B1(n_129),
.B2(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_158),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_127),
.B(n_114),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_117),
.B(n_26),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_132),
.C(n_124),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_146),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_186),
.B(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_185),
.B1(n_164),
.B2(n_173),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_188),
.B(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_148),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.C(n_189),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_101),
.B(n_79),
.C(n_77),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_117),
.C(n_54),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_101),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_101),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_0),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_196),
.B1(n_178),
.B2(n_186),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_202),
.B(n_41),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_170),
.B1(n_175),
.B2(n_165),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_165),
.C(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_204),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_4),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_174),
.C(n_48),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_19),
.B1(n_22),
.B2(n_77),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_79),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_187),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_212),
.C(n_197),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_202),
.B(n_198),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_214),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_193),
.B(n_206),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_79),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_200),
.C(n_6),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_222),
.B(n_225),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_226),
.Y(n_231)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_199),
.B(n_217),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_9),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_5),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_200),
.B(n_6),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_208),
.B1(n_216),
.B2(n_9),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_232),
.B(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_5),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_8),
.B(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_13),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_231),
.B(n_12),
.C(n_13),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_10),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_12),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_10),
.B(n_12),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.C(n_235),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_240),
.B(n_13),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_244),
.Y(n_246)
);


endmodule