module real_jpeg_23425_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_39),
.B1(n_65),
.B2(n_70),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_53),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_3),
.A2(n_30),
.B(n_33),
.C(n_245),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_185),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_3),
.B(n_65),
.C(n_68),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_185),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_3),
.A2(n_102),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_36),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_5),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_89),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_89),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_5),
.A2(n_65),
.B1(n_70),
.B2(n_89),
.Y(n_205)
);

INVx8_ASAP7_75t_SL g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_43),
.B1(n_56),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_7),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_145),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_7),
.A2(n_65),
.B1(n_70),
.B2(n_145),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_10),
.A2(n_56),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_81),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_81),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_10),
.A2(n_65),
.B1(n_70),
.B2(n_81),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_55),
.B1(n_65),
.B2(n_70),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_12),
.A2(n_43),
.B1(n_51),
.B2(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_12),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_120),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_120),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_12),
.A2(n_65),
.B1(n_70),
.B2(n_120),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_13),
.A2(n_45),
.B1(n_56),
.B2(n_175),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_175),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_13),
.A2(n_65),
.B1(n_70),
.B2(n_175),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_15),
.A2(n_46),
.B1(n_65),
.B2(n_70),
.Y(n_193)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_16),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_16),
.A2(n_103),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_16),
.A2(n_103),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_95),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_21),
.B(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_37),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_24),
.A2(n_36),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_24),
.A2(n_36),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_24),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_25),
.A2(n_26),
.B1(n_93),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_25),
.A2(n_26),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_25),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_25),
.A2(n_214),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_26),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_26),
.A2(n_141),
.B(n_200),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_28),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_27),
.A2(n_31),
.B(n_185),
.Y(n_245)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_28),
.B(n_266),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_SL g196 ( 
.A(n_33),
.B(n_50),
.C(n_58),
.Y(n_196)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_34),
.A2(n_49),
.B(n_186),
.C(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_36),
.B(n_201),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_52),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_44),
.B(n_185),
.Y(n_186)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_47),
.A2(n_147),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_47),
.A2(n_53),
.B1(n_144),
.B2(n_217),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_78),
.B1(n_79),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_88),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_52),
.B(n_119),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_52),
.A2(n_117),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_57),
.Y(n_184)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_75),
.C(n_77),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_75),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_87),
.C(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_62),
.A2(n_86),
.B1(n_91),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_71),
.B(n_73),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_71),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_71),
.B1(n_111),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_63),
.B(n_181),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_63),
.A2(n_71),
.B1(n_240),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_64),
.A2(n_74),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_64),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_64),
.A2(n_126),
.B1(n_139),
.B2(n_179),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_64),
.B(n_185),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_64),
.A2(n_180),
.B(n_255),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_70),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_71),
.B(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_90),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_83),
.A2(n_87),
.B1(n_157),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_87),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_91),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI31xp33_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_158),
.A3(n_164),
.B(n_345),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_148),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_98),
.B(n_148),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_121),
.C(n_129),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_99),
.A2(n_121),
.B1(n_122),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_99),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_113),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_101),
.B(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_101),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B(n_108),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_108),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_102),
.A2(n_192),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_102),
.A2(n_105),
.B1(n_134),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_102),
.A2(n_274),
.B(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_103),
.B(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_106),
.B(n_185),
.Y(n_278)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B(n_128),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_126),
.A2(n_239),
.B(n_241),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_126),
.A2(n_241),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_129),
.A2(n_130),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.C(n_142),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_131),
.A2(n_132),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_133),
.Y(n_317)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_135),
.A2(n_248),
.B(n_272),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_140),
.B(n_142),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_159),
.A2(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_160),
.B(n_163),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_338),
.B(n_344),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_328),
.B(n_337),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_226),
.B(n_311),
.C(n_327),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_209),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_168),
.B(n_209),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_187),
.C(n_197),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_169),
.A2(n_170),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_182),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_177),
.C(n_182),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B(n_186),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_187),
.A2(n_188),
.B1(n_197),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_194),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_197),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.C(n_204),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_218),
.B1(n_219),
.B2(n_225),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_210),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.CI(n_215),
.CON(n_210),
.SN(n_210)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_212),
.C(n_215),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_220),
.B(n_224),
.C(n_225),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_221),
.B(n_223),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_304),
.B(n_310),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_259),
.B(n_303),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_251),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_231),
.B(n_251),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_250),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_232),
.B(n_238),
.C(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.C(n_256),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_256),
.B1(n_257),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_297),
.B(n_302),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_287),
.B(n_296),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_275),
.B(n_286),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_282),
.B(n_285),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_326),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_323),
.C(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_333),
.C(n_336),
.Y(n_343)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_343),
.Y(n_344)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);


endmodule