module fake_jpeg_3513_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_5),
.Y(n_78)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_18),
.A2(n_3),
.B(n_5),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_15),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_20),
.B1(n_25),
.B2(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_80),
.B1(n_51),
.B2(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_36),
.A2(n_24),
.B1(n_13),
.B2(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_7),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_5),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_42),
.B1(n_40),
.B2(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_69),
.B1(n_65),
.B2(n_64),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_88),
.B1(n_93),
.B2(n_101),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_49),
.B1(n_13),
.B2(n_15),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_41),
.B1(n_45),
.B2(n_15),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_74),
.B1(n_73),
.B2(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_6),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_6),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_104),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_7),
.B1(n_8),
.B2(n_73),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_77),
.B(n_75),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_74),
.C(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_114),
.B1(n_122),
.B2(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_83),
.B1(n_102),
.B2(n_99),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_53),
.B1(n_69),
.B2(n_64),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_53),
.B1(n_65),
.B2(n_55),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_90),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_89),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_122),
.B1(n_114),
.B2(n_109),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_133),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_100),
.B(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_136),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_93),
.B1(n_104),
.B2(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_91),
.C(n_94),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_110),
.B1(n_118),
.B2(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_146),
.B1(n_141),
.B2(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_135),
.B(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_154),
.B1(n_152),
.B2(n_148),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_125),
.B1(n_124),
.B2(n_129),
.C(n_118),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_96),
.A3(n_126),
.B1(n_95),
.B2(n_86),
.C1(n_143),
.C2(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_123),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_159),
.B(n_152),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_144),
.B1(n_127),
.B2(n_130),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_158),
.B(n_157),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_113),
.B1(n_119),
.B2(n_105),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_159),
.C(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.C(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_113),
.C(n_119),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_162),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_170),
.B(n_105),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);


endmodule