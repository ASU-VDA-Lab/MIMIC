module fake_jpeg_1991_n_258 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_1),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_64),
.C(n_26),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_51),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_67),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_2),
.C(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_64),
.Y(n_108)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_99),
.Y(n_129)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_17),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_102),
.C(n_51),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_38),
.B1(n_36),
.B2(n_22),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_104),
.B1(n_61),
.B2(n_52),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_38),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_18),
.B1(n_23),
.B2(n_30),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_130),
.Y(n_159)
);

OR2x2_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_51),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_46),
.B1(n_44),
.B2(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_104),
.B1(n_83),
.B2(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_68),
.B(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_14),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_3),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_57),
.B1(n_30),
.B2(n_56),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_18),
.B1(n_27),
.B2(n_50),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_73),
.B1(n_100),
.B2(n_18),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_50),
.C(n_51),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_134),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_50),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_82),
.B(n_77),
.C(n_18),
.D(n_27),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_4),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_148),
.B1(n_113),
.B2(n_135),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_157),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_83),
.B(n_100),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_103),
.B1(n_101),
.B2(n_73),
.Y(n_148)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_80),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_80),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_101),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_122),
.B1(n_82),
.B2(n_77),
.Y(n_175)
);

AO21x1_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_136),
.B(n_131),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_116),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_157),
.A3(n_139),
.B1(n_149),
.B2(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_170),
.B1(n_175),
.B2(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_173),
.Y(n_200)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_134),
.B1(n_132),
.B2(n_119),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_133),
.B1(n_125),
.B2(n_106),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_160),
.B1(n_146),
.B2(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_182),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_114),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_140),
.C(n_128),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_106),
.B1(n_124),
.B2(n_135),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_152),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_118),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_148),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_162),
.B(n_150),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_150),
.B(n_143),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_185),
.B(n_181),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_159),
.B(n_144),
.C(n_158),
.D(n_142),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_190),
.B(n_177),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_201),
.C(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_166),
.B1(n_180),
.B2(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_140),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_155),
.C(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_214),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_213),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_198),
.B1(n_192),
.B2(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_219),
.B1(n_200),
.B2(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_170),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_181),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_168),
.C(n_138),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_204),
.C(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_227),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_196),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_229),
.Y(n_231)
);

OR2x6_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_194),
.C(n_190),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_193),
.C(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_218),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_197),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_225),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_216),
.C(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_207),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_224),
.C(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_243),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_245),
.B(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_220),
.C(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_234),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_203),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_203),
.C(n_5),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_239),
.Y(n_250)
);

O2A1O1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_250),
.A2(n_244),
.B(n_203),
.C(n_10),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_247),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_253),
.B1(n_203),
.B2(n_6),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_5),
.Y(n_258)
);


endmodule