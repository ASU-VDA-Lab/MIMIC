module fake_jpeg_14343_n_203 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx11_ASAP7_75t_SL g82 ( 
.A(n_46),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_0),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_93),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_1),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_72),
.Y(n_122)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_110),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_73),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_117),
.B1(n_123),
.B2(n_128),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_89),
.B1(n_87),
.B2(n_73),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_57),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_73),
.B1(n_64),
.B2(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_70),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_133),
.C(n_96),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_63),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_130),
.B(n_132),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_84),
.B1(n_85),
.B2(n_61),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_84),
.B1(n_85),
.B2(n_61),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_34),
.B1(n_52),
.B2(n_51),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_75),
.B(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_58),
.B1(n_80),
.B2(n_79),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_62),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_66),
.A3(n_60),
.B1(n_82),
.B2(n_76),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_137),
.B(n_145),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_60),
.B(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2x1p5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_16),
.Y(n_164)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_151),
.B(n_15),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_116),
.B1(n_124),
.B2(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_148),
.B1(n_156),
.B2(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_151)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2x1_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_16),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_13),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_14),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_171),
.B1(n_141),
.B2(n_155),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_36),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_170),
.C(n_30),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_167),
.B(n_140),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_19),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_153),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_20),
.C(n_25),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_184),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_152),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_181),
.C(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_183),
.Y(n_189)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_163),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_161),
.A3(n_162),
.B1(n_166),
.B2(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_171),
.C(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_181),
.C(n_167),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_177),
.Y(n_194)
);

FAx1_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_194),
.CI(n_188),
.CON(n_196),
.SN(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_189),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_186),
.B1(n_173),
.B2(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_38),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_170),
.C(n_44),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_42),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_45),
.Y(n_203)
);


endmodule