module fake_jpeg_12369_n_75 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

OR2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_22),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_1),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_2),
.B(n_3),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_12),
.C(n_21),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_55),
.C(n_58),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_2),
.B(n_3),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_56),
.B(n_5),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_13),
.B1(n_20),
.B2(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_43),
.B(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_65),
.B1(n_8),
.B2(n_10),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_66),
.B1(n_64),
.B2(n_24),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_64),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_68),
.CI(n_15),
.CON(n_73),
.SN(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_18),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_73),
.Y(n_75)
);


endmodule