module fake_jpeg_24049_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_22),
.B(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_34),
.Y(n_37)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_1),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_20),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_16),
.B(n_23),
.Y(n_36)
);

XNOR2x1_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_24),
.B1(n_32),
.B2(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_12),
.B1(n_18),
.B2(n_21),
.Y(n_53)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_50),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_27),
.C(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_51),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_31),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_37),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_62),
.C(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_58),
.B1(n_51),
.B2(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_76),
.B1(n_69),
.B2(n_67),
.Y(n_86)
);

NAND2x1_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_58),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_72),
.B(n_46),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_55),
.B1(n_45),
.B2(n_47),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.C(n_63),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_45),
.C(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_75),
.C(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_87),
.C(n_77),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_82),
.B(n_93),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_92),
.B(n_78),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_74),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_80),
.B(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_27),
.B1(n_4),
.B2(n_7),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_25),
.C(n_44),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_107),
.B(n_102),
.C(n_105),
.D(n_103),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_2),
.Y(n_111)
);


endmodule