module real_aes_6984_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_0), .A2(n_13), .B1(n_161), .B2(n_163), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_1), .Y(n_87) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_2), .A2(n_75), .B1(n_154), .B2(n_157), .Y(n_153) );
INVx1_ASAP7_75t_L g267 ( .A(n_3), .Y(n_267) );
AOI21xp33_ASAP7_75t_L g247 ( .A1(n_4), .A2(n_205), .B(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g188 ( .A(n_6), .Y(n_188) );
AND2x6_ASAP7_75t_L g210 ( .A(n_6), .B(n_186), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_6), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_7), .A2(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g254 ( .A(n_8), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_9), .B(n_298), .Y(n_297) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_10), .A2(n_28), .B1(n_93), .B2(n_94), .Y(n_92) );
INVx1_ASAP7_75t_L g203 ( .A(n_11), .Y(n_203) );
INVx1_ASAP7_75t_L g312 ( .A(n_12), .Y(n_312) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_14), .A2(n_30), .B1(n_93), .B2(n_97), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_15), .B(n_218), .Y(n_323) );
INVx1_ASAP7_75t_L g534 ( .A(n_15), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_16), .B(n_205), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_17), .B(n_226), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_18), .A2(n_26), .B1(n_138), .B2(n_140), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_19), .A2(n_310), .B(n_311), .C(n_313), .Y(n_309) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_20), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_21), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_22), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_23), .B(n_252), .Y(n_269) );
INVx1_ASAP7_75t_L g241 ( .A(n_24), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_25), .A2(n_49), .B1(n_145), .B2(n_148), .Y(n_144) );
INVx2_ASAP7_75t_L g208 ( .A(n_27), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g172 ( .A1(n_29), .A2(n_47), .B1(n_173), .B2(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_29), .Y(n_174) );
OAI221xp5_ASAP7_75t_L g179 ( .A1(n_30), .A2(n_40), .B1(n_48), .B2(n_180), .C(n_181), .Y(n_179) );
INVxp67_ASAP7_75t_L g182 ( .A(n_30), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_31), .A2(n_210), .B(n_213), .C(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g239 ( .A(n_32), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_33), .A2(n_73), .B1(n_116), .B2(n_120), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_34), .B(n_252), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_34), .A2(n_82), .B1(n_83), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_34), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_35), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_36), .B(n_205), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_37), .A2(n_213), .B1(n_235), .B2(n_237), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_38), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_39), .Y(n_264) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_40), .A2(n_58), .B1(n_93), .B2(n_97), .Y(n_102) );
INVxp67_ASAP7_75t_L g183 ( .A(n_40), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_41), .A2(n_222), .B(n_251), .C(n_253), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_42), .Y(n_326) );
INVx1_ASAP7_75t_L g249 ( .A(n_43), .Y(n_249) );
INVx1_ASAP7_75t_L g186 ( .A(n_44), .Y(n_186) );
INVx1_ASAP7_75t_L g202 ( .A(n_45), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_46), .Y(n_180) );
INVx1_ASAP7_75t_L g173 ( .A(n_47), .Y(n_173) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_48), .A2(n_63), .B1(n_93), .B2(n_94), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_SL g217 ( .A1(n_50), .A2(n_218), .B(n_219), .C(n_222), .Y(n_217) );
INVxp67_ASAP7_75t_L g220 ( .A(n_51), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_52), .A2(n_70), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_52), .Y(n_170) );
INVx1_ASAP7_75t_L g81 ( .A(n_53), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_54), .Y(n_245) );
INVx1_ASAP7_75t_L g319 ( .A(n_55), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_56), .A2(n_82), .B1(n_83), .B2(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_56), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_57), .A2(n_210), .B(n_213), .C(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_59), .B(n_268), .Y(n_281) );
INVx2_ASAP7_75t_L g200 ( .A(n_60), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_61), .B(n_218), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_62), .A2(n_210), .B(n_213), .C(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_64), .B(n_256), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_65), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_66), .A2(n_210), .B(n_213), .C(n_295), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_67), .Y(n_302) );
INVx1_ASAP7_75t_L g216 ( .A(n_68), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_69), .Y(n_308) );
INVx1_ASAP7_75t_L g171 ( .A(n_70), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_70), .B(n_268), .Y(n_296) );
INVx1_ASAP7_75t_L g93 ( .A(n_71), .Y(n_93) );
INVx1_ASAP7_75t_L g95 ( .A(n_71), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_72), .B(n_198), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_74), .A2(n_205), .B(n_211), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_76), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_176), .B1(n_189), .B2(n_514), .C(n_522), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_167), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_135), .Y(n_84) );
NOR3xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_108), .C(n_124), .Y(n_85) );
OAI22xp5_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_88), .B1(n_103), .B2(n_104), .Y(n_86) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
OR2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
INVx2_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
OR2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_96), .Y(n_90) );
AND2x2_ASAP7_75t_L g107 ( .A(n_91), .B(n_96), .Y(n_107) );
AND2x2_ASAP7_75t_L g143 ( .A(n_91), .B(n_131), .Y(n_143) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g111 ( .A(n_92), .B(n_96), .Y(n_111) );
AND2x2_ASAP7_75t_L g119 ( .A(n_92), .B(n_102), .Y(n_119) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_95), .Y(n_97) );
INVx2_ASAP7_75t_L g131 ( .A(n_96), .Y(n_131) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
NAND2x1p5_ASAP7_75t_L g106 ( .A(n_99), .B(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g162 ( .A(n_99), .B(n_143), .Y(n_162) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_101), .Y(n_99) );
INVx1_ASAP7_75t_L g113 ( .A(n_100), .Y(n_113) );
INVx1_ASAP7_75t_L g118 ( .A(n_100), .Y(n_118) );
INVx1_ASAP7_75t_L g123 ( .A(n_100), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_100), .B(n_102), .Y(n_151) );
AND2x2_ASAP7_75t_L g112 ( .A(n_101), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g142 ( .A(n_102), .B(n_123), .Y(n_142) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g156 ( .A(n_107), .B(n_112), .Y(n_156) );
AND2x2_ASAP7_75t_L g159 ( .A(n_107), .B(n_142), .Y(n_159) );
OAI21xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_114), .B(n_115), .Y(n_108) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x4_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_L g138 ( .A(n_112), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g147 ( .A(n_112), .B(n_143), .Y(n_147) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g130 ( .A(n_118), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g129 ( .A(n_119), .B(n_130), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_119), .B(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_132), .B2(n_133), .Y(n_124) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_152), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_144), .Y(n_136) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x4_ASAP7_75t_L g149 ( .A(n_143), .B(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x6_ASAP7_75t_L g165 ( .A(n_151), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_160), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx8_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx6_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B1(n_172), .B2(n_175), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_172), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
AND3x1_ASAP7_75t_SL g178 ( .A(n_179), .B(n_184), .C(n_187), .Y(n_178) );
INVxp67_ASAP7_75t_L g528 ( .A(n_179), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx1_ASAP7_75t_SL g530 ( .A(n_184), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_184), .A2(n_517), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_184), .Y(n_540) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_185), .B(n_188), .Y(n_533) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_SL g539 ( .A(n_187), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_191), .B(n_451), .Y(n_190) );
NOR4xp25_ASAP7_75t_L g191 ( .A(n_192), .B(n_381), .C(n_412), .D(n_431), .Y(n_191) );
NAND4xp25_ASAP7_75t_L g192 ( .A(n_193), .B(n_339), .C(n_354), .D(n_372), .Y(n_192) );
AOI222xp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_274), .B1(n_315), .B2(n_327), .C1(n_332), .C2(n_334), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_257), .Y(n_194) );
INVx1_ASAP7_75t_L g395 ( .A(n_195), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_228), .Y(n_195) );
AND2x2_ASAP7_75t_L g258 ( .A(n_196), .B(n_246), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_196), .B(n_261), .Y(n_424) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g331 ( .A(n_197), .B(n_230), .Y(n_331) );
AND2x2_ASAP7_75t_L g340 ( .A(n_197), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g366 ( .A(n_197), .Y(n_366) );
AND2x2_ASAP7_75t_L g387 ( .A(n_197), .B(n_230), .Y(n_387) );
BUFx2_ASAP7_75t_L g410 ( .A(n_197), .Y(n_410) );
AND2x2_ASAP7_75t_L g434 ( .A(n_197), .B(n_231), .Y(n_434) );
AND2x2_ASAP7_75t_L g498 ( .A(n_197), .B(n_246), .Y(n_498) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_204), .B(n_225), .Y(n_197) );
INVx4_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_200), .B(n_201), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
BUFx2_ASAP7_75t_L g306 ( .A(n_205), .Y(n_306) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_206), .B(n_210), .Y(n_243) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_209), .Y(n_206) );
INVx1_ASAP7_75t_L g519 ( .A(n_207), .Y(n_519) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g214 ( .A(n_208), .Y(n_214) );
INVx1_ASAP7_75t_L g236 ( .A(n_208), .Y(n_236) );
INVx1_ASAP7_75t_L g215 ( .A(n_209), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_209), .Y(n_218) );
INVx3_ASAP7_75t_L g221 ( .A(n_209), .Y(n_221) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_209), .Y(n_238) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_209), .Y(n_252) );
INVx4_ASAP7_75t_SL g224 ( .A(n_210), .Y(n_224) );
BUFx3_ASAP7_75t_L g516 ( .A(n_210), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_216), .B(n_217), .C(n_224), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_212), .A2(n_224), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_212), .A2(n_224), .B(n_308), .C(n_309), .Y(n_307) );
INVx5_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_214), .Y(n_223) );
BUFx3_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_221), .B(n_254), .Y(n_253) );
INVx5_ASAP7_75t_L g268 ( .A(n_221), .Y(n_268) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_224), .A2(n_234), .B1(n_242), .B2(n_243), .Y(n_233) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_226), .A2(n_247), .B(n_255), .Y(n_246) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_SL g287 ( .A(n_227), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g399 ( .A(n_228), .B(n_330), .Y(n_399) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_229), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_246), .Y(n_229) );
OR2x2_ASAP7_75t_L g359 ( .A(n_230), .B(n_262), .Y(n_359) );
AND2x2_ASAP7_75t_L g371 ( .A(n_230), .B(n_330), .Y(n_371) );
BUFx2_ASAP7_75t_L g503 ( .A(n_230), .Y(n_503) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g260 ( .A(n_231), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g353 ( .A(n_231), .B(n_262), .Y(n_353) );
AND2x2_ASAP7_75t_L g406 ( .A(n_231), .B(n_246), .Y(n_406) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_231), .Y(n_442) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_244), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_232), .B(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_232), .A2(n_263), .B(n_271), .Y(n_262) );
INVx2_ASAP7_75t_L g286 ( .A(n_232), .Y(n_286) );
INVx2_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_237) );
INVx2_ASAP7_75t_L g240 ( .A(n_238), .Y(n_240) );
INVx4_ASAP7_75t_L g310 ( .A(n_238), .Y(n_310) );
INVx2_ASAP7_75t_L g521 ( .A(n_240), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_243), .A2(n_264), .B(n_265), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_243), .A2(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g329 ( .A(n_246), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g341 ( .A(n_246), .Y(n_341) );
INVx2_ASAP7_75t_L g352 ( .A(n_246), .Y(n_352) );
BUFx2_ASAP7_75t_L g376 ( .A(n_246), .Y(n_376) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_246), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx4_ASAP7_75t_L g298 ( .A(n_252), .Y(n_298) );
INVx1_ASAP7_75t_L g273 ( .A(n_256), .Y(n_273) );
INVx2_ASAP7_75t_L g292 ( .A(n_256), .Y(n_292) );
OA21x2_ASAP7_75t_L g304 ( .A1(n_256), .A2(n_305), .B(n_314), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AOI332xp33_ASAP7_75t_L g354 ( .A1(n_258), .A2(n_355), .A3(n_359), .B1(n_360), .B2(n_364), .B3(n_367), .C1(n_368), .C2(n_370), .Y(n_354) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_258), .B(n_330), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_258), .B(n_344), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_SL g372 ( .A1(n_259), .A2(n_373), .B(n_376), .C(n_377), .Y(n_372) );
AND2x2_ASAP7_75t_L g511 ( .A(n_259), .B(n_352), .Y(n_511) );
INVx3_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g408 ( .A(n_260), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g413 ( .A(n_260), .B(n_410), .Y(n_413) );
INVx1_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
AND2x2_ASAP7_75t_L g447 ( .A(n_261), .B(n_406), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_261), .B(n_387), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_261), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_261), .B(n_365), .Y(n_473) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g330 ( .A(n_262), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_269), .C(n_270), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_273), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_273), .B(n_326), .Y(n_325) );
OAI31xp33_ASAP7_75t_L g512 ( .A1(n_274), .A2(n_433), .A3(n_440), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_289), .Y(n_274) );
AND2x2_ASAP7_75t_L g315 ( .A(n_275), .B(n_316), .Y(n_315) );
NAND2x1_ASAP7_75t_SL g335 ( .A(n_275), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_275), .Y(n_422) );
AND2x2_ASAP7_75t_L g427 ( .A(n_275), .B(n_338), .Y(n_427) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_276), .A2(n_340), .B(n_342), .C(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g356 ( .A(n_276), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g369 ( .A(n_276), .Y(n_369) );
AND2x2_ASAP7_75t_L g375 ( .A(n_276), .B(n_317), .Y(n_375) );
INVx2_ASAP7_75t_L g393 ( .A(n_276), .Y(n_393) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_358), .Y(n_404) );
AND2x2_ASAP7_75t_L g436 ( .A(n_276), .B(n_394), .Y(n_436) );
AND2x2_ASAP7_75t_L g440 ( .A(n_276), .B(n_363), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_276), .B(n_289), .Y(n_445) );
AND2x2_ASAP7_75t_L g479 ( .A(n_276), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_276), .B(n_382), .Y(n_513) );
OR2x6_ASAP7_75t_L g276 ( .A(n_277), .B(n_287), .Y(n_276) );
AOI21xp5_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_279), .B(n_286), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_283), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_283), .A2(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_289), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g421 ( .A(n_289), .Y(n_421) );
AND2x2_ASAP7_75t_L g483 ( .A(n_289), .B(n_404), .Y(n_483) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_303), .Y(n_289) );
OR2x2_ASAP7_75t_L g337 ( .A(n_290), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g347 ( .A(n_290), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_290), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g455 ( .A(n_290), .Y(n_455) );
AND2x2_ASAP7_75t_L g472 ( .A(n_290), .B(n_317), .Y(n_472) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g363 ( .A(n_291), .B(n_303), .Y(n_363) );
AND2x2_ASAP7_75t_L g392 ( .A(n_291), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g403 ( .A(n_291), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_291), .B(n_358), .Y(n_494) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_301), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_300), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g316 ( .A(n_304), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
AND2x2_ASAP7_75t_L g394 ( .A(n_304), .B(n_358), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_310), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g496 ( .A(n_315), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_316), .Y(n_500) );
INVx2_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_324), .B(n_325), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_329), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_329), .B(n_434), .Y(n_492) );
OR2x2_ASAP7_75t_L g333 ( .A(n_330), .B(n_331), .Y(n_333) );
INVx1_ASAP7_75t_SL g385 ( .A(n_330), .Y(n_385) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_336), .A2(n_389), .B1(n_391), .B2(n_395), .C(n_396), .Y(n_388) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g416 ( .A(n_337), .B(n_380), .Y(n_416) );
INVx2_ASAP7_75t_L g348 ( .A(n_338), .Y(n_348) );
INVx1_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_338), .B(n_358), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_338), .B(n_361), .Y(n_468) );
INVx1_ASAP7_75t_L g476 ( .A(n_338), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_340), .B(n_344), .Y(n_390) );
AND2x4_ASAP7_75t_L g365 ( .A(n_341), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g478 ( .A(n_344), .B(n_434), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_347), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g486 ( .A(n_348), .Y(n_486) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g386 ( .A(n_352), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g458 ( .A(n_352), .B(n_434), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_352), .B(n_371), .Y(n_464) );
AOI322xp5_ASAP7_75t_L g418 ( .A1(n_353), .A2(n_387), .A3(n_394), .B1(n_419), .B2(n_422), .C1(n_423), .C2(n_425), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_353), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g484 ( .A(n_356), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
INVx2_ASAP7_75t_L g361 ( .A(n_358), .Y(n_361) );
INVx1_ASAP7_75t_L g420 ( .A(n_358), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_359), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g456 ( .A(n_361), .B(n_369), .Y(n_456) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g368 ( .A(n_363), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g411 ( .A(n_363), .B(n_404), .Y(n_411) );
AND2x2_ASAP7_75t_L g415 ( .A(n_363), .B(n_375), .Y(n_415) );
OAI21xp33_ASAP7_75t_SL g425 ( .A1(n_364), .A2(n_426), .B(n_428), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_364), .A2(n_496), .B1(n_497), .B2(n_499), .Y(n_495) );
INVx3_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g370 ( .A(n_365), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_365), .B(n_385), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_367), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g507 ( .A(n_374), .Y(n_507) );
INVx4_ASAP7_75t_L g380 ( .A(n_375), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_375), .B(n_402), .Y(n_450) );
INVx1_ASAP7_75t_SL g462 ( .A(n_376), .Y(n_462) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_380), .B(n_476), .Y(n_475) );
OAI211xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_383), .B(n_388), .C(n_405), .Y(n_381) );
OAI221xp5_ASAP7_75t_SL g501 ( .A1(n_383), .A2(n_421), .B1(n_500), .B2(n_502), .C(n_504), .Y(n_501) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_385), .B(n_498), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g477 ( .A1(n_386), .A2(n_463), .A3(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g467 ( .A(n_392), .Y(n_467) );
AND2x2_ASAP7_75t_L g480 ( .A(n_394), .B(n_403), .Y(n_480) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_404), .B(n_507), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_417), .C(n_418), .Y(n_412) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_413), .A2(n_482), .B(n_484), .C(n_487), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_416), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_427), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g471 ( .A(n_427), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_437), .C(n_446), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_435), .A2(n_445), .B1(n_509), .B2(n_510), .C(n_512), .Y(n_508) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_441), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_448), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_SL g509 ( .A(n_448), .Y(n_509) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NOR4xp25_ASAP7_75t_L g451 ( .A(n_452), .B(n_481), .C(n_501), .D(n_508), .Y(n_451) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_457), .B(n_459), .C(n_477), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B(n_465), .C(n_469), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g488 ( .A(n_466), .Y(n_488) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
OR2x2_ASAP7_75t_L g499 ( .A(n_467), .B(n_500), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_491), .B2(n_493), .C(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_498), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI322xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .A3(n_529), .B1(n_531), .B2(n_534), .C1(n_535), .C2(n_537), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
endmodule