module fake_netlist_6_2303_n_1596 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1596);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1596;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_47),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_1),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_37),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_56),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_44),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_98),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_84),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_128),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_115),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_38),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_102),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_7),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_17),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_29),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_99),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_45),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_41),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_12),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_20),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_34),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_25),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_33),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_72),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_63),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_38),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_68),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_80),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_85),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_88),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_140),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_40),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_104),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_73),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_51),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_13),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_97),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_122),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_114),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_67),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_37),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_49),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_22),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_59),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_109),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_44),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_113),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_30),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_91),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_43),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_21),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_9),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_126),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_14),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_48),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_137),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_54),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_141),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_41),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_0),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_28),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_52),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_110),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_61),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_240),
.B(n_0),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_149),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_173),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_180),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_164),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_175),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_167),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_182),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_194),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_194),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_183),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_194),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_201),
.B(n_2),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_171),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_153),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_188),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_206),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_207),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_201),
.B(n_2),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_R g338 ( 
.A(n_159),
.B(n_161),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_209),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_165),
.B(n_3),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_187),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_199),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_220),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_222),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_227),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_232),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_213),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_181),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_255),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_300),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_280),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_269),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_184),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_234),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_203),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_241),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_238),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_239),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_212),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_269),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_219),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_237),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_250),
.B(n_4),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_260),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_243),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_246),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_251),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_284),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_304),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_153),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_313),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_170),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_306),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_363),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_316),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_307),
.A2(n_252),
.B(n_170),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_309),
.B(n_252),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_150),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_312),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_312),
.A2(n_155),
.B(n_151),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_325),
.B(n_159),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_314),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_337),
.B(n_161),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_310),
.Y(n_411)
);

AND3x1_ASAP7_75t_L g412 ( 
.A(n_302),
.B(n_176),
.C(n_168),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_318),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_322),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_177),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_327),
.B(n_166),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_166),
.Y(n_422)
);

OA21x2_ASAP7_75t_L g423 ( 
.A1(n_361),
.A2(n_179),
.B(n_178),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_358),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_373),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_332),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_331),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_365),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_334),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_362),
.B(n_202),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_331),
.A2(n_189),
.B(n_185),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_344),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_335),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_391),
.B(n_336),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_367),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_385),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_385),
.B(n_400),
.Y(n_449)
);

INVx4_ASAP7_75t_SL g450 ( 
.A(n_402),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_315),
.Y(n_451)
);

CKINVDCx6p67_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_339),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_391),
.B(n_158),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_343),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_403),
.Y(n_458)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_412),
.B(n_154),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_346),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_347),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_340),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_412),
.B(n_154),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_407),
.B(n_348),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_407),
.B(n_349),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_345),
.C(n_366),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_396),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_410),
.B(n_359),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_403),
.B(n_154),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_410),
.B(n_364),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_403),
.B(n_372),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_419),
.B(n_374),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_429),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_375),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_368),
.Y(n_482)
);

BUFx4f_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_426),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_422),
.B(n_371),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_404),
.B(n_231),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_402),
.B(n_154),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_426),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_429),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_417),
.B(n_371),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_233),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_381),
.B(n_376),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_390),
.A2(n_283),
.B1(n_226),
.B2(n_215),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_423),
.B(n_154),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_384),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_414),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_393),
.A2(n_256),
.B1(n_224),
.B2(n_223),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_408),
.B(n_162),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_411),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_413),
.B(n_377),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_415),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_392),
.B(n_420),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx4_ASAP7_75t_SL g514 ( 
.A(n_402),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_408),
.B(n_263),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_392),
.B(n_376),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_399),
.A2(n_369),
.B1(n_377),
.B2(n_162),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_408),
.B(n_264),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_272),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_392),
.B(n_157),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_427),
.B(n_333),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_397),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_430),
.A2(n_354),
.B1(n_353),
.B2(n_351),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_409),
.B(n_275),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_427),
.B(n_156),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_431),
.B(n_195),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_402),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_431),
.B(n_200),
.Y(n_533)
);

INVx4_ASAP7_75t_SL g534 ( 
.A(n_409),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_409),
.B(n_162),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_432),
.B(n_210),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_L g538 ( 
.A1(n_435),
.A2(n_285),
.B1(n_160),
.B2(n_157),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_433),
.B(n_162),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_379),
.B(n_214),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_438),
.B(n_204),
.C(n_208),
.Y(n_544)
);

BUFx4f_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_399),
.A2(n_162),
.B1(n_192),
.B2(n_262),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_397),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_380),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_436),
.B(n_174),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_436),
.B(n_228),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_399),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_380),
.B(n_235),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_382),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_399),
.A2(n_192),
.B1(n_257),
.B2(n_271),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_382),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_406),
.B(n_245),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_434),
.B(n_274),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_406),
.A2(n_192),
.B1(n_278),
.B2(n_291),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_386),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_406),
.B(n_248),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_388),
.B(n_389),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_388),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_401),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_477),
.B(n_519),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_530),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_446),
.B(n_350),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_477),
.B(n_401),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_L g576 ( 
.A(n_446),
.B(n_287),
.C(n_258),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_519),
.B(n_448),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_497),
.B(n_169),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_508),
.B(n_389),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_532),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_453),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_467),
.B(n_398),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_459),
.A2(n_441),
.B1(n_192),
.B2(n_286),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_L g586 ( 
.A(n_456),
.B(n_169),
.C(n_172),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_398),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_497),
.B(n_172),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_512),
.B(n_434),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_458),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_474),
.B(n_418),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_509),
.B(n_225),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_479),
.B(n_225),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_449),
.B(n_428),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_485),
.B(n_428),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_455),
.B(n_418),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_485),
.B(n_445),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_483),
.A2(n_441),
.B(n_428),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_505),
.B(n_274),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_457),
.B(n_442),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_547),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_456),
.B(n_292),
.C(n_293),
.Y(n_603)
);

INVx8_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

BUFx6f_ASAP7_75t_SL g605 ( 
.A(n_501),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_459),
.A2(n_441),
.B1(n_192),
.B2(n_286),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_479),
.B(n_292),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_452),
.B(n_160),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_SL g610 ( 
.A(n_466),
.B(n_299),
.C(n_301),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_505),
.A2(n_394),
.B(n_434),
.C(n_443),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_549),
.A2(n_163),
.B1(n_236),
.B2(n_294),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_460),
.B(n_293),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_466),
.A2(n_442),
.B(n_301),
.C(n_299),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_478),
.A2(n_247),
.B1(n_186),
.B2(n_190),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_461),
.B(n_549),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_470),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_473),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_540),
.B(n_191),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_540),
.B(n_193),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_522),
.B(n_544),
.C(n_538),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_488),
.A2(n_512),
.B1(n_447),
.B2(n_465),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_L g626 ( 
.A1(n_465),
.A2(n_298),
.B1(n_297),
.B2(n_295),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_L g627 ( 
.A(n_522),
.B(n_254),
.C(n_197),
.Y(n_627)
);

AND2x4_ASAP7_75t_SL g628 ( 
.A(n_501),
.B(n_202),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_571),
.B(n_205),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_511),
.B(n_55),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_447),
.B(n_202),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_547),
.B(n_274),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_564),
.Y(n_635)
);

BUFx8_ASAP7_75t_L g636 ( 
.A(n_526),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_537),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_484),
.B(n_163),
.Y(n_639)
);

BUFx8_ASAP7_75t_L g640 ( 
.A(n_548),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_525),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_527),
.B(n_57),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_504),
.B(n_211),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_547),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_546),
.B(n_217),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_570),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_546),
.B(n_218),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_555),
.B(n_541),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_492),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_447),
.B(n_221),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_555),
.B(n_541),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_565),
.A2(n_298),
.B1(n_297),
.B2(n_295),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_492),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_516),
.B(n_268),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_267),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_551),
.B(n_273),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_482),
.B(n_261),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_566),
.B(n_4),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_565),
.A2(n_294),
.B1(n_236),
.B2(n_288),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_541),
.B(n_289),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_516),
.A2(n_493),
.B1(n_535),
.B2(n_513),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_517),
.B(n_281),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_537),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_558),
.A2(n_279),
.B1(n_277),
.B2(n_276),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_541),
.B(n_259),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_518),
.B(n_524),
.Y(n_667)
);

INVx8_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_553),
.B(n_253),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_516),
.B(n_244),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g671 ( 
.A(n_481),
.B(n_242),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_451),
.B(n_230),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_554),
.B(n_5),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_451),
.B(n_10),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_558),
.B(n_58),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_559),
.B(n_12),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_486),
.B(n_15),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_500),
.B(n_539),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_525),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_496),
.B(n_18),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_65),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_561),
.B(n_21),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_569),
.B(n_70),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_451),
.Y(n_685)
);

BUFx12f_ASAP7_75t_SL g686 ( 
.A(n_531),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_531),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_561),
.B(n_136),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_472),
.B(n_26),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_560),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_26),
.C(n_27),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_561),
.B(n_71),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_560),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_563),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_531),
.A2(n_129),
.B1(n_124),
.B2(n_123),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_536),
.B(n_111),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_543),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_533),
.B(n_34),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_510),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_533),
.B(n_35),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_498),
.B(n_35),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_533),
.B(n_39),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_552),
.B(n_39),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_552),
.A2(n_568),
.B1(n_562),
.B2(n_515),
.Y(n_704)
);

BUFx6f_ASAP7_75t_SL g705 ( 
.A(n_563),
.Y(n_705)
);

AND2x4_ASAP7_75t_SL g706 ( 
.A(n_552),
.B(n_103),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_SL g707 ( 
.A(n_454),
.B(n_42),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_562),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_556),
.B(n_48),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_562),
.A2(n_75),
.B1(n_82),
.B2(n_49),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_619),
.B(n_545),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_652),
.A2(n_499),
.B(n_523),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_572),
.B(n_550),
.Y(n_714)
);

AOI21x1_ASAP7_75t_L g715 ( 
.A1(n_599),
.A2(n_520),
.B(n_521),
.Y(n_715)
);

NOR2x1_ASAP7_75t_L g716 ( 
.A(n_602),
.B(n_528),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_585),
.A2(n_568),
.B1(n_567),
.B2(n_557),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_622),
.A2(n_568),
.B(n_476),
.C(n_557),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_634),
.B(n_567),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_578),
.A2(n_487),
.B(n_476),
.C(n_550),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_678),
.A2(n_494),
.B(n_503),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_598),
.B(n_542),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_613),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_641),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_635),
.B(n_542),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_638),
.B(n_487),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_589),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_575),
.A2(n_599),
.B(n_595),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_585),
.A2(n_495),
.B1(n_490),
.B2(n_462),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_635),
.A2(n_475),
.B1(n_469),
.B2(n_463),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_621),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_596),
.A2(n_692),
.B(n_688),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_573),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_577),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_613),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_667),
.B(n_502),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_502),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_634),
.B(n_502),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_681),
.B(n_454),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_641),
.B(n_450),
.Y(n_740)
);

AOI21x1_ASAP7_75t_L g741 ( 
.A1(n_661),
.A2(n_666),
.B(n_656),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_607),
.A2(n_463),
.B1(n_491),
.B2(n_489),
.Y(n_742)
);

AO21x1_ASAP7_75t_L g743 ( 
.A1(n_683),
.A2(n_507),
.B(n_450),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_625),
.A2(n_463),
.B1(n_491),
.B2(n_489),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_574),
.B(n_463),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_683),
.A2(n_507),
.B(n_536),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_607),
.A2(n_491),
.B1(n_489),
.B2(n_506),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_450),
.B(n_514),
.C(n_536),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_675),
.A2(n_506),
.B(n_514),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_611),
.A2(n_536),
.B(n_506),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_579),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_583),
.B(n_514),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_600),
.B(n_534),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_613),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_646),
.A2(n_536),
.B(n_534),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_657),
.B(n_662),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_645),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_687),
.B(n_658),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_576),
.A2(n_624),
.B1(n_610),
.B2(n_644),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_629),
.B(n_623),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_684),
.A2(n_693),
.B(n_690),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_616),
.B(n_590),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_648),
.A2(n_615),
.B(n_624),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_SL g766 ( 
.A(n_605),
.B(n_705),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_699),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_576),
.A2(n_698),
.B(n_680),
.C(n_677),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_616),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_639),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_620),
.B(n_616),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_663),
.B(n_630),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_647),
.B(n_581),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_671),
.B(n_626),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_702),
.B(n_594),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_664),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_606),
.B(n_608),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_606),
.B(n_584),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_676),
.B(n_580),
.Y(n_779)
);

CKINVDCx10_ASAP7_75t_R g780 ( 
.A(n_605),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_593),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_653),
.A2(n_660),
.B(n_588),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_700),
.A2(n_654),
.B(n_642),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_618),
.A2(n_650),
.B(n_669),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_686),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_696),
.A2(n_632),
.B(n_651),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_685),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_655),
.A2(n_670),
.B(n_592),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_614),
.A2(n_631),
.B(n_706),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_L g790 ( 
.A1(n_597),
.A2(n_587),
.B(n_601),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_626),
.B(n_643),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_676),
.B(n_700),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_653),
.A2(n_660),
.B1(n_710),
.B2(n_708),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_591),
.B(n_689),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_703),
.A2(n_673),
.B(n_603),
.C(n_586),
.Y(n_796)
);

OAI21xp33_ASAP7_75t_L g797 ( 
.A1(n_617),
.A2(n_665),
.B(n_612),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_637),
.B(n_627),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_637),
.A2(n_695),
.B(n_664),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_664),
.A2(n_668),
.B(n_604),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_707),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_668),
.A2(n_604),
.B(n_627),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_633),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_633),
.B(n_628),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_586),
.A2(n_603),
.B(n_633),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_609),
.B(n_674),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_674),
.A2(n_697),
.B(n_612),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_674),
.A2(n_697),
.B(n_659),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_659),
.A2(n_708),
.B(n_691),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_659),
.Y(n_810)
);

AOI21x1_ASAP7_75t_L g811 ( 
.A1(n_701),
.A2(n_691),
.B(n_705),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_636),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_694),
.B(n_701),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_701),
.A2(n_640),
.B(n_483),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_640),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_R g817 ( 
.A(n_694),
.B(n_397),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_613),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_649),
.A2(n_652),
.B(n_678),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_619),
.B(n_641),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_649),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_572),
.B(n_619),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_572),
.B(n_619),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_641),
.Y(n_828)
);

CKINVDCx10_ASAP7_75t_R g829 ( 
.A(n_605),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_572),
.A2(n_578),
.B(n_466),
.C(n_598),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_641),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_589),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_574),
.B(n_498),
.C(n_479),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_619),
.B(n_391),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_572),
.A2(n_619),
.B(n_477),
.C(n_622),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_589),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_664),
.B(n_668),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_599),
.A2(n_692),
.B(n_688),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_649),
.A2(n_652),
.B(n_678),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_649),
.A2(n_652),
.B(n_678),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_599),
.A2(n_692),
.B(n_688),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_572),
.B(n_619),
.Y(n_843)
);

AOI21xp33_ASAP7_75t_L g844 ( 
.A1(n_644),
.A2(n_391),
.B(n_477),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_572),
.A2(n_578),
.B(n_466),
.C(n_598),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_619),
.B(n_391),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_613),
.B(n_616),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_572),
.A2(n_619),
.B1(n_477),
.B2(n_635),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_574),
.B(n_498),
.C(n_479),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_599),
.A2(n_692),
.B(n_688),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_599),
.A2(n_692),
.B(n_688),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_572),
.A2(n_678),
.B1(n_578),
.B2(n_704),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_619),
.B(n_391),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_572),
.A2(n_619),
.B1(n_477),
.B2(n_635),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_572),
.A2(n_578),
.B(n_466),
.C(n_598),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_583),
.B(n_391),
.Y(n_860)
);

AOI21xp33_ASAP7_75t_L g861 ( 
.A1(n_644),
.A2(n_391),
.B(n_477),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_602),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_649),
.A2(n_545),
.B(n_483),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_572),
.A2(n_578),
.B(n_466),
.C(n_598),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_634),
.B(n_391),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_589),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_572),
.B(n_619),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_602),
.B(n_645),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_L g869 ( 
.A(n_638),
.B(n_508),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_649),
.A2(n_652),
.B(n_678),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_641),
.Y(n_871)
);

CKINVDCx8_ASAP7_75t_R g872 ( 
.A(n_780),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_835),
.B(n_847),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_834),
.A2(n_850),
.B1(n_844),
.B2(n_861),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_759),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_856),
.B(n_826),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_763),
.A2(n_713),
.B(n_784),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_733),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_794),
.A2(n_761),
.B1(n_793),
.B2(n_712),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_827),
.B(n_843),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_790),
.B(n_778),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_765),
.A2(n_792),
.B(n_831),
.Y(n_882)
);

AND3x4_ASAP7_75t_L g883 ( 
.A(n_806),
.B(n_798),
.C(n_868),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_867),
.B(n_849),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_854),
.A2(n_728),
.B(n_820),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_836),
.B(n_722),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_820),
.A2(n_841),
.B(n_840),
.Y(n_887)
);

AND2x2_ASAP7_75t_SL g888 ( 
.A(n_803),
.B(n_815),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_857),
.B(n_758),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_762),
.B(n_845),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_734),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_782),
.A2(n_797),
.B(n_768),
.C(n_859),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_840),
.A2(n_870),
.B(n_841),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_779),
.B(n_824),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_745),
.B(n_719),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_772),
.B(n_725),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_870),
.A2(n_864),
.B(n_765),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_776),
.B(n_838),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_860),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_SL g900 ( 
.A1(n_717),
.A2(n_718),
.B(n_742),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_724),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_711),
.A2(n_818),
.B(n_816),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_731),
.B(n_760),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_822),
.A2(n_825),
.B(n_863),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_775),
.B(n_777),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_823),
.A2(n_852),
.B(n_830),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_738),
.B(n_833),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_723),
.B(n_724),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_846),
.A2(n_858),
.B(n_855),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_866),
.B(n_821),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_751),
.Y(n_911)
);

OAI21x1_ASAP7_75t_SL g912 ( 
.A1(n_786),
.A2(n_789),
.B(n_799),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_753),
.B(n_727),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_837),
.B(n_714),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_809),
.B(n_788),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_770),
.A2(n_774),
.B(n_754),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_770),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_756),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_791),
.A2(n_807),
.B1(n_796),
.B2(n_717),
.Y(n_919)
);

BUFx2_ASAP7_75t_SL g920 ( 
.A(n_869),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_721),
.A2(n_720),
.B(n_746),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_808),
.A2(n_742),
.B1(n_746),
.B2(n_805),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_817),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_767),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_SL g925 ( 
.A(n_723),
.B(n_724),
.Y(n_925)
);

OA22x2_ASAP7_75t_L g926 ( 
.A1(n_810),
.A2(n_795),
.B1(n_806),
.B2(n_798),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_787),
.B(n_773),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_721),
.A2(n_729),
.B(n_757),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_773),
.B(n_862),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_764),
.B(n_819),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_764),
.B(n_819),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_748),
.A2(n_783),
.B(n_757),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_736),
.B(n_755),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_783),
.A2(n_750),
.B(n_749),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_755),
.B(n_771),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_804),
.B(n_811),
.Y(n_936)
);

AOI221x1_ASAP7_75t_L g937 ( 
.A1(n_801),
.A2(n_729),
.B1(n_802),
.B2(n_730),
.C(n_744),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_781),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_747),
.A2(n_842),
.B(n_853),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_716),
.B(n_752),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_776),
.B(n_838),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_723),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_747),
.A2(n_737),
.B(n_739),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_828),
.B(n_871),
.Y(n_944)
);

OAI21x1_ASAP7_75t_SL g945 ( 
.A1(n_743),
.A2(n_814),
.B(n_750),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_813),
.B(n_785),
.C(n_803),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_839),
.A2(n_851),
.B(n_740),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_871),
.A2(n_832),
.B1(n_828),
.B2(n_723),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_848),
.A2(n_871),
.B(n_832),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_726),
.A2(n_832),
.B(n_828),
.C(n_803),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_838),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_735),
.B(n_769),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_766),
.A2(n_812),
.B(n_769),
.C(n_815),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_815),
.B(n_829),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_849),
.B(n_857),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_865),
.B(n_634),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_844),
.A2(n_861),
.B(n_790),
.C(n_836),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_815),
.Y(n_958)
);

OA21x2_ASAP7_75t_L g959 ( 
.A1(n_721),
.A2(n_732),
.B(n_728),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_835),
.B(n_847),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_834),
.A2(n_850),
.B1(n_861),
.B2(n_844),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_860),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_849),
.B(n_857),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_865),
.B(n_634),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_753),
.B(n_801),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_847),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_835),
.B(n_847),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_731),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_728),
.A2(n_652),
.B(n_649),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_731),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_793),
.A2(n_572),
.B1(n_761),
.B2(n_836),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_844),
.A2(n_861),
.B(n_790),
.C(n_836),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_741),
.A2(n_715),
.B(n_714),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_728),
.A2(n_652),
.B(n_649),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_776),
.B(n_868),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_827),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_724),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_800),
.B(n_838),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_860),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_815),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_826),
.B(n_827),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_835),
.B(n_847),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_854),
.A2(n_728),
.B(n_820),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_844),
.A2(n_861),
.B(n_782),
.C(n_836),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_844),
.A2(n_861),
.B(n_782),
.C(n_836),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_849),
.B(n_857),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_835),
.B(n_847),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_733),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_SL g989 ( 
.A1(n_717),
.A2(n_572),
.B(n_718),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_835),
.B(n_847),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_815),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_844),
.A2(n_861),
.B(n_782),
.C(n_836),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_793),
.A2(n_572),
.B1(n_761),
.B2(n_836),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_728),
.A2(n_652),
.B(n_649),
.Y(n_994)
);

INVx6_ASAP7_75t_L g995 ( 
.A(n_815),
.Y(n_995)
);

INVx3_ASAP7_75t_SL g996 ( 
.A(n_815),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_976),
.B(n_981),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_901),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_873),
.A2(n_967),
.B(n_987),
.C(n_966),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_956),
.B(n_964),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_898),
.B(n_941),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_890),
.A2(n_915),
.B(n_989),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_881),
.B(n_962),
.Y(n_1003)
);

AOI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_960),
.A2(n_990),
.B(n_982),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_876),
.B(n_905),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_898),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_879),
.A2(n_961),
.B1(n_874),
.B2(n_979),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_941),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_975),
.B(n_978),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_955),
.A2(n_963),
.B1(n_986),
.B2(n_993),
.Y(n_1010)
);

INVx8_ASAP7_75t_L g1011 ( 
.A(n_991),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_962),
.B(n_979),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_978),
.B(n_926),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_872),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_896),
.B(n_880),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_924),
.Y(n_1016)
);

CKINVDCx16_ASAP7_75t_R g1017 ( 
.A(n_923),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_891),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_971),
.A2(n_993),
.B1(n_889),
.B2(n_919),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_911),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_969),
.A2(n_994),
.B(n_974),
.Y(n_1021)
);

AO21x2_ASAP7_75t_L g1022 ( 
.A1(n_939),
.A2(n_921),
.B(n_885),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_888),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_L g1024 ( 
.A(n_972),
.B(n_957),
.C(n_971),
.Y(n_1024)
);

CKINVDCx6p67_ASAP7_75t_R g1025 ( 
.A(n_996),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_927),
.B(n_976),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_899),
.B(n_929),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_900),
.A2(n_983),
.B(n_885),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_917),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_981),
.B(n_918),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_884),
.B(n_895),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_988),
.B(n_968),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_938),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_926),
.B(n_970),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_894),
.B(n_914),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_975),
.B(n_978),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_958),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_958),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_920),
.B(n_908),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_903),
.Y(n_1040)
);

NAND2x1_ASAP7_75t_L g1041 ( 
.A(n_925),
.B(n_912),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_951),
.B(n_946),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_983),
.A2(n_886),
.B(n_909),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_886),
.A2(n_959),
.B(n_902),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_892),
.B(n_984),
.Y(n_1045)
);

INVx3_ASAP7_75t_SL g1046 ( 
.A(n_995),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_901),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_916),
.B(n_936),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_985),
.A2(n_992),
.B1(n_919),
.B2(n_928),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_980),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_930),
.B(n_931),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_935),
.B(n_910),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_901),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_951),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_933),
.Y(n_1055)
);

NAND2x1_ASAP7_75t_L g1056 ( 
.A(n_965),
.B(n_977),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_977),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_897),
.A2(n_922),
.B(n_921),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_953),
.B(n_950),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_883),
.B(n_922),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_882),
.B(n_897),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_944),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_954),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_934),
.A2(n_932),
.B(n_947),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_943),
.A2(n_887),
.B(n_893),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_SL g1066 ( 
.A1(n_937),
.A2(n_948),
.B(n_893),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_907),
.B(n_913),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_940),
.B(n_952),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_977),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_965),
.B(n_949),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_945),
.A2(n_947),
.B(n_948),
.C(n_942),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_942),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_965),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_973),
.B(n_965),
.C(n_906),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_904),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_877),
.A2(n_741),
.B(n_715),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_875),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_976),
.B(n_981),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_881),
.B(n_790),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_923),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_901),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_878),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_978),
.B(n_800),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_890),
.A2(n_732),
.B(n_915),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_924),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_957),
.A2(n_861),
.B(n_844),
.C(n_879),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_898),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_881),
.A2(n_850),
.B1(n_834),
.B2(n_844),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_962),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_978),
.B(n_800),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_976),
.B(n_981),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_898),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_898),
.B(n_941),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_976),
.B(n_981),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_957),
.A2(n_861),
.B(n_844),
.C(n_879),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_873),
.A2(n_966),
.B(n_960),
.Y(n_1096)
);

CKINVDCx6p67_ASAP7_75t_R g1097 ( 
.A(n_996),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_875),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_971),
.A2(n_993),
.B(n_972),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_956),
.B(n_964),
.Y(n_1100)
);

AND2x6_ASAP7_75t_L g1101 ( 
.A(n_915),
.B(n_879),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_SL g1102 ( 
.A1(n_957),
.A2(n_574),
.B(n_587),
.C(n_584),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_956),
.B(n_964),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_971),
.A2(n_993),
.B(n_972),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_901),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_956),
.B(n_964),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_876),
.B(n_881),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_878),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_924),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_976),
.B(n_981),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_879),
.A2(n_873),
.B1(n_966),
.B2(n_960),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_976),
.B(n_981),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_901),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1055),
.B(n_1010),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1047),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1016),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_1013),
.B(n_1083),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1020),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1089),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_1071),
.A2(n_1070),
.B(n_1035),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1047),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1079),
.A2(n_1060),
.B1(n_1088),
.B2(n_1111),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1085),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_997),
.B(n_1078),
.Y(n_1124)
);

BUFx4_ASAP7_75t_SL g1125 ( 
.A(n_1050),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1005),
.B(n_1107),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1109),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1111),
.A2(n_1007),
.B1(n_1096),
.B2(n_1060),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1018),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1012),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1013),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1089),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_1078),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_1043),
.A2(n_1002),
.B(n_1044),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1080),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1049),
.A2(n_1045),
.B(n_1028),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1096),
.B(n_999),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1046),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_L g1139 ( 
.A(n_1001),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1091),
.B(n_1094),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1029),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1077),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1003),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_1059),
.B(n_1009),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1076),
.A2(n_1021),
.B(n_1084),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1082),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_SL g1148 ( 
.A1(n_1049),
.A2(n_1099),
.B1(n_1104),
.B2(n_1101),
.Y(n_1148)
);

INVx6_ASAP7_75t_SL g1149 ( 
.A(n_1039),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1004),
.B(n_1026),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1004),
.B(n_1015),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1063),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1091),
.A2(n_1094),
.B1(n_1110),
.B2(n_1112),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1032),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1024),
.A2(n_1095),
.B(n_1086),
.Y(n_1155)
);

INVx4_ASAP7_75t_SL g1156 ( 
.A(n_1101),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1101),
.A2(n_1019),
.B1(n_1104),
.B2(n_1099),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1013),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1110),
.B(n_1112),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1047),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_1101),
.A2(n_1058),
.B1(n_1048),
.B2(n_1059),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1072),
.Y(n_1162)
);

BUFx4_ASAP7_75t_R g1163 ( 
.A(n_1054),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1056),
.B(n_1009),
.Y(n_1164)
);

BUFx4f_ASAP7_75t_SL g1165 ( 
.A(n_1025),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1036),
.B(n_1073),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1108),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1097),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1033),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1098),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1037),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1031),
.A2(n_1068),
.B1(n_1106),
.B2(n_1103),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1062),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1000),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1030),
.B(n_1100),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1023),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1036),
.A2(n_1034),
.B1(n_1042),
.B2(n_1011),
.Y(n_1177)
);

CKINVDCx10_ASAP7_75t_R g1178 ( 
.A(n_1017),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1040),
.A2(n_1051),
.B1(n_1042),
.B2(n_1067),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1083),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1064),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1038),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1001),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_1011),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1052),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1022),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1102),
.B(n_1087),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1074),
.A2(n_1061),
.B(n_1065),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1011),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1006),
.B(n_1008),
.Y(n_1191)
);

BUFx2_ASAP7_75t_R g1192 ( 
.A(n_1070),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1090),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1093),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_998),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_998),
.Y(n_1196)
);

INVx5_ASAP7_75t_L g1197 ( 
.A(n_998),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1022),
.B(n_1066),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_1053),
.B(n_1057),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_1113),
.A2(n_1053),
.B(n_1057),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1069),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1069),
.A2(n_1081),
.B(n_1105),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1105),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1012),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1016),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1016),
.Y(n_1206)
);

BUFx2_ASAP7_75t_R g1207 ( 
.A(n_1014),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1005),
.B(n_1107),
.Y(n_1208)
);

AO21x1_ASAP7_75t_L g1209 ( 
.A1(n_1049),
.A2(n_957),
.B(n_971),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1041),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1046),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1016),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1013),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1079),
.A2(n_834),
.B1(n_850),
.B2(n_574),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1055),
.B(n_1010),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1016),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1187),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1181),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1193),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1189),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1146),
.A2(n_1209),
.B(n_1157),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1135),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1117),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1136),
.A2(n_1134),
.B(n_1148),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1124),
.B(n_1133),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1134),
.Y(n_1226)
);

INVxp33_ASAP7_75t_L g1227 ( 
.A(n_1154),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1162),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1137),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1124),
.B(n_1133),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1117),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_1186),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1117),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1198),
.A2(n_1120),
.B(n_1188),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1198),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1155),
.B(n_1131),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1140),
.B(n_1159),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1162),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1140),
.B(n_1159),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1153),
.B(n_1186),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1180),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1136),
.B(n_1158),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1193),
.B(n_1210),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1119),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1155),
.B(n_1161),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1155),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1114),
.B(n_1215),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1131),
.B(n_1213),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1129),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1147),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1213),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1114),
.B(n_1215),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_1122),
.B(n_1151),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1150),
.B(n_1123),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1167),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1144),
.B(n_1130),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1132),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1169),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1184),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1204),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1145),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1199),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1208),
.B(n_1214),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1173),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1116),
.A2(n_1216),
.B(n_1118),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1172),
.A2(n_1179),
.B(n_1191),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1156),
.B(n_1121),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1164),
.A2(n_1166),
.B(n_1212),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1127),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1205),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1206),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1156),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1156),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1141),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1178),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1145),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1145),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1202),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1164),
.A2(n_1166),
.B(n_1200),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1145),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1229),
.B(n_1175),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1278),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1278),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1235),
.B(n_1174),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1253),
.A2(n_1152),
.B1(n_1192),
.B2(n_1139),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1222),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1235),
.B(n_1143),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1246),
.B(n_1177),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1229),
.B(n_1176),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1262),
.Y(n_1290)
);

NOR2x1_ASAP7_75t_L g1291 ( 
.A(n_1220),
.B(n_1121),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1218),
.B(n_1203),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1262),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1240),
.B(n_1195),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1263),
.B(n_1149),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1234),
.Y(n_1296)
);

OR2x2_ASAP7_75t_SL g1297 ( 
.A(n_1234),
.B(n_1163),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1245),
.B(n_1201),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1219),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1224),
.A2(n_1196),
.B(n_1149),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1240),
.B(n_1201),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1226),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1245),
.B(n_1194),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1217),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1221),
.B(n_1234),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1232),
.B(n_1115),
.Y(n_1306)
);

NAND2x1_ASAP7_75t_L g1307 ( 
.A(n_1242),
.B(n_1160),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1236),
.B(n_1115),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1221),
.B(n_1183),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1221),
.B(n_1183),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1234),
.B(n_1183),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_L g1312 ( 
.A(n_1265),
.B(n_1160),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1234),
.B(n_1183),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1263),
.A2(n_1139),
.B(n_1197),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1298),
.B(n_1247),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1285),
.A2(n_1224),
.B(n_1266),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1298),
.B(n_1247),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1295),
.A2(n_1253),
.B1(n_1231),
.B2(n_1233),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1298),
.B(n_1252),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1303),
.B(n_1252),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1289),
.A2(n_1227),
.B1(n_1260),
.B2(n_1244),
.C(n_1238),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1295),
.B(n_1253),
.C(n_1266),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1281),
.B(n_1289),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1281),
.B(n_1257),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1285),
.B(n_1253),
.C(n_1257),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1287),
.B(n_1228),
.Y(n_1326)
);

AOI211xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1311),
.A2(n_1236),
.B(n_1273),
.C(n_1272),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1302),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1311),
.B(n_1313),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1314),
.A2(n_1288),
.B(n_1231),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1294),
.A2(n_1260),
.B1(n_1238),
.B2(n_1274),
.C(n_1254),
.Y(n_1331)
);

OAI221xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1296),
.A2(n_1248),
.B1(n_1242),
.B2(n_1256),
.C(n_1251),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1287),
.B(n_1254),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1287),
.B(n_1232),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1314),
.A2(n_1253),
.B1(n_1288),
.B2(n_1261),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1308),
.Y(n_1336)
);

NOR3xp33_ASAP7_75t_L g1337 ( 
.A(n_1294),
.B(n_1268),
.C(n_1273),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1301),
.B(n_1256),
.C(n_1271),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1284),
.B(n_1225),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1284),
.B(n_1225),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1301),
.B(n_1270),
.C(n_1269),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1306),
.B(n_1270),
.C(n_1269),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1284),
.B(n_1237),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1305),
.A2(n_1251),
.B1(n_1230),
.B2(n_1239),
.C(n_1271),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1306),
.B(n_1237),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1300),
.A2(n_1223),
.B1(n_1242),
.B2(n_1259),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1312),
.A2(n_1268),
.B(n_1279),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1312),
.B(n_1248),
.C(n_1255),
.Y(n_1348)
);

OAI221xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1296),
.A2(n_1242),
.B1(n_1230),
.B2(n_1239),
.C(n_1280),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1296),
.B(n_1255),
.C(n_1258),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1292),
.B(n_1264),
.Y(n_1351)
);

OAI221xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1305),
.A2(n_1242),
.B1(n_1280),
.B2(n_1277),
.C(n_1276),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1313),
.B(n_1241),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1305),
.A2(n_1267),
.B(n_1243),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1291),
.A2(n_1268),
.B(n_1279),
.Y(n_1355)
);

OAI211xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1308),
.A2(n_1168),
.B(n_1135),
.C(n_1249),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1291),
.B(n_1250),
.C(n_1249),
.Y(n_1357)
);

OAI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1307),
.A2(n_1211),
.B1(n_1138),
.B2(n_1272),
.C(n_1267),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1328),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1323),
.B(n_1282),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1329),
.B(n_1309),
.Y(n_1361)
);

NOR2xp67_ASAP7_75t_SL g1362 ( 
.A(n_1325),
.B(n_1219),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1328),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1336),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1351),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1329),
.B(n_1309),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1350),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1353),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1315),
.B(n_1310),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1324),
.B(n_1282),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1350),
.B(n_1283),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1315),
.B(n_1310),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1356),
.B(n_1308),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1342),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1342),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1358),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1317),
.B(n_1310),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1338),
.B(n_1283),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1341),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1338),
.B(n_1290),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1357),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1317),
.B(n_1290),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1341),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1345),
.B(n_1290),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1334),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1357),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1344),
.B(n_1304),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1347),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1326),
.B(n_1293),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1348),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1348),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1359),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1361),
.B(n_1319),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1361),
.B(n_1319),
.Y(n_1394)
);

NOR4xp75_ASAP7_75t_L g1395 ( 
.A(n_1387),
.B(n_1355),
.C(n_1307),
.D(n_1299),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1385),
.B(n_1320),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1382),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1379),
.B(n_1333),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1381),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1379),
.B(n_1339),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1376),
.B(n_1337),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1363),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1363),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1320),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1364),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1366),
.B(n_1354),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1407)
);

AOI211x1_ASAP7_75t_L g1408 ( 
.A1(n_1362),
.A2(n_1325),
.B(n_1322),
.C(n_1340),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1383),
.B(n_1343),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1364),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1366),
.B(n_1369),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_SL g1413 ( 
.A(n_1376),
.B(n_1322),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1370),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1368),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1383),
.B(n_1297),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1370),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1370),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1381),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1378),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1378),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1385),
.B(n_1321),
.Y(n_1427)
);

NOR2xp67_ASAP7_75t_L g1428 ( 
.A(n_1410),
.B(n_1391),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1405),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1411),
.Y(n_1430)
);

NAND2x1p5_ASAP7_75t_L g1431 ( 
.A(n_1413),
.B(n_1362),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1423),
.B(n_1386),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1399),
.B(n_1386),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1393),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1427),
.B(n_1376),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1393),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1414),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1394),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1414),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1412),
.B(n_1372),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1404),
.B(n_1372),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1398),
.B(n_1387),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1419),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1417),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1389),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1401),
.A2(n_1316),
.B(n_1390),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1419),
.B(n_1391),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1400),
.B(n_1389),
.Y(n_1448)
);

NAND3xp33_ASAP7_75t_L g1449 ( 
.A(n_1413),
.B(n_1362),
.C(n_1388),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1417),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1420),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1404),
.B(n_1377),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1397),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1400),
.B(n_1389),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1409),
.B(n_1384),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_SL g1457 ( 
.A(n_1410),
.B(n_1388),
.C(n_1373),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1409),
.B(n_1384),
.Y(n_1458)
);

OAI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1401),
.A2(n_1390),
.B(n_1330),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1422),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1422),
.B(n_1367),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1412),
.B(n_1377),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1401),
.B(n_1365),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1395),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1416),
.B(n_1332),
.Y(n_1465)
);

OAI21xp33_ASAP7_75t_L g1466 ( 
.A1(n_1416),
.A2(n_1330),
.B(n_1373),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1443),
.B(n_1424),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1443),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1460),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1454),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1460),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1428),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1435),
.B(n_1275),
.Y(n_1473)
);

NAND2xp33_ASAP7_75t_L g1474 ( 
.A(n_1459),
.B(n_1367),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1429),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1424),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1433),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1431),
.A2(n_1403),
.B(n_1402),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1430),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1433),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1466),
.A2(n_1318),
.B1(n_1407),
.B2(n_1418),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1431),
.B(n_1440),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1406),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1462),
.B(n_1406),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1464),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1439),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1464),
.B(n_1407),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1444),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1425),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1450),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1451),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1425),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1461),
.B(n_1432),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1449),
.B(n_1426),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_1465),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1434),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1497),
.A2(n_1408),
.B1(n_1446),
.B2(n_1432),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1487),
.B(n_1436),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1475),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1497),
.A2(n_1465),
.B1(n_1457),
.B2(n_1463),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1475),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1474),
.A2(n_1442),
.B(n_1286),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1487),
.A2(n_1438),
.B1(n_1418),
.B2(n_1455),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1472),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1472),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

AOI321xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1477),
.A2(n_1445),
.A3(n_1448),
.B1(n_1456),
.B2(n_1458),
.C(n_1397),
.Y(n_1510)
);

AOI22x1_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_1190),
.B1(n_1182),
.B2(n_1171),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1481),
.A2(n_1331),
.B(n_1378),
.C(n_1327),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1487),
.A2(n_1452),
.B1(n_1441),
.B2(n_1286),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1479),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1479),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1495),
.B(n_1396),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1495),
.B(n_1426),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1471),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1471),
.B(n_1346),
.C(n_1349),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1394),
.Y(n_1521)
);

OAI31xp33_ASAP7_75t_L g1522 ( 
.A1(n_1481),
.A2(n_1371),
.A3(n_1380),
.B(n_1352),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1480),
.A2(n_1360),
.B1(n_1415),
.B2(n_1421),
.C(n_1392),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1513),
.B(n_1473),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1507),
.B(n_1489),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1499),
.A2(n_1489),
.B1(n_1496),
.B2(n_1482),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1508),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1468),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1514),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1514),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1502),
.A2(n_1480),
.B1(n_1469),
.B2(n_1496),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1521),
.B(n_1505),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1505),
.A2(n_1470),
.B1(n_1496),
.B2(n_1486),
.Y(n_1535)
);

NAND2x1_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1482),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1511),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1518),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1517),
.B(n_1470),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1506),
.B(n_1470),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1533),
.A2(n_1512),
.B1(n_1520),
.B2(n_1496),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_SL g1544 ( 
.A(n_1526),
.B(n_1535),
.C(n_1542),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1528),
.A2(n_1522),
.B(n_1494),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1525),
.A2(n_1510),
.B(n_1516),
.C(n_1515),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1532),
.A2(n_1211),
.B(n_1138),
.Y(n_1548)
);

OAI21xp33_ASAP7_75t_L g1549 ( 
.A1(n_1535),
.A2(n_1496),
.B(n_1482),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1536),
.Y(n_1550)
);

AOI211xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1542),
.A2(n_1529),
.B(n_1531),
.C(n_1541),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1530),
.A2(n_1478),
.B(n_1483),
.Y(n_1552)
);

OAI221xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1534),
.A2(n_1523),
.B1(n_1476),
.B2(n_1491),
.C(n_1494),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1546),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1550),
.Y(n_1555)
);

NOR2xp67_ASAP7_75t_L g1556 ( 
.A(n_1552),
.B(n_1538),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1551),
.B(n_1549),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1544),
.A2(n_1524),
.B1(n_1540),
.B2(n_1486),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1545),
.B(n_1539),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1543),
.A2(n_1498),
.B1(n_1483),
.B2(n_1485),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1547),
.B(n_1537),
.C(n_1168),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1553),
.B(n_1486),
.C(n_1467),
.Y(n_1562)
);

NOR3x1_ASAP7_75t_L g1563 ( 
.A(n_1548),
.B(n_1491),
.C(n_1467),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1544),
.A2(n_1488),
.B(n_1484),
.Y(n_1564)
);

NAND4xp75_ASAP7_75t_L g1565 ( 
.A(n_1556),
.B(n_1488),
.C(n_1484),
.D(n_1490),
.Y(n_1565)
);

OAI211xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1561),
.A2(n_1476),
.B(n_1467),
.C(n_1490),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1557),
.A2(n_1493),
.B(n_1492),
.Y(n_1567)
);

NOR3xp33_ASAP7_75t_L g1568 ( 
.A(n_1559),
.B(n_1190),
.C(n_1476),
.Y(n_1568)
);

OAI211xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1558),
.A2(n_1492),
.B(n_1493),
.C(n_1498),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1554),
.B(n_1152),
.C(n_1185),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1565),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1568),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1569),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1566),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1570),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1567),
.Y(n_1576)
);

XNOR2xp5_ASAP7_75t_L g1577 ( 
.A(n_1575),
.B(n_1555),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1575),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1573),
.B(n_1564),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1574),
.B(n_1562),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1576),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1577),
.Y(n_1582)
);

INVx3_ASAP7_75t_SL g1583 ( 
.A(n_1578),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1581),
.B(n_1576),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1584),
.Y(n_1585)
);

NAND4xp25_ASAP7_75t_SL g1586 ( 
.A(n_1585),
.B(n_1579),
.C(n_1580),
.D(n_1571),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1586),
.A2(n_1582),
.B1(n_1572),
.B2(n_1583),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1586),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1587),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1588),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1590),
.A2(n_1560),
.B(n_1563),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1589),
.Y(n_1592)
);

NAND4xp25_ASAP7_75t_L g1593 ( 
.A(n_1592),
.B(n_1170),
.C(n_1142),
.D(n_1165),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1593),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_R g1595 ( 
.A1(n_1594),
.A2(n_1591),
.B1(n_1185),
.B2(n_1125),
.C(n_1207),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1595),
.A2(n_1591),
.B(n_1171),
.C(n_1142),
.Y(n_1596)
);


endmodule