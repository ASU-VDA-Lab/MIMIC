module real_aes_222_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g577 ( .A(n_0), .B(n_232), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g155 ( .A(n_2), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_3), .B(n_514), .Y(n_513) );
NAND2xp33_ASAP7_75t_SL g569 ( .A(n_4), .B(n_172), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_5), .B(n_216), .Y(n_224) );
INVx1_ASAP7_75t_L g562 ( .A(n_6), .Y(n_562) );
INVx1_ASAP7_75t_L g163 ( .A(n_7), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
AOI22xp5_ASAP7_75t_SL g121 ( .A1(n_9), .A2(n_122), .B1(n_123), .B2(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_9), .Y(n_122) );
OAI22x1_ASAP7_75t_R g124 ( .A1(n_10), .A2(n_79), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_10), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_11), .Y(n_189) );
AND2x2_ASAP7_75t_L g511 ( .A(n_12), .B(n_204), .Y(n_511) );
INVx2_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_14), .Y(n_113) );
INVx1_ASAP7_75t_L g233 ( .A(n_15), .Y(n_233) );
AOI221x1_ASAP7_75t_L g565 ( .A1(n_16), .A2(n_176), .B1(n_516), .B2(n_566), .C(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_17), .B(n_514), .Y(n_549) );
INVx1_ASAP7_75t_L g117 ( .A(n_18), .Y(n_117) );
INVx1_ASAP7_75t_L g230 ( .A(n_19), .Y(n_230) );
INVx1_ASAP7_75t_SL g245 ( .A(n_20), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_21), .B(n_166), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_22), .A2(n_30), .B1(n_502), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_22), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_23), .Y(n_837) );
AOI33xp33_ASAP7_75t_L g270 ( .A1(n_24), .A2(n_53), .A3(n_150), .B1(n_158), .B2(n_271), .B3(n_272), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_25), .A2(n_516), .B(n_517), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_26), .B(n_232), .Y(n_518) );
AOI221xp5_ASAP7_75t_SL g541 ( .A1(n_27), .A2(n_44), .B1(n_514), .B2(n_516), .C(n_542), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_28), .A2(n_104), .B1(n_119), .B2(n_814), .C1(n_816), .C2(n_839), .Y(n_103) );
OAI21xp5_ASAP7_75t_L g816 ( .A1(n_28), .A2(n_817), .B(n_832), .Y(n_816) );
INVx1_ASAP7_75t_L g835 ( .A(n_28), .Y(n_835) );
INVx1_ASAP7_75t_L g181 ( .A(n_29), .Y(n_181) );
NOR3xp33_ASAP7_75t_L g134 ( .A(n_30), .B(n_135), .C(n_326), .Y(n_134) );
INVx1_ASAP7_75t_SL g502 ( .A(n_30), .Y(n_502) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_31), .A2(n_91), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g205 ( .A(n_31), .B(n_91), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_32), .B(n_235), .Y(n_553) );
INVxp67_ASAP7_75t_L g564 ( .A(n_33), .Y(n_564) );
AND2x2_ASAP7_75t_L g537 ( .A(n_34), .B(n_203), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_35), .B(n_156), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_36), .A2(n_516), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_37), .B(n_235), .Y(n_543) );
INVx1_ASAP7_75t_L g149 ( .A(n_38), .Y(n_149) );
AND2x2_ASAP7_75t_L g161 ( .A(n_38), .B(n_152), .Y(n_161) );
AND2x2_ASAP7_75t_L g172 ( .A(n_38), .B(n_155), .Y(n_172) );
OR2x6_ASAP7_75t_L g115 ( .A(n_39), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_40), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_41), .B(n_156), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_42), .A2(n_177), .B1(n_212), .B2(n_216), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_43), .B(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_45), .A2(n_83), .B1(n_147), .B2(n_516), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_46), .B(n_166), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_47), .B(n_232), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_48), .B(n_143), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_49), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_50), .Y(n_215) );
AND2x2_ASAP7_75t_L g580 ( .A(n_51), .B(n_203), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_52), .B(n_203), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_54), .B(n_166), .Y(n_201) );
INVx1_ASAP7_75t_L g154 ( .A(n_55), .Y(n_154) );
INVx1_ASAP7_75t_L g168 ( .A(n_55), .Y(n_168) );
AND2x2_ASAP7_75t_L g202 ( .A(n_56), .B(n_203), .Y(n_202) );
AOI221xp5_ASAP7_75t_L g146 ( .A1(n_57), .A2(n_75), .B1(n_147), .B2(n_156), .C(n_162), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_58), .B(n_156), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_59), .B(n_514), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_60), .B(n_177), .Y(n_191) );
AOI21xp5_ASAP7_75t_SL g254 ( .A1(n_61), .A2(n_147), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g528 ( .A(n_62), .B(n_203), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_63), .B(n_235), .Y(n_578) );
INVx1_ASAP7_75t_L g227 ( .A(n_64), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_65), .B(n_232), .Y(n_526) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_66), .B(n_204), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_67), .A2(n_516), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g200 ( .A(n_68), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_235), .Y(n_519) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_70), .B(n_143), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_71), .A2(n_147), .B(n_199), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_72), .A2(n_121), .B1(n_806), .B2(n_810), .Y(n_805) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
INVx1_ASAP7_75t_L g170 ( .A(n_73), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_74), .B(n_156), .Y(n_273) );
AND2x2_ASAP7_75t_L g247 ( .A(n_76), .B(n_176), .Y(n_247) );
INVx1_ASAP7_75t_L g228 ( .A(n_77), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_78), .A2(n_147), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_80), .A2(n_147), .B(n_218), .C(n_222), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_81), .B(n_514), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_82), .A2(n_86), .B1(n_156), .B2(n_514), .Y(n_590) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_85), .B(n_176), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_87), .A2(n_147), .B1(n_268), .B2(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_88), .B(n_232), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_89), .B(n_232), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_90), .A2(n_516), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g256 ( .A(n_92), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_93), .B(n_235), .Y(n_525) );
AND2x2_ASAP7_75t_L g274 ( .A(n_94), .B(n_176), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_95), .A2(n_179), .B(n_180), .C(n_183), .Y(n_178) );
INVxp67_ASAP7_75t_L g567 ( .A(n_96), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_97), .B(n_514), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_98), .B(n_235), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_99), .A2(n_516), .B(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g110 ( .A(n_100), .Y(n_110) );
BUFx2_ASAP7_75t_SL g843 ( .A(n_100), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_101), .B(n_166), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g827 ( .A1(n_102), .A2(n_828), .B1(n_829), .B2(n_831), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_102), .Y(n_828) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_111), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_SL g815 ( .A(n_108), .B(n_110), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_108), .A2(n_841), .B(n_844), .Y(n_840) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g821 ( .A(n_112), .Y(n_821) );
BUFx2_ASAP7_75t_L g838 ( .A(n_112), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_SL g132 ( .A(n_113), .B(n_115), .Y(n_132) );
OR2x6_ASAP7_75t_SL g804 ( .A(n_113), .B(n_114), .Y(n_804) );
OR2x2_ASAP7_75t_L g813 ( .A(n_113), .B(n_115), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_805), .Y(n_120) );
INVxp33_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B1(n_504), .B2(n_802), .Y(n_128) );
CKINVDCx6p67_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
CKINVDCx11_ASAP7_75t_R g809 ( .A(n_130), .Y(n_809) );
INVx3_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
AOI211xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_397), .B(n_500), .C(n_503), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_134), .A2(n_397), .B(n_500), .Y(n_807) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_136), .A2(n_398), .B(n_502), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_136), .B(n_475), .Y(n_825) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_304), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_287), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_206), .B1(n_248), .B2(n_262), .C(n_277), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_193), .Y(n_139) );
NAND2x1_ASAP7_75t_SL g313 ( .A(n_140), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g340 ( .A(n_140), .B(n_310), .Y(n_340) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_140), .Y(n_386) );
AND2x2_ASAP7_75t_L g394 ( .A(n_140), .B(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g498 ( .A(n_140), .Y(n_498) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_174), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_142), .Y(n_276) );
INVx1_ASAP7_75t_L g292 ( .A(n_142), .Y(n_292) );
AND2x4_ASAP7_75t_L g299 ( .A(n_142), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g309 ( .A(n_142), .B(n_174), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_142), .B(n_295), .Y(n_336) );
INVx1_ASAP7_75t_L g347 ( .A(n_142), .Y(n_347) );
INVxp67_ASAP7_75t_L g381 ( .A(n_142), .Y(n_381) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_173), .Y(n_142) );
INVx2_ASAP7_75t_SL g222 ( .A(n_143), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_143), .A2(n_549), .B(n_550), .Y(n_548) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_145), .B(n_205), .Y(n_204) );
AND2x4_ASAP7_75t_L g216 ( .A(n_145), .B(n_205), .Y(n_216) );
INVxp67_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_147), .A2(n_156), .B1(n_561), .B2(n_563), .Y(n_560) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
NOR2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx1_ASAP7_75t_L g272 ( .A(n_150), .Y(n_272) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x6_ASAP7_75t_L g164 ( .A(n_151), .B(n_158), .Y(n_164) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g232 ( .A(n_152), .B(n_167), .Y(n_232) );
AND2x6_ASAP7_75t_L g516 ( .A(n_153), .B(n_161), .Y(n_516) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx2_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
AND2x4_ASAP7_75t_L g235 ( .A(n_154), .B(n_169), .Y(n_235) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_155), .Y(n_159) );
INVx1_ASAP7_75t_L g192 ( .A(n_156), .Y(n_192) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_160), .Y(n_156) );
INVx1_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVxp33_ASAP7_75t_L g271 ( .A(n_158), .Y(n_271) );
INVx1_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B(n_165), .C(n_171), .Y(n_162) );
INVxp67_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_164), .A2(n_171), .B(n_200), .C(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_164), .A2(n_182), .B1(n_227), .B2(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_164), .A2(n_171), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_164), .A2(n_171), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
AND2x4_ASAP7_75t_L g514 ( .A(n_166), .B(n_172), .Y(n_514) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_171), .A2(n_219), .B(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_171), .B(n_216), .Y(n_236) );
INVx1_ASAP7_75t_L g268 ( .A(n_171), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_171), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_171), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_171), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_171), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_171), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_171), .A2(n_577), .B(n_578), .Y(n_576) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_172), .Y(n_183) );
INVx2_ASAP7_75t_L g264 ( .A(n_174), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_174), .B(n_195), .Y(n_280) );
INVx1_ASAP7_75t_L g298 ( .A(n_174), .Y(n_298) );
INVx1_ASAP7_75t_L g345 ( .A(n_174), .Y(n_345) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_186), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .B1(n_184), .B2(n_185), .Y(n_175) );
INVx3_ASAP7_75t_L g185 ( .A(n_176), .Y(n_185) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_177), .B(n_188), .Y(n_187) );
AOI21x1_ASAP7_75t_L g573 ( .A1(n_177), .A2(n_574), .B(n_580), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_182), .B(n_216), .C(n_569), .Y(n_568) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_185), .A2(n_196), .B(n_202), .Y(n_195) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_185), .A2(n_196), .B(n_202), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_193), .B(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_L g334 ( .A(n_193), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_193), .B(n_299), .Y(n_353) );
INVx1_ASAP7_75t_L g362 ( .A(n_193), .Y(n_362) );
AND2x2_ASAP7_75t_L g410 ( .A(n_193), .B(n_309), .Y(n_410) );
OR2x2_ASAP7_75t_L g453 ( .A(n_193), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g293 ( .A(n_194), .B(n_294), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_194), .B(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g275 ( .A(n_195), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_195), .B(n_295), .Y(n_373) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_195), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_203), .Y(n_240) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_203), .A2(n_541), .B(n_545), .Y(n_540) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_237), .Y(n_207) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_208), .B(n_332), .Y(n_377) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g339 ( .A(n_209), .B(n_330), .Y(n_339) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_223), .Y(n_209) );
INVx1_ASAP7_75t_L g259 ( .A(n_210), .Y(n_259) );
AND2x4_ASAP7_75t_L g285 ( .A(n_210), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g289 ( .A(n_210), .Y(n_289) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_210), .Y(n_325) );
AND2x2_ASAP7_75t_L g495 ( .A(n_210), .B(n_251), .Y(n_495) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_217), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .C(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_254), .B(n_258), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_216), .A2(n_513), .B(n_515), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_216), .B(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_216), .B(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_216), .B(n_567), .Y(n_566) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_222), .A2(n_266), .B(n_274), .Y(n_265) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_222), .A2(n_266), .B(n_274), .Y(n_295) );
AOI21x1_ASAP7_75t_L g588 ( .A1(n_222), .A2(n_589), .B(n_592), .Y(n_588) );
INVx3_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
INVx2_ASAP7_75t_L g303 ( .A(n_223), .Y(n_303) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_223), .B(n_251), .Y(n_320) );
AND2x2_ASAP7_75t_L g358 ( .A(n_223), .B(n_239), .Y(n_358) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_229), .B(n_236), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B1(n_233), .B2(n_234), .Y(n_229) );
INVxp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVxp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g432 ( .A(n_237), .Y(n_432) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g261 ( .A(n_238), .Y(n_261) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
INVx1_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
INVx1_ASAP7_75t_L g390 ( .A(n_239), .Y(n_390) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_239), .Y(n_409) );
OR2x2_ASAP7_75t_L g415 ( .A(n_239), .B(n_251), .Y(n_415) );
AND2x2_ASAP7_75t_L g459 ( .A(n_239), .B(n_286), .Y(n_459) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_240), .A2(n_522), .B(n_528), .Y(n_521) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_240), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_240), .A2(n_531), .B(n_537), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_260), .Y(n_249) );
AND2x2_ASAP7_75t_L g301 ( .A(n_250), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g455 ( .A(n_250), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g460 ( .A(n_250), .Y(n_460) );
AND2x2_ASAP7_75t_L g472 ( .A(n_250), .B(n_358), .Y(n_472) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
INVx4_ASAP7_75t_L g283 ( .A(n_251), .Y(n_283) );
INVx2_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_251), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_251), .B(n_391), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_251), .B(n_261), .Y(n_464) );
AND2x2_ASAP7_75t_L g490 ( .A(n_251), .B(n_303), .Y(n_490) );
OR2x6_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x4_ASAP7_75t_L g392 ( .A(n_259), .B(n_283), .Y(n_392) );
AND2x2_ASAP7_75t_L g319 ( .A(n_260), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g337 ( .A(n_260), .B(n_324), .Y(n_337) );
INVx1_ASAP7_75t_L g371 ( .A(n_260), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_260), .B(n_285), .Y(n_427) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_261), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_262), .A2(n_344), .B1(n_488), .B2(n_491), .Y(n_487) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_275), .Y(n_262) );
INVx1_ASAP7_75t_L g417 ( .A(n_263), .Y(n_417) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_264), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g440 ( .A(n_264), .B(n_312), .Y(n_440) );
NOR2xp67_ASAP7_75t_L g449 ( .A(n_264), .B(n_312), .Y(n_449) );
INVx2_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
AND2x4_ASAP7_75t_L g310 ( .A(n_265), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_276), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_279), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g384 ( .A(n_279), .B(n_299), .Y(n_384) );
INVx2_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g422 ( .A(n_280), .B(n_336), .Y(n_422) );
INVxp33_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g403 ( .A(n_282), .Y(n_403) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x4_ASAP7_75t_SL g324 ( .A(n_283), .B(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_283), .Y(n_349) );
INVx2_ASAP7_75t_L g413 ( .A(n_284), .Y(n_413) );
NAND2xp33_ASAP7_75t_SL g488 ( .A(n_284), .B(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g354 ( .A(n_285), .B(n_333), .Y(n_354) );
AND2x2_ASAP7_75t_L g288 ( .A(n_286), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g391 ( .A(n_286), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B1(n_296), .B2(n_301), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
INVx1_ASAP7_75t_L g370 ( .A(n_289), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_290), .A2(n_329), .B1(n_334), .B2(n_337), .Y(n_328) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g454 ( .A(n_291), .Y(n_454) );
BUFx3_ASAP7_75t_L g419 ( .A(n_292), .Y(n_419) );
INVx1_ASAP7_75t_L g442 ( .A(n_293), .Y(n_442) );
AND2x2_ASAP7_75t_L g380 ( .A(n_294), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g447 ( .A(n_294), .B(n_312), .Y(n_447) );
INVx1_ASAP7_75t_L g481 ( .A(n_294), .Y(n_481) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_296), .A2(n_319), .B(n_321), .Y(n_318) );
OA21x2_ASAP7_75t_L g352 ( .A1(n_296), .A2(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g429 ( .A(n_298), .Y(n_429) );
AND2x2_ASAP7_75t_L g446 ( .A(n_298), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g436 ( .A(n_299), .B(n_395), .Y(n_436) );
AND2x2_ASAP7_75t_L g439 ( .A(n_299), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g448 ( .A(n_299), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g393 ( .A(n_302), .B(n_392), .Y(n_393) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_303), .B(n_332), .Y(n_331) );
NAND2x1_ASAP7_75t_L g407 ( .A(n_303), .B(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_315), .B(n_318), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_313), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_308), .A2(n_324), .B1(n_349), .B2(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_312), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_314), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_314), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g456 ( .A(n_317), .Y(n_456) );
AND2x2_ASAP7_75t_L g443 ( .A(n_320), .B(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_R g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_324), .B(n_407), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_326), .Y(n_501) );
OR3x2_ASAP7_75t_L g824 ( .A(n_326), .B(n_399), .C(n_825), .Y(n_824) );
NAND3x1_ASAP7_75t_SL g326 ( .A(n_327), .B(n_341), .C(n_355), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_338), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_329), .A2(n_439), .B1(n_441), .B2(n_443), .Y(n_438) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_330), .B(n_369), .Y(n_383) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_335), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g404 ( .A(n_335), .B(n_345), .Y(n_404) );
AND2x2_ASAP7_75t_L g428 ( .A(n_335), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_339), .A2(n_435), .B(n_436), .Y(n_434) );
AND2x2_ASAP7_75t_L g486 ( .A(n_339), .B(n_365), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_340), .A2(n_493), .B1(n_496), .B2(n_499), .Y(n_492) );
AOI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_348), .B(n_352), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
BUFx2_ASAP7_75t_L g462 ( .A(n_345), .Y(n_462) );
INVx1_ASAP7_75t_SL g469 ( .A(n_345), .Y(n_469) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_346), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_375), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_358), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_358), .B(n_369), .Y(n_450) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_372), .Y(n_363) );
OR2x6_ASAP7_75t_L g420 ( .A(n_365), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g470 ( .A(n_373), .Y(n_470) );
OR2x2_ASAP7_75t_L g497 ( .A(n_373), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_374), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_385), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_382), .B2(n_384), .Y(n_376) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_379), .Y(n_477) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_393), .B2(n_394), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_473), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_423), .C(n_451), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_411), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_405), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_416), .B1(n_420), .B2(n_422), .Y(n_411) );
NAND2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_413), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_415), .B(n_421), .Y(n_491) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx3_ASAP7_75t_L g479 ( .A(n_419), .Y(n_479) );
INVx2_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_437), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_434), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_433), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_445), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_440), .B(n_481), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B(n_457), .C(n_466), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_454), .A2(n_485), .B(n_487), .C(n_492), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B1(n_463), .B2(n_465), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI21xp5_ASAP7_75t_SL g500 ( .A1(n_473), .A2(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_476), .B(n_484), .Y(n_475) );
AOI21xp33_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_478), .B(n_482), .Y(n_476) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVxp33_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_503), .B(n_809), .Y(n_808) );
AO22x2_ASAP7_75t_L g806 ( .A1(n_504), .A2(n_803), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_713), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_635), .C(n_685), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_602), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_538), .B1(n_555), .B2(n_585), .C(n_594), .Y(n_508) );
INVx1_ASAP7_75t_SL g684 ( .A(n_509), .Y(n_684) );
AND2x4_ASAP7_75t_SL g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g606 ( .A(n_510), .Y(n_606) );
OR2x2_ASAP7_75t_L g628 ( .A(n_510), .B(n_619), .Y(n_628) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_510), .Y(n_643) );
INVx5_ASAP7_75t_L g650 ( .A(n_510), .Y(n_650) );
AND2x4_ASAP7_75t_L g656 ( .A(n_510), .B(n_530), .Y(n_656) );
AND2x2_ASAP7_75t_SL g659 ( .A(n_510), .B(n_587), .Y(n_659) );
OR2x2_ASAP7_75t_L g668 ( .A(n_510), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g675 ( .A(n_510), .B(n_521), .Y(n_675) );
AND2x2_ASAP7_75t_L g776 ( .A(n_510), .B(n_529), .Y(n_776) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx3_ASAP7_75t_SL g627 ( .A(n_520), .Y(n_627) );
AND2x2_ASAP7_75t_L g671 ( .A(n_520), .B(n_587), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_520), .A2(n_675), .B(n_676), .Y(n_674) );
AND2x2_ASAP7_75t_L g712 ( .A(n_520), .B(n_650), .Y(n_712) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_529), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_521), .B(n_530), .Y(n_593) );
OR2x2_ASAP7_75t_L g597 ( .A(n_521), .B(n_530), .Y(n_597) );
INVx1_ASAP7_75t_L g605 ( .A(n_521), .Y(n_605) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
INVx2_ASAP7_75t_L g625 ( .A(n_521), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_521), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g734 ( .A(n_521), .B(n_619), .Y(n_734) );
AND2x2_ASAP7_75t_L g749 ( .A(n_521), .B(n_587), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_530), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_538), .B(n_742), .Y(n_741) );
NOR2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_546), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g571 ( .A(n_540), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_540), .B(n_547), .Y(n_600) );
INVx1_ASAP7_75t_L g610 ( .A(n_540), .Y(n_610) );
INVx2_ASAP7_75t_L g633 ( .A(n_540), .Y(n_633) );
INVx2_ASAP7_75t_L g639 ( .A(n_540), .Y(n_639) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_540), .Y(n_709) );
OR2x2_ASAP7_75t_L g740 ( .A(n_540), .B(n_547), .Y(n_740) );
OR2x2_ASAP7_75t_L g756 ( .A(n_546), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_SL g558 ( .A(n_547), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g583 ( .A(n_547), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g620 ( .A(n_547), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g632 ( .A(n_547), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g645 ( .A(n_547), .B(n_611), .Y(n_645) );
OR2x2_ASAP7_75t_L g653 ( .A(n_547), .B(n_559), .Y(n_653) );
INVx2_ASAP7_75t_L g680 ( .A(n_547), .Y(n_680) );
INVx1_ASAP7_75t_L g698 ( .A(n_547), .Y(n_698) );
NOR2xp33_ASAP7_75t_R g731 ( .A(n_547), .B(n_572), .Y(n_731) );
OR2x6_ASAP7_75t_L g547 ( .A(n_548), .B(n_554), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_581), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_556), .A2(n_623), .B1(n_626), .B2(n_629), .Y(n_622) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_570), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g637 ( .A(n_558), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g672 ( .A(n_558), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g751 ( .A(n_558), .B(n_729), .Y(n_751) );
INVx3_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
AND2x4_ASAP7_75t_L g611 ( .A(n_559), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_559), .B(n_572), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_559), .B(n_633), .Y(n_678) );
AND2x2_ASAP7_75t_L g683 ( .A(n_559), .B(n_680), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_559), .B(n_571), .Y(n_720) );
INVx1_ASAP7_75t_L g790 ( .A(n_559), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_559), .B(n_708), .Y(n_801) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .Y(n_559) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g582 ( .A(n_572), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_572), .B(n_584), .Y(n_601) );
INVx2_ASAP7_75t_L g612 ( .A(n_572), .Y(n_612) );
AND2x2_ASAP7_75t_L g638 ( .A(n_572), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g654 ( .A(n_572), .B(n_633), .Y(n_654) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_572), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_572), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g743 ( .A(n_572), .Y(n_743) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_582), .B(n_610), .Y(n_621) );
AOI221x1_ASAP7_75t_SL g715 ( .A1(n_583), .A2(n_716), .B1(n_719), .B2(n_721), .C(n_725), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_583), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g773 ( .A(n_583), .B(n_638), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_583), .B(n_795), .Y(n_794) );
OR2x2_ASAP7_75t_L g704 ( .A(n_584), .B(n_632), .Y(n_704) );
AND2x2_ASAP7_75t_L g742 ( .A(n_584), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_593), .Y(n_586) );
AND2x2_ASAP7_75t_L g595 ( .A(n_587), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g690 ( .A(n_587), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_587), .B(n_606), .Y(n_695) );
AND2x4_ASAP7_75t_L g724 ( .A(n_587), .B(n_625), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_587), .B(n_656), .Y(n_760) );
OR2x2_ASAP7_75t_L g778 ( .A(n_587), .B(n_709), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_587), .B(n_669), .Y(n_788) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g619 ( .A(n_588), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g644 ( .A(n_593), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_593), .A2(n_652), .B1(n_655), .B2(n_657), .Y(n_651) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVx2_ASAP7_75t_L g607 ( .A(n_595), .Y(n_607) );
AND2x2_ASAP7_75t_L g746 ( .A(n_596), .B(n_606), .Y(n_746) );
AND2x2_ASAP7_75t_L g792 ( .A(n_596), .B(n_659), .Y(n_792) );
AND2x2_ASAP7_75t_L g797 ( .A(n_596), .B(n_648), .Y(n_797) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI32xp33_ASAP7_75t_L g766 ( .A1(n_598), .A2(n_668), .A3(n_748), .B1(n_767), .B2(n_769), .Y(n_766) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
AOI211xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_608), .B(n_613), .C(n_622), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_605), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_606), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g786 ( .A(n_606), .Y(n_786) );
AND2x2_ASAP7_75t_L g696 ( .A(n_608), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_SL g608 ( .A(n_609), .B(n_611), .Y(n_608) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_609), .Y(n_796) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_610), .Y(n_665) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_610), .Y(n_765) );
INVx1_ASAP7_75t_L g662 ( .A(n_611), .Y(n_662) );
AND2x2_ASAP7_75t_L g728 ( .A(n_611), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_611), .B(n_739), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_620), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_615), .A2(n_695), .B(n_696), .Y(n_694) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g624 ( .A(n_619), .B(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_624), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g755 ( .A(n_624), .Y(n_755) );
AND2x2_ASAP7_75t_L g785 ( .A(n_624), .B(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_625), .Y(n_762) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_627), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g702 ( .A(n_628), .Y(n_702) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g661 ( .A(n_632), .B(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_633), .Y(n_729) );
AND2x2_ASAP7_75t_L g738 ( .A(n_634), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_658), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_640), .B1(n_645), .B2(n_646), .C(n_651), .Y(n_636) );
INVx1_ASAP7_75t_L g757 ( .A(n_638), .Y(n_757) );
INVxp33_ASAP7_75t_SL g789 ( .A(n_638), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_640), .A2(n_736), .B(n_744), .Y(n_735) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_644), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g657 ( .A(n_645), .Y(n_657) );
AND2x2_ASAP7_75t_L g692 ( .A(n_645), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g711 ( .A(n_645), .B(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_645), .A2(n_773), .B1(n_774), .B2(n_777), .Y(n_772) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OR2x2_ASAP7_75t_L g667 ( .A(n_648), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_648), .B(n_656), .Y(n_706) );
AND2x4_ASAP7_75t_L g723 ( .A(n_650), .B(n_669), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_650), .B(n_724), .Y(n_770) );
AND2x2_ASAP7_75t_L g782 ( .A(n_650), .B(n_734), .Y(n_782) );
NAND2xp33_ASAP7_75t_L g767 ( .A(n_652), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g710 ( .A(n_653), .Y(n_710) );
INVx1_ASAP7_75t_L g781 ( .A(n_654), .Y(n_781) );
INVx2_ASAP7_75t_SL g733 ( .A(n_656), .Y(n_733) );
AOI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B(n_663), .C(n_681), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_667), .B(n_670), .C(n_674), .Y(n_663) );
OR2x6_ASAP7_75t_SL g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
INVx1_ASAP7_75t_SL g718 ( .A(n_668), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_668), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_673), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_677), .A2(n_760), .B1(n_761), .B2(n_763), .Y(n_759) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_691), .B(n_694), .C(n_699), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_711), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g791 ( .A1(n_710), .A2(n_792), .B1(n_793), .B2(n_797), .C1(n_798), .C2(n_800), .Y(n_791) );
INVx2_ASAP7_75t_L g726 ( .A(n_712), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_752), .C(n_771), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_735), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_723), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_724), .B(n_786), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_730), .B2(n_732), .Y(n_725) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVxp33_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_733), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_741), .A2(n_745), .B1(n_747), .B2(n_750), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
OAI211xp5_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_756), .B(n_758), .C(n_766), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_779), .C(n_791), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B(n_790), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_789), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx9p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_819), .B(n_835), .Y(n_834) );
BUFx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
INVxp67_ASAP7_75t_L g833 ( .A(n_822), .Y(n_833) );
AOI22x1_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_826), .B2(n_827), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g831 ( .A(n_829), .Y(n_831) );
AOI21xp33_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B(n_836), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx2_ASAP7_75t_L g844 ( .A(n_838), .Y(n_844) );
INVx1_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
CKINVDCx11_ASAP7_75t_R g841 ( .A(n_842), .Y(n_841) );
CKINVDCx8_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
endmodule