module real_jpeg_31533_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_536, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_536;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_0),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_1),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_1),
.A2(n_53),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22x1_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_53),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_1),
.A2(n_53),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_2),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_2),
.B(n_522),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_5),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_6),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_6),
.A2(n_173),
.B1(n_283),
.B2(n_359),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_6),
.A2(n_247),
.B1(n_283),
.B2(n_426),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_6),
.A2(n_283),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_7),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_28),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_8),
.A2(n_28),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_8),
.A2(n_28),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_13),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_99),
.B1(n_125),
.B2(n_129),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g236 ( 
.A1(n_13),
.A2(n_99),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_13),
.B(n_210),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_13),
.B(n_106),
.Y(n_452)
);

OAI32xp33_ASAP7_75t_L g470 ( 
.A1(n_13),
.A2(n_417),
.A3(n_471),
.B1(n_476),
.B2(n_482),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_520),
.B(n_532),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_15),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_194),
.B(n_519),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_180),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_18),
.B(n_180),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_153),
.C(n_165),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_20),
.A2(n_153),
.B1(n_154),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_20),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B(n_46),
.Y(n_21)
);

OAI21x1_ASAP7_75t_SL g182 ( 
.A1(n_22),
.A2(n_162),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_27),
.Y(n_159)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_27),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_27),
.Y(n_344)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_35),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_35),
.A2(n_56),
.B(n_156),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2x1p5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_36),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_36),
.B(n_280),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_38),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_38),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_40),
.Y(n_341)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_41),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_42),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_42),
.Y(n_175)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_46),
.B(n_287),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_47),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_56),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_48),
.B(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_52),
.Y(n_161)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_56),
.B(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_56),
.B(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_59),
.Y(n_282)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_61),
.Y(n_348)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_103),
.B2(n_152),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_68),
.A2(n_69),
.B1(n_368),
.B2(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_154),
.C(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_69),
.B(n_190),
.C(n_193),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_69),
.B(n_168),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_69),
.B(n_367),
.C(n_368),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_84),
.B(n_97),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_70),
.B(n_97),
.Y(n_207)
);

NAND2x1p5_ASAP7_75t_L g251 ( 
.A(n_70),
.B(n_209),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_70),
.B(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_70),
.B(n_425),
.Y(n_437)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_71),
.B(n_99),
.Y(n_497)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_78),
.Y(n_234)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_78),
.Y(n_241)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_83),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_84),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_84),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_84),
.B(n_97),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_84),
.B(n_425),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_93),
.B2(n_96),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_89),
.Y(n_216)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_89),
.Y(n_429)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_157),
.B(n_160),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_99),
.B(n_164),
.Y(n_390)
);

AOI32xp33_ASAP7_75t_L g416 ( 
.A1(n_99),
.A2(n_417),
.A3(n_419),
.B1(n_421),
.B2(n_422),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_99),
.B(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_99),
.B(n_230),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_101),
.Y(n_246)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_102),
.Y(n_418)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_132),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_105),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_123),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_106),
.A2(n_132),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_106),
.B(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AO21x2_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_139),
.B(n_147),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_116),
.B2(n_120),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21x1_ASAP7_75t_L g185 ( 
.A1(n_124),
.A2(n_138),
.B(n_186),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_124),
.B(n_138),
.Y(n_276)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_133),
.B(n_369),
.Y(n_368)
);

NAND2x1_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_137),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_142),
.Y(n_420)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_147),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_155),
.B(n_317),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_156),
.B(n_163),
.Y(n_287)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_160),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_162),
.B(n_279),
.Y(n_361)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_166),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_176),
.B(n_177),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_170),
.Y(n_337)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_177),
.B(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_178),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_182),
.B(n_187),
.C(n_189),
.Y(n_529)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g301 ( 
.A(n_184),
.B(n_302),
.C(n_315),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_185),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_295),
.B(n_516),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_255),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_196),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_252),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_197),
.B(n_252),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_217),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_199),
.B(n_202),
.Y(n_294)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_203),
.A2(n_204),
.B(n_206),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_207),
.B(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_208),
.B(n_262),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_208),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_210),
.B(n_483),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_217),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_223),
.B2(n_536),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_219),
.B(n_223),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_220),
.A2(n_221),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_242),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_222),
.A2(n_223),
.B1(n_416),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2x2_ASAP7_75t_SL g321 ( 
.A(n_223),
.B(n_242),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_223),
.B(n_416),
.Y(n_415)
);

AO21x2_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_235),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_228),
.A2(n_306),
.B(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_229),
.B(n_236),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_229),
.B(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_230),
.Y(n_493)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_238),
.Y(n_458)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx4f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_250),
.B(n_251),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_251),
.B(n_303),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_251),
.B(n_424),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_293),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_256),
.B(n_293),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_288),
.C(n_289),
.Y(n_256)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_273),
.C(n_277),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_320),
.Y(n_319)
);

OAI21x1_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2x2_ASAP7_75t_SL g374 ( 
.A(n_264),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

AND2x4_ASAP7_75t_SL g454 ( 
.A(n_265),
.B(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_268),
.A2(n_306),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_268),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_269),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_271),
.Y(n_460)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_271),
.Y(n_475)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_271),
.Y(n_481)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_278),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_276),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_404),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_326),
.B(n_403),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g405 ( 
.A(n_298),
.B(n_397),
.C(n_406),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_322),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_299),
.B(n_322),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_318),
.C(n_321),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_301),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_302),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_303),
.B(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_311),
.B(n_455),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_378),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_321),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_379),
.B(n_397),
.C(n_402),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_370),
.Y(n_327)
);

NAND2x1_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_370),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_362),
.C(n_365),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_355),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_361),
.C(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_336),
.Y(n_386)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx4f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI31xp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.A3(n_342),
.B(n_345),
.Y(n_336)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx11_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_349),
.B(n_354),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_366),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_374),
.C(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_395),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_395),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.C(n_387),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_383),
.B(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_388),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.C(n_391),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_400),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_432),
.B(n_515),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_430),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_430),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.C(n_423),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_412),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_423),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_447),
.B(n_514),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_444),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_434),
.B(n_444),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.C(n_441),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_435),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_462)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_463),
.B(n_513),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_449),
.B(n_461),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.C(n_453),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_450),
.A2(n_451),
.B1(n_452),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_493),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_460),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_464),
.A2(n_489),
.B(n_512),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_468),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_488),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_488),
.Y(n_494)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_495),
.B(n_511),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_494),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_499),
.B(n_510),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_498),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_509),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_526),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_526),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_529),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);


endmodule