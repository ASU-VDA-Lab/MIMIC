module fake_jpeg_3045_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_43),
.B1(n_38),
.B2(n_51),
.Y(n_61)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_0),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_69),
.B1(n_47),
.B2(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_53),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.C(n_47),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_39),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_49),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_39),
.B1(n_52),
.B2(n_51),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_58),
.B1(n_49),
.B2(n_52),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_84),
.B2(n_5),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_38),
.B(n_57),
.C(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_68),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_50),
.B1(n_45),
.B2(n_48),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_83),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_3),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_63),
.C(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_67),
.C(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_110),
.B1(n_118),
.B2(n_24),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_112),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_23),
.B1(n_36),
.B2(n_11),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_7),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_9),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_17),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_37),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_18),
.B(n_19),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_108),
.B(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_20),
.C(n_22),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_133),
.C(n_26),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_27),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_143),
.B(n_145),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_133),
.B1(n_122),
.B2(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_146),
.B1(n_141),
.B2(n_136),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_134),
.C(n_138),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_147),
.A2(n_148),
.B1(n_127),
.B2(n_125),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_125),
.B(n_117),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_111),
.B1(n_140),
.B2(n_32),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_155),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_28),
.Y(n_157)
);


endmodule