module fake_jpeg_315_n_680 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_10),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_22),
.B(n_10),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_68),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_10),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_79),
.B(n_113),
.Y(n_213)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_91),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_92),
.Y(n_217)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_52),
.B(n_0),
.CON(n_95),
.SN(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_95),
.A2(n_24),
.B(n_26),
.C(n_37),
.Y(n_161)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_126),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_102),
.Y(n_222)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_9),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_46),
.Y(n_119)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_9),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_124),
.Y(n_201)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_27),
.B(n_41),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_27),
.B(n_29),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_50),
.C(n_51),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_142),
.B(n_1),
.C(n_5),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_29),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_157),
.B(n_175),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_161),
.B(n_11),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_30),
.B1(n_50),
.B2(n_46),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_162),
.A2(n_172),
.B1(n_186),
.B2(n_187),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_68),
.A2(n_51),
.B1(n_121),
.B2(n_50),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_44),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_119),
.A2(n_51),
.B1(n_41),
.B2(n_44),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_182),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_102),
.B(n_26),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_185),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_62),
.A2(n_30),
.B1(n_42),
.B2(n_37),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_42),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_70),
.A2(n_43),
.B1(n_49),
.B2(n_30),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_60),
.A2(n_46),
.B1(n_43),
.B2(n_32),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_28),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_188),
.B(n_192),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_75),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_191),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_116),
.B(n_28),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_95),
.A2(n_43),
.B1(n_49),
.B2(n_46),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_32),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_196),
.B(n_206),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_69),
.A2(n_35),
.B1(n_49),
.B2(n_48),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_94),
.A2(n_49),
.B1(n_48),
.B2(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_74),
.A2(n_35),
.B1(n_49),
.B2(n_57),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_211),
.B(n_212),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_82),
.B(n_12),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_84),
.A2(n_48),
.B1(n_34),
.B2(n_12),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_97),
.B1(n_89),
.B2(n_88),
.Y(n_230)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_120),
.B1(n_109),
.B2(n_107),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_223),
.A2(n_225),
.B1(n_230),
.B2(n_292),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_168),
.A2(n_92),
.B1(n_100),
.B2(n_99),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_227),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_106),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_228),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_161),
.A2(n_34),
.B(n_14),
.C(n_18),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_229),
.B(n_7),
.Y(n_326)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_147),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_232),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_251),
.Y(n_321)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

INVx11_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_235),
.Y(n_346)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_236),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_172),
.A2(n_193),
.B1(n_186),
.B2(n_200),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_237),
.A2(n_240),
.B1(n_243),
.B2(n_256),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_198),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_238),
.Y(n_324)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_239),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_132),
.A2(n_213),
.B1(n_199),
.B2(n_187),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_241),
.Y(n_362)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_87),
.B1(n_34),
.B2(n_3),
.Y(n_243)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_151),
.A2(n_11),
.B(n_17),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_258),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_134),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_247),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_173),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_253),
.A2(n_171),
.B1(n_220),
.B2(n_159),
.Y(n_339)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_254),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_202),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_183),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_260),
.B1(n_149),
.B2(n_130),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_158),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_259),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_190),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_131),
.Y(n_262)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_263),
.Y(n_360)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_135),
.Y(n_264)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_SL g320 ( 
.A(n_265),
.B(n_209),
.C(n_7),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_197),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_277),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_279),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_195),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_298),
.B1(n_184),
.B2(n_208),
.Y(n_304)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_293),
.C(n_214),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_140),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_276),
.Y(n_311)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_166),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_158),
.B(n_5),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_280),
.Y(n_319)
);

INVx5_ASAP7_75t_SL g279 ( 
.A(n_138),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_168),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

BUFx4f_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_284),
.Y(n_328)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_283),
.Y(n_355)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_138),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_288),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g286 ( 
.A1(n_203),
.A2(n_5),
.B(n_6),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_300),
.Y(n_361)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_143),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_290),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_150),
.B(n_218),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_164),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_291),
.B(n_294),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_174),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_139),
.B(n_6),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_217),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_295),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_143),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_297),
.Y(n_356)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_177),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_145),
.A2(n_7),
.B1(n_146),
.B2(n_173),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_141),
.Y(n_300)
);

CKINVDCx6p67_ASAP7_75t_R g301 ( 
.A(n_141),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_302),
.B1(n_209),
.B2(n_177),
.Y(n_347)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_304),
.B(n_339),
.Y(n_394)
);

OAI21xp33_ASAP7_75t_L g383 ( 
.A1(n_306),
.A2(n_320),
.B(n_326),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_224),
.A2(n_189),
.B1(n_184),
.B2(n_208),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_307),
.B(n_317),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_313),
.A2(n_342),
.B1(n_349),
.B2(n_352),
.Y(n_364)
);

OR2x4_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_154),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_228),
.B(n_169),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_337),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_226),
.A2(n_220),
.B1(n_140),
.B2(n_171),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_334),
.A2(n_340),
.B1(n_339),
.B2(n_331),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_287),
.B(n_170),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_228),
.A2(n_130),
.B1(n_149),
.B2(n_159),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_179),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_350),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_237),
.A2(n_163),
.B1(n_165),
.B2(n_177),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_163),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_250),
.A2(n_299),
.B1(n_275),
.B2(n_265),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_250),
.A2(n_165),
.B1(n_265),
.B2(n_274),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_354),
.A2(n_357),
.B1(n_292),
.B2(n_288),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_257),
.A2(n_260),
.B1(n_244),
.B2(n_268),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_278),
.B(n_239),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_301),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_317),
.A2(n_243),
.B1(n_256),
.B2(n_279),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_365),
.A2(n_398),
.B(n_399),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_366),
.A2(n_370),
.B1(n_402),
.B2(n_403),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_314),
.A2(n_342),
.B(n_361),
.C(n_318),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_367),
.A2(n_375),
.B(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_321),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_369),
.B(n_380),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_331),
.A2(n_269),
.B1(n_273),
.B2(n_263),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_371),
.B(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_271),
.C(n_234),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_314),
.A2(n_301),
.B(n_285),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_328),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_242),
.C(n_291),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_377),
.B(n_384),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_255),
.B1(n_249),
.B2(n_248),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_379),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_310),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_302),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_314),
.A2(n_301),
.B(n_292),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_281),
.B1(n_294),
.B2(n_238),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_238),
.B1(n_276),
.B2(n_272),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_352),
.A2(n_227),
.B1(n_261),
.B2(n_295),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_390),
.B(n_393),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_392),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_319),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_282),
.C(n_259),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_324),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_400),
.Y(n_427)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_245),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_283),
.C(n_235),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_322),
.B(n_233),
.C(n_241),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_322),
.B(n_231),
.C(n_232),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_404),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_349),
.A2(n_297),
.B1(n_254),
.B2(n_236),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_358),
.A2(n_326),
.B1(n_305),
.B2(n_356),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_252),
.C(n_267),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_311),
.A2(n_363),
.B1(n_344),
.B2(n_343),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_359),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_330),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_409),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_375),
.A2(n_385),
.B(n_367),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_413),
.A2(n_436),
.B(n_437),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_364),
.A2(n_311),
.B1(n_363),
.B2(n_360),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_422),
.A2(n_449),
.B1(n_388),
.B2(n_370),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_365),
.A2(n_351),
.B(n_329),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_435),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_409),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_367),
.A2(n_405),
.B(n_390),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_367),
.A2(n_355),
.B(n_351),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_329),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_444),
.Y(n_466)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_406),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_382),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_343),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_316),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_381),
.B(n_316),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_445),
.B(n_327),
.Y(n_472)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_447),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_366),
.A2(n_348),
.B1(n_359),
.B2(n_323),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_364),
.A2(n_360),
.B1(n_335),
.B2(n_332),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_450),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_384),
.C(n_446),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_454),
.C(n_468),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_451),
.A2(n_405),
.B1(n_371),
.B2(n_394),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_453),
.A2(n_424),
.B1(n_438),
.B2(n_450),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_374),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g522 ( 
.A(n_455),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_436),
.B(n_382),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_462),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_461),
.A2(n_473),
.B1(n_475),
.B2(n_420),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_436),
.B(n_377),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_412),
.B(n_383),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_463),
.B(n_467),
.Y(n_513)
);

AO22x1_ASAP7_75t_L g464 ( 
.A1(n_442),
.A2(n_398),
.B1(n_367),
.B2(n_394),
.Y(n_464)
);

AOI22x1_ASAP7_75t_L g515 ( 
.A1(n_464),
.A2(n_423),
.B1(n_449),
.B2(n_372),
.Y(n_515)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_465),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_412),
.B(n_400),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_393),
.C(n_404),
.Y(n_468)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_394),
.B1(n_398),
.B2(n_389),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_398),
.B1(n_402),
.B2(n_387),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_309),
.Y(n_476)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_416),
.B(n_401),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_477),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_416),
.B(n_323),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_478),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_399),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_437),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_309),
.C(n_348),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_483),
.C(n_484),
.Y(n_505)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_482),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_432),
.B(n_303),
.C(n_315),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_427),
.B(n_303),
.C(n_315),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

OAI32xp33_ASAP7_75t_L g488 ( 
.A1(n_444),
.A2(n_372),
.A3(n_378),
.B1(n_325),
.B2(n_410),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_488),
.B(n_426),
.Y(n_491)
);

OAI31xp33_ASAP7_75t_L g539 ( 
.A1(n_491),
.A2(n_512),
.A3(n_515),
.B(n_470),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_453),
.A2(n_469),
.B1(n_473),
.B2(n_460),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_492),
.A2(n_493),
.B1(n_501),
.B2(n_511),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_413),
.B1(n_414),
.B2(n_437),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_486),
.A2(n_414),
.B(n_413),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_496),
.A2(n_499),
.B(n_456),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_502),
.B1(n_479),
.B2(n_475),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_498),
.B(n_500),
.C(n_507),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_486),
.A2(n_421),
.B1(n_440),
.B2(n_419),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_427),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_460),
.A2(n_414),
.B1(n_422),
.B2(n_421),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_457),
.A2(n_448),
.B1(n_445),
.B2(n_419),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_454),
.B(n_433),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_457),
.B(n_433),
.Y(n_508)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_466),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_519),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_422),
.B1(n_449),
.B2(n_420),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_423),
.B(n_419),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_461),
.A2(n_417),
.B1(n_435),
.B2(n_447),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_514),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_468),
.B(n_417),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_362),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_471),
.B(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_462),
.B(n_418),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_464),
.A2(n_441),
.B1(n_424),
.B2(n_439),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_520),
.A2(n_525),
.B1(n_482),
.B2(n_431),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_487),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_480),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_526),
.B(n_537),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_504),
.Y(n_528)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_459),
.Y(n_531)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_471),
.Y(n_532)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_532),
.Y(n_567)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_517),
.Y(n_533)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_533),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_535),
.A2(n_539),
.B(n_556),
.Y(n_580)
);

CKINVDCx14_ASAP7_75t_R g565 ( 
.A(n_536),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_491),
.A2(n_488),
.B(n_481),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_483),
.B1(n_470),
.B2(n_458),
.Y(n_538)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_538),
.Y(n_576)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_540),
.Y(n_571)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_503),
.Y(n_543)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_543),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_490),
.B(n_484),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_544),
.Y(n_572)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_520),
.Y(n_545)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_545),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_511),
.A2(n_485),
.B1(n_418),
.B2(n_430),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_547),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_513),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_492),
.A2(n_430),
.B1(n_474),
.B2(n_465),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_548),
.B(n_549),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_522),
.B(n_525),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_550),
.B(n_498),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_524),
.B(n_434),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_552),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_505),
.B(n_434),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_493),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_505),
.C(n_501),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_555),
.Y(n_579)
);

AOI322xp5_ASAP7_75t_L g555 ( 
.A1(n_512),
.A2(n_431),
.A3(n_407),
.B1(n_379),
.B2(n_332),
.C1(n_338),
.C2(n_327),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_518),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_325),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_557),
.B(n_495),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_561),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_507),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_500),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_568),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_544),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_494),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_535),
.B(n_489),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_581),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_494),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_496),
.B(n_515),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_582),
.A2(n_515),
.B(n_541),
.Y(n_602)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_516),
.C(n_519),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_585),
.B(n_551),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_538),
.C(n_526),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_586),
.B(n_591),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_546),
.Y(n_588)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_566),
.Y(n_589)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_589),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_598),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_532),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_563),
.C(n_585),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_594),
.Y(n_620)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_567),
.Y(n_593)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_593),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_562),
.A2(n_534),
.B1(n_549),
.B2(n_545),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_531),
.B1(n_537),
.B2(n_565),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_607),
.B1(n_580),
.B2(n_560),
.Y(n_614)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_596),
.B(n_600),
.Y(n_625)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_583),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_562),
.A2(n_541),
.B1(n_537),
.B2(n_540),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_601),
.A2(n_582),
.B1(n_580),
.B2(n_576),
.Y(n_610)
);

OAI321xp33_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_604),
.A3(n_537),
.B1(n_569),
.B2(n_529),
.C(n_575),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_568),
.B(n_530),
.C(n_489),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_573),
.C(n_576),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_575),
.B(n_556),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_562),
.A2(n_527),
.B1(n_529),
.B2(n_533),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_606),
.B(n_608),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_584),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_579),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_561),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_621),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_610),
.A2(n_614),
.B1(n_619),
.B2(n_628),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_601),
.A2(n_527),
.B1(n_571),
.B2(n_570),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_611),
.B(n_627),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_612),
.B(n_599),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_569),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_618),
.B(n_623),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_587),
.B(n_559),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_586),
.B(n_577),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_592),
.B(n_548),
.C(n_554),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_626),
.B(n_588),
.C(n_605),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_594),
.B(n_499),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_602),
.A2(n_578),
.B1(n_574),
.B2(n_543),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_620),
.A2(n_588),
.B1(n_604),
.B2(n_597),
.Y(n_629)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_628),
.Y(n_630)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_630),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_603),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_634),
.B(n_638),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_625),
.A2(n_600),
.B(n_597),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_635),
.A2(n_618),
.B(n_617),
.Y(n_647)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_616),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_636),
.A2(n_642),
.B1(n_643),
.B2(n_615),
.Y(n_645)
);

MAJx2_ASAP7_75t_L g637 ( 
.A(n_612),
.B(n_605),
.C(n_606),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_SL g651 ( 
.A(n_637),
.B(n_617),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_613),
.A2(n_542),
.B(n_528),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_639),
.A2(n_640),
.B(n_641),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_616),
.B(n_599),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_622),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_624),
.Y(n_643)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_645),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_647),
.B(n_648),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_638),
.B(n_626),
.C(n_609),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_637),
.C(n_644),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_650),
.B(n_632),
.C(n_630),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_651),
.B(n_655),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_633),
.A2(n_627),
.B(n_621),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_654),
.A2(n_635),
.B(n_631),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_644),
.B(n_557),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_633),
.B(n_495),
.C(n_506),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_656),
.B(n_632),
.C(n_506),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_650),
.B(n_639),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_659),
.Y(n_669)
);

MAJx2_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_661),
.C(n_651),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_653),
.B(n_630),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_662),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_653),
.B(n_630),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_664),
.B(n_646),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_666),
.B(n_667),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_665),
.A2(n_652),
.B(n_649),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_670),
.B(n_661),
.C(n_649),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_672),
.B(n_673),
.C(n_668),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_669),
.B(n_660),
.C(n_648),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_674),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_SL g675 ( 
.A1(n_671),
.A2(n_663),
.B(n_655),
.C(n_355),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_663),
.C(n_675),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_677),
.A2(n_338),
.B(n_346),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_346),
.C(n_362),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_679),
.B(n_327),
.Y(n_680)
);


endmodule