module real_aes_1203_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g529 ( .A(n_0), .B(n_226), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_1), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_2), .Y(n_831) );
INVx1_ASAP7_75t_L g160 ( .A(n_3), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_4), .B(n_532), .Y(n_551) );
NAND2xp33_ASAP7_75t_SL g522 ( .A(n_5), .B(n_181), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_6), .B(n_194), .Y(n_217) );
INVx1_ASAP7_75t_L g514 ( .A(n_7), .Y(n_514) );
INVx1_ASAP7_75t_L g251 ( .A(n_8), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_9), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_10), .Y(n_268) );
AND2x2_ASAP7_75t_L g549 ( .A(n_11), .B(n_150), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_12), .A2(n_796), .B1(n_803), .B2(n_805), .Y(n_802) );
INVx2_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
AND3x1_ASAP7_75t_L g113 ( .A(n_14), .B(n_35), .C(n_114), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_14), .Y(n_129) );
INVx1_ASAP7_75t_L g227 ( .A(n_15), .Y(n_227) );
AOI221x1_ASAP7_75t_L g517 ( .A1(n_16), .A2(n_183), .B1(n_518), .B2(n_520), .C(n_521), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_17), .B(n_532), .Y(n_585) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_18), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g133 ( .A(n_18), .Y(n_133) );
INVx1_ASAP7_75t_L g224 ( .A(n_19), .Y(n_224) );
INVx1_ASAP7_75t_SL g172 ( .A(n_20), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_21), .B(n_175), .Y(n_197) );
AOI33xp33_ASAP7_75t_L g242 ( .A1(n_22), .A2(n_49), .A3(n_157), .B1(n_168), .B2(n_243), .B3(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_23), .A2(n_520), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_24), .B(n_226), .Y(n_554) );
AOI221xp5_ASAP7_75t_SL g594 ( .A1(n_25), .A2(n_40), .B1(n_520), .B2(n_532), .C(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g261 ( .A(n_26), .Y(n_261) );
OR2x2_ASAP7_75t_L g152 ( .A(n_27), .B(n_91), .Y(n_152) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_27), .A2(n_91), .B(n_151), .Y(n_185) );
INVxp67_ASAP7_75t_L g516 ( .A(n_28), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_29), .B(n_229), .Y(n_589) );
AND2x2_ASAP7_75t_L g543 ( .A(n_30), .B(n_149), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_31), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_32), .A2(n_520), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_33), .B(n_229), .Y(n_596) );
AND2x2_ASAP7_75t_L g162 ( .A(n_34), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g167 ( .A(n_34), .Y(n_167) );
AND2x2_ASAP7_75t_L g181 ( .A(n_34), .B(n_160), .Y(n_181) );
OR2x6_ASAP7_75t_L g131 ( .A(n_35), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_36), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_37), .B(n_155), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_38), .A2(n_184), .B1(n_190), .B2(n_194), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_39), .B(n_199), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_41), .A2(n_83), .B1(n_165), .B2(n_520), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_42), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_43), .B(n_226), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_44), .B(n_201), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_45), .B(n_175), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
AND2x2_ASAP7_75t_L g533 ( .A(n_47), .B(n_149), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_48), .B(n_149), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_50), .B(n_175), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_51), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_51), .A2(n_63), .B1(n_440), .B2(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g158 ( .A(n_52), .Y(n_158) );
INVx1_ASAP7_75t_L g177 ( .A(n_52), .Y(n_177) );
AOI22x1_ASAP7_75t_L g796 ( .A1(n_53), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_53), .Y(n_797) );
AND2x2_ASAP7_75t_L g293 ( .A(n_54), .B(n_149), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_55), .A2(n_76), .B1(n_155), .B2(n_165), .C(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_56), .B(n_155), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_57), .B(n_532), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_58), .A2(n_808), .B(n_823), .Y(n_807) );
INVx1_ASAP7_75t_L g826 ( .A(n_58), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_59), .B(n_184), .Y(n_270) );
AOI21xp5_ASAP7_75t_SL g206 ( .A1(n_60), .A2(n_165), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g570 ( .A(n_61), .B(n_149), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_229), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_63), .Y(n_821) );
INVx1_ASAP7_75t_L g220 ( .A(n_64), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_65), .B(n_226), .Y(n_568) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_66), .B(n_150), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_67), .A2(n_520), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g291 ( .A(n_68), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_69), .B(n_229), .Y(n_555) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_70), .B(n_201), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_71), .A2(n_103), .B1(n_800), .B2(n_801), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_71), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_72), .A2(n_165), .B(n_290), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_73), .A2(n_819), .B1(n_820), .B2(n_822), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_73), .Y(n_819) );
INVx1_ASAP7_75t_L g163 ( .A(n_74), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_74), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_75), .B(n_155), .Y(n_245) );
AND2x2_ASAP7_75t_L g182 ( .A(n_77), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g221 ( .A(n_78), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_79), .A2(n_165), .B(n_171), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_80), .A2(n_165), .B(n_196), .C(n_200), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_81), .A2(n_86), .B1(n_155), .B2(n_532), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_82), .B(n_532), .Y(n_569) );
INVx1_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_85), .B(n_183), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_87), .A2(n_165), .B1(n_240), .B2(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_88), .B(n_226), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_89), .B(n_226), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_90), .A2(n_520), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g208 ( .A(n_92), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_93), .B(n_229), .Y(n_567) );
AND2x2_ASAP7_75t_L g246 ( .A(n_94), .B(n_183), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_95), .A2(n_259), .B(n_260), .C(n_262), .Y(n_258) );
INVxp67_ASAP7_75t_L g519 ( .A(n_96), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_97), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_98), .B(n_229), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_99), .A2(n_520), .B(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_100), .Y(n_126) );
BUFx2_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_102), .B(n_175), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_103), .Y(n_801) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_830), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_107), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_111), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_134), .B1(n_807), .B2(n_828), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
CKINVDCx11_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g829 ( .A(n_120), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_125), .A2(n_824), .B(n_825), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g827 ( .A(n_127), .Y(n_827) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g811 ( .A(n_128), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x6_ASAP7_75t_SL g504 ( .A(n_129), .B(n_131), .Y(n_504) );
OR2x6_ASAP7_75t_SL g795 ( .A(n_129), .B(n_130), .Y(n_795) );
OR2x2_ASAP7_75t_L g806 ( .A(n_129), .B(n_131), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_796), .B(n_802), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_503), .B1(n_505), .B2(n_793), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_138), .A2(n_503), .B1(n_506), .B2(n_804), .Y(n_803) );
AND3x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_497), .C(n_500), .Y(n_138) );
NAND5xp2_ASAP7_75t_L g139 ( .A(n_140), .B(n_397), .C(n_427), .D(n_441), .E(n_467), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_141), .A2(n_440), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g815 ( .A(n_141), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_346), .Y(n_141) );
NOR3xp33_ASAP7_75t_SL g142 ( .A(n_143), .B(n_294), .C(n_328), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_211), .B(n_233), .C(n_272), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_186), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_146), .B(n_284), .Y(n_349) );
AND2x2_ASAP7_75t_L g436 ( .A(n_146), .B(n_214), .Y(n_436) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g232 ( .A(n_147), .B(n_203), .Y(n_232) );
INVx1_ASAP7_75t_L g274 ( .A(n_147), .Y(n_274) );
INVx2_ASAP7_75t_L g279 ( .A(n_147), .Y(n_279) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_147), .Y(n_307) );
INVx1_ASAP7_75t_L g321 ( .A(n_147), .Y(n_321) );
AND2x2_ASAP7_75t_L g325 ( .A(n_147), .B(n_216), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_147), .B(n_215), .Y(n_406) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_153), .B(n_182), .Y(n_147) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_148), .A2(n_537), .B(n_543), .Y(n_536) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_148), .A2(n_564), .B(n_570), .Y(n_563) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_148), .A2(n_537), .B(n_543), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_149), .Y(n_148) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_149), .A2(n_594), .B(n_598), .Y(n_593) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x4_ASAP7_75t_L g194 ( .A(n_151), .B(n_152), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_164), .Y(n_153) );
INVx1_ASAP7_75t_L g271 ( .A(n_155), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_155), .A2(n_165), .B1(n_513), .B2(n_515), .Y(n_512) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_161), .Y(n_155) );
INVx1_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
OR2x6_ASAP7_75t_L g173 ( .A(n_157), .B(n_169), .Y(n_173) );
INVxp33_ASAP7_75t_L g243 ( .A(n_157), .Y(n_243) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g170 ( .A(n_158), .B(n_160), .Y(n_170) );
AND2x4_ASAP7_75t_L g229 ( .A(n_158), .B(n_178), .Y(n_229) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x6_ASAP7_75t_L g520 ( .A(n_162), .B(n_170), .Y(n_520) );
INVx2_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
AND2x6_ASAP7_75t_L g226 ( .A(n_163), .B(n_176), .Y(n_226) );
INVxp67_ASAP7_75t_L g269 ( .A(n_165), .Y(n_269) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
NOR2x1p5_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g244 ( .A(n_168), .Y(n_244) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_180), .Y(n_171) );
INVx2_ASAP7_75t_L g199 ( .A(n_173), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_173), .A2(n_180), .B(n_208), .C(n_209), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_173), .A2(n_220), .B1(n_221), .B2(n_222), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_173), .A2(n_180), .B(n_251), .C(n_252), .Y(n_250) );
INVxp67_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_173), .A2(n_180), .B(n_291), .C(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
AND2x4_ASAP7_75t_L g532 ( .A(n_175), .B(n_181), .Y(n_532) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_197), .B(n_198), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_180), .B(n_194), .Y(n_230) );
INVx1_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_180), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_180), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_180), .A2(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_180), .A2(n_567), .B(n_568), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_180), .A2(n_588), .B(n_589), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_180), .A2(n_596), .B(n_597), .Y(n_595) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_183), .A2(n_258), .B1(n_263), .B2(n_264), .Y(n_257) );
INVx3_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_184), .B(n_267), .Y(n_266) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_184), .A2(n_526), .B(n_533), .Y(n_525) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_185), .Y(n_201) );
AND2x4_ASAP7_75t_SL g186 ( .A(n_187), .B(n_202), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g231 ( .A(n_188), .Y(n_231) );
AND2x2_ASAP7_75t_L g275 ( .A(n_188), .B(n_216), .Y(n_275) );
AND2x2_ASAP7_75t_L g296 ( .A(n_188), .B(n_203), .Y(n_296) );
INVx1_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
AND2x4_ASAP7_75t_L g386 ( .A(n_188), .B(n_215), .Y(n_386) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_195), .Y(n_188) );
NOR3xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .C(n_193), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_194), .A2(n_206), .B(n_210), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_194), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_194), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_194), .B(n_519), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_194), .B(n_222), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_194), .A2(n_551), .B(n_552), .Y(n_550) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_200), .A2(n_238), .B(n_246), .Y(n_237) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_200), .A2(n_238), .B(n_246), .Y(n_301) );
AOI21x1_ASAP7_75t_L g558 ( .A1(n_200), .A2(n_559), .B(n_562), .Y(n_558) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_201), .A2(n_249), .B(n_253), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_201), .A2(n_585), .B(n_586), .Y(n_584) );
AND2x4_ASAP7_75t_L g402 ( .A(n_202), .B(n_319), .Y(n_402) );
OR2x2_ASAP7_75t_L g443 ( .A(n_202), .B(n_444), .Y(n_443) );
NOR2xp67_ASAP7_75t_SL g462 ( .A(n_202), .B(n_335), .Y(n_462) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_202), .B(n_394), .Y(n_480) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2x1_ASAP7_75t_SL g280 ( .A(n_203), .B(n_216), .Y(n_280) );
AND2x4_ASAP7_75t_L g318 ( .A(n_203), .B(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_203), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_203), .B(n_278), .Y(n_356) );
INVx2_ASAP7_75t_L g370 ( .A(n_203), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_203), .B(n_322), .Y(n_392) );
AND2x2_ASAP7_75t_L g484 ( .A(n_203), .B(n_342), .Y(n_484) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2x1_ASAP7_75t_L g212 ( .A(n_213), .B(n_232), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_214), .B(n_321), .Y(n_335) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_214), .B(n_324), .Y(n_344) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_231), .Y(n_214) );
INVx1_ASAP7_75t_L g322 ( .A(n_215), .Y(n_322) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g342 ( .A(n_216), .Y(n_342) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_223), .B(n_230), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_222), .B(n_261), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B1(n_227), .B2(n_228), .Y(n_223) );
INVxp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g375 ( .A(n_231), .Y(n_375) );
INVx2_ASAP7_75t_SL g420 ( .A(n_232), .Y(n_420) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_254), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_235), .B(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g366 ( .A(n_235), .Y(n_366) );
AND2x2_ASAP7_75t_L g490 ( .A(n_235), .B(n_315), .Y(n_490) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_247), .Y(n_235) );
AND2x4_ASAP7_75t_L g303 ( .A(n_236), .B(n_285), .Y(n_303) );
INVx1_ASAP7_75t_L g314 ( .A(n_236), .Y(n_314) );
AND2x2_ASAP7_75t_L g345 ( .A(n_236), .B(n_300), .Y(n_345) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_237), .B(n_248), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_237), .B(n_286), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_239), .B(n_245), .Y(n_238) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
AND2x4_ASAP7_75t_L g351 ( .A(n_248), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g363 ( .A(n_248), .Y(n_363) );
INVx1_ASAP7_75t_L g405 ( .A(n_248), .Y(n_405) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_248), .Y(n_417) );
AND2x2_ASAP7_75t_L g433 ( .A(n_248), .B(n_256), .Y(n_433) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g380 ( .A(n_255), .B(n_338), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_255), .Y(n_382) );
AND2x2_ASAP7_75t_L g403 ( .A(n_255), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g282 ( .A(n_256), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g310 ( .A(n_256), .Y(n_310) );
INVx2_ASAP7_75t_L g316 ( .A(n_256), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_256), .B(n_286), .Y(n_331) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_265), .Y(n_256) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_287), .B(n_293), .Y(n_286) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_264), .A2(n_287), .B(n_293), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B1(n_270), .B2(n_271), .Y(n_265) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_281), .Y(n_272) );
INVx1_ASAP7_75t_L g412 ( .A(n_273), .Y(n_412) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g332 ( .A(n_275), .Y(n_332) );
AND2x2_ASAP7_75t_L g388 ( .A(n_275), .B(n_324), .Y(n_388) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_277), .B(n_318), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_277), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g409 ( .A(n_277), .B(n_402), .Y(n_409) );
AND2x2_ASAP7_75t_L g483 ( .A(n_277), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_278), .Y(n_471) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_279), .Y(n_391) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_305), .Y(n_304) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_280), .A2(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx3_ASAP7_75t_L g378 ( .A(n_282), .Y(n_378) );
NAND2x1_ASAP7_75t_SL g422 ( .A(n_282), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g425 ( .A(n_282), .B(n_303), .Y(n_425) );
AND2x2_ASAP7_75t_L g337 ( .A(n_284), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g474 ( .A(n_284), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g485 ( .A(n_284), .B(n_433), .Y(n_485) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_285), .B(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g416 ( .A(n_286), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_308), .B(n_311), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B1(n_303), .B2(n_304), .Y(n_295) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g432 ( .A(n_298), .B(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_298), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_298), .B(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g315 ( .A(n_300), .B(n_316), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_300), .B(n_316), .Y(n_396) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_300), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
AND2x2_ASAP7_75t_L g360 ( .A(n_301), .B(n_316), .Y(n_360) );
INVx1_ASAP7_75t_L g423 ( .A(n_301), .Y(n_423) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2x1_ASAP7_75t_L g341 ( .A(n_306), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g453 ( .A(n_309), .B(n_338), .Y(n_453) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_310), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g438 ( .A(n_310), .B(n_345), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_317), .B1(n_323), .B2(n_326), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g446 ( .A(n_313), .B(n_447), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g476 ( .A(n_316), .B(n_363), .Y(n_476) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx2_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
OAI21xp33_ASAP7_75t_SL g489 ( .A1(n_318), .A2(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_321), .Y(n_479) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_SL g421 ( .A1(n_324), .A2(n_422), .B(n_424), .C(n_426), .Y(n_421) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_325), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g426 ( .A(n_325), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_325), .B(n_402), .Y(n_466) );
INVx1_ASAP7_75t_SL g333 ( .A(n_326), .Y(n_333) );
AND2x2_ASAP7_75t_L g414 ( .A(n_327), .B(n_351), .Y(n_414) );
INVx1_ASAP7_75t_L g459 ( .A(n_327), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_333), .B2(n_334), .C(n_336), .Y(n_328) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_329), .Y(n_448) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g496 ( .A(n_331), .B(n_339), .Y(n_496) );
OR2x2_ASAP7_75t_L g355 ( .A(n_332), .B(n_356), .Y(n_355) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_332), .B(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_332), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g494 ( .A(n_332), .B(n_391), .Y(n_494) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI32xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .A3(n_343), .B1(n_344), .B2(n_345), .Y(n_336) );
INVx1_ASAP7_75t_L g357 ( .A(n_338), .Y(n_357) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_340), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g452 ( .A(n_341), .Y(n_452) );
OAI22xp33_ASAP7_75t_SL g434 ( .A1(n_343), .A2(n_435), .B1(n_437), .B2(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g465 ( .A(n_344), .Y(n_465) );
AOI211x1_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_353), .B(n_354), .C(n_371), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_348), .B(n_433), .Y(n_439) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g395 ( .A(n_351), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g461 ( .A(n_351), .Y(n_461) );
OAI222xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B1(n_358), .B2(n_364), .C1(n_365), .C2(n_367), .Y(n_354) );
INVxp67_ASAP7_75t_L g451 ( .A(n_355), .Y(n_451) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_359), .B(n_444), .Y(n_491) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g407 ( .A(n_360), .B(n_404), .Y(n_407) );
INVx3_ASAP7_75t_L g447 ( .A(n_362), .Y(n_447) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g385 ( .A(n_370), .B(n_386), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B1(n_379), .B2(n_384), .C(n_387), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_373), .A2(n_430), .B(n_432), .Y(n_429) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g383 ( .A(n_377), .Y(n_383) );
OR2x2_ASAP7_75t_L g487 ( .A(n_378), .B(n_423), .Y(n_487) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_381), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_384), .A2(n_413), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_385), .A2(n_457), .B(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g394 ( .A(n_386), .Y(n_394) );
OAI31xp33_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .A3(n_393), .B(n_395), .Y(n_387) );
INVx1_ASAP7_75t_L g445 ( .A(n_389), .Y(n_445) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_410), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_398), .B(n_410), .C(n_429), .D(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_408), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B1(n_406), .B2(n_407), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_403), .B(n_423), .Y(n_431) );
INVx1_ASAP7_75t_SL g444 ( .A(n_406), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_421), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_415), .B2(n_418), .Y(n_411) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_420), .A2(n_483), .B1(n_485), .B2(n_486), .Y(n_482) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_434), .C(n_440), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_440), .A2(n_501), .B(n_502), .Y(n_500) );
INVxp33_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
AND2x2_ASAP7_75t_L g814 ( .A(n_441), .B(n_467), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_446), .A2(n_469), .B(n_472), .Y(n_468) );
INVx2_ASAP7_75t_L g456 ( .A(n_447), .Y(n_456) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_454), .C(n_463), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_457), .B1(n_460), .B2(n_462), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVxp33_ASAP7_75t_SL g502 ( .A(n_467), .Y(n_502) );
NOR3x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_481), .C(n_488), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_477), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_489), .B(n_492), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g816 ( .A(n_498), .Y(n_816) );
CKINVDCx11_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_670), .Y(n_506) );
NOR4xp25_ASAP7_75t_L g507 ( .A(n_508), .B(n_613), .C(n_652), .D(n_659), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_534), .B1(n_571), .B2(n_580), .C(n_599), .Y(n_508) );
OR2x2_ASAP7_75t_L g743 ( .A(n_509), .B(n_605), .Y(n_743) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g658 ( .A(n_510), .B(n_583), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_510), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_510), .B(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_523), .Y(n_510) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_511), .B(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g604 ( .A(n_511), .Y(n_604) );
AND2x2_ASAP7_75t_L g639 ( .A(n_511), .B(n_612), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_511), .B(n_524), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_511), .B(n_606), .Y(n_691) );
OR2x2_ASAP7_75t_L g769 ( .A(n_511), .B(n_583), .Y(n_769) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .Y(n_511) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g591 ( .A(n_524), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_524), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g617 ( .A(n_524), .Y(n_617) );
OR2x2_ASAP7_75t_L g622 ( .A(n_524), .B(n_606), .Y(n_622) );
AND2x2_ASAP7_75t_L g635 ( .A(n_524), .B(n_593), .Y(n_635) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_524), .Y(n_638) );
INVx1_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_524), .B(n_604), .Y(n_715) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_544), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g579 ( .A(n_536), .B(n_563), .Y(n_579) );
AND2x4_ASAP7_75t_L g609 ( .A(n_536), .B(n_548), .Y(n_609) );
INVx2_ASAP7_75t_L g643 ( .A(n_536), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_536), .B(n_563), .Y(n_701) );
AND2x2_ASAP7_75t_L g748 ( .A(n_536), .B(n_577), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g736 ( .A1(n_544), .A2(n_608), .B1(n_651), .B2(n_711), .C1(n_737), .C2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
AND2x2_ASAP7_75t_L g655 ( .A(n_546), .B(n_575), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_546), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g784 ( .A(n_546), .B(n_624), .Y(n_784) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_547), .A2(n_615), .B(n_619), .Y(n_614) );
AND2x2_ASAP7_75t_L g695 ( .A(n_547), .B(n_578), .Y(n_695) );
OR2x2_ASAP7_75t_L g720 ( .A(n_547), .B(n_579), .Y(n_720) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx5_ASAP7_75t_L g574 ( .A(n_548), .Y(n_574) );
AND2x2_ASAP7_75t_L g661 ( .A(n_548), .B(n_643), .Y(n_661) );
AND2x2_ASAP7_75t_L g687 ( .A(n_548), .B(n_563), .Y(n_687) );
OR2x2_ASAP7_75t_L g690 ( .A(n_548), .B(n_577), .Y(n_690) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_548), .Y(n_708) );
AND2x4_ASAP7_75t_SL g765 ( .A(n_548), .B(n_642), .Y(n_765) );
OR2x2_ASAP7_75t_L g774 ( .A(n_548), .B(n_601), .Y(n_774) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g607 ( .A(n_556), .Y(n_607) );
AOI221xp5_ASAP7_75t_SL g725 ( .A1(n_556), .A2(n_609), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_725) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_563), .Y(n_556) );
OR2x2_ASAP7_75t_L g664 ( .A(n_557), .B(n_634), .Y(n_664) );
OR2x2_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g700 ( .A(n_557), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g706 ( .A(n_557), .B(n_625), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_557), .B(n_689), .Y(n_718) );
INVx2_ASAP7_75t_L g731 ( .A(n_557), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_557), .B(n_609), .Y(n_752) );
AND2x2_ASAP7_75t_L g756 ( .A(n_557), .B(n_578), .Y(n_756) );
AND2x2_ASAP7_75t_L g764 ( .A(n_557), .B(n_765), .Y(n_764) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_558), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_563), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_577), .Y(n_608) );
INVx2_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
AND2x4_ASAP7_75t_L g642 ( .A(n_563), .B(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_563), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g754 ( .A(n_573), .B(n_576), .Y(n_754) );
AND2x4_ASAP7_75t_L g600 ( .A(n_574), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g641 ( .A(n_574), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g668 ( .A(n_574), .B(n_608), .Y(n_668) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g772 ( .A(n_576), .B(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g624 ( .A(n_577), .B(n_625), .Y(n_624) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_578), .A2(n_645), .B(n_651), .Y(n_644) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_591), .Y(n_581) );
INVx1_ASAP7_75t_SL g698 ( .A(n_582), .Y(n_698) );
AND2x2_ASAP7_75t_L g728 ( .A(n_582), .B(n_638), .Y(n_728) );
AND2x4_ASAP7_75t_L g739 ( .A(n_582), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g605 ( .A(n_583), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g612 ( .A(n_583), .Y(n_612) );
AND2x4_ASAP7_75t_L g618 ( .A(n_583), .B(n_604), .Y(n_618) );
INVx2_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
INVx1_ASAP7_75t_L g678 ( .A(n_583), .Y(n_678) );
OR2x2_ASAP7_75t_L g699 ( .A(n_583), .B(n_683), .Y(n_699) );
OR2x2_ASAP7_75t_L g713 ( .A(n_583), .B(n_593), .Y(n_713) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_583), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_583), .B(n_635), .Y(n_785) );
OR2x6_ASAP7_75t_L g583 ( .A(n_584), .B(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g630 ( .A(n_591), .Y(n_630) );
AND2x2_ASAP7_75t_L g763 ( .A(n_591), .B(n_629), .Y(n_763) );
AND2x2_ASAP7_75t_L g788 ( .A(n_591), .B(n_618), .Y(n_788) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g606 ( .A(n_593), .Y(n_606) );
BUFx3_ASAP7_75t_L g648 ( .A(n_593), .Y(n_648) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_593), .Y(n_675) );
INVx1_ASAP7_75t_L g684 ( .A(n_593), .Y(n_684) );
AOI33xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .A3(n_607), .B1(n_608), .B2(n_609), .B3(n_610), .Y(n_599) );
AOI21x1_ASAP7_75t_SL g702 ( .A1(n_600), .A2(n_624), .B(n_686), .Y(n_702) );
INVx2_ASAP7_75t_L g732 ( .A(n_600), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_600), .B(n_731), .Y(n_738) );
AND2x2_ASAP7_75t_L g686 ( .A(n_601), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g649 ( .A(n_604), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g750 ( .A(n_605), .Y(n_750) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_606), .Y(n_740) );
OAI32xp33_ASAP7_75t_L g789 ( .A1(n_607), .A2(n_609), .A3(n_785), .B1(n_790), .B2(n_792), .Y(n_789) );
AND2x2_ASAP7_75t_L g707 ( .A(n_608), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g697 ( .A(n_609), .Y(n_697) );
AND2x2_ASAP7_75t_L g762 ( .A(n_609), .B(n_706), .Y(n_762) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_623), .B1(n_626), .B2(n_640), .C(n_644), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_617), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_618), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_618), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_618), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .C(n_636), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_628), .A2(n_690), .B1(n_730), .B2(n_733), .Y(n_729) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g633 ( .A(n_629), .Y(n_633) );
NOR2x1p5_ASAP7_75t_L g647 ( .A(n_629), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_629), .Y(n_669) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI322xp33_ASAP7_75t_L g696 ( .A1(n_632), .A2(n_674), .A3(n_697), .B1(n_698), .B2(n_699), .C1(n_700), .C2(n_702), .Y(n_696) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_653), .B(n_654), .C(n_656), .Y(n_652) );
OR2x2_ASAP7_75t_L g744 ( .A(n_634), .B(n_698), .Y(n_744) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g651 ( .A(n_635), .B(n_639), .Y(n_651) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g657 ( .A(n_641), .B(n_658), .Y(n_657) );
INVx3_ASAP7_75t_SL g689 ( .A(n_642), .Y(n_689) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_646), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_SL g693 ( .A(n_649), .Y(n_693) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_650), .Y(n_735) );
OR2x6_ASAP7_75t_SL g790 ( .A(n_653), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_658), .A2(n_781), .B(n_782), .C(n_789), .Y(n_780) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_662), .B(n_665), .C(n_669), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_660), .A2(n_672), .B(n_679), .C(n_703), .Y(n_671) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_716), .C(n_760), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_675), .Y(n_767) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g722 ( .A(n_678), .Y(n_722) );
NOR3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_692), .C(n_696), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_688), .B2(n_691), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g724 ( .A(n_684), .Y(n_724) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_684), .Y(n_791) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_SL g777 ( .A(n_690), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OR2x2_ASAP7_75t_L g727 ( .A(n_693), .B(n_713), .Y(n_727) );
OR2x2_ASAP7_75t_L g778 ( .A(n_693), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g776 ( .A(n_701), .Y(n_776) );
OR2x2_ASAP7_75t_L g792 ( .A(n_701), .B(n_731), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B(n_709), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g717 ( .A1(n_704), .A2(n_718), .A3(n_719), .B(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g749 ( .A(n_714), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND4xp25_ASAP7_75t_SL g716 ( .A(n_717), .B(n_725), .C(n_736), .D(n_741), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_724), .Y(n_759) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVxp67_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B1(n_749), .B2(n_751), .C(n_753), .Y(n_741) );
NAND2xp33_ASAP7_75t_SL g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g786 ( .A(n_745), .Y(n_786) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g781 ( .A(n_755), .Y(n_781) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_780), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_764), .B2(n_766), .C(n_770), .Y(n_761) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
AOI21xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_775), .B(n_778), .Y(n_770) );
INVxp33_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B1(n_786), .B2(n_787), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_794), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_812), .Y(n_824) );
XNOR2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .Y(n_812) );
NAND3x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_816), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_820), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
endmodule