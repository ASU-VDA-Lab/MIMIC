module fake_netlist_1_11342_n_680 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_680);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_680;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_621;
wire n_342;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_582;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_19), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_76), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_83), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_55), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_32), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_80), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_73), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_86), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_6), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_35), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_10), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_84), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_12), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_17), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_2), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_57), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_21), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_66), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_22), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_19), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_3), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
BUFx5_ASAP7_75t_L g121 ( .A(n_33), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_23), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_6), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_1), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_112), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_100), .B(n_0), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_103), .B(n_1), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_121), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_102), .Y(n_130) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_92), .A2(n_43), .B(n_82), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_121), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_88), .B(n_2), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_95), .B(n_3), .Y(n_136) );
OAI22x1_ASAP7_75t_R g137 ( .A1(n_87), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_108), .A2(n_44), .B(n_81), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_125), .A2(n_4), .B1(n_5), .B2(n_8), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_120), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_125), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_87), .B(n_9), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_121), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_98), .B(n_11), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_127), .B(n_106), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_145), .B(n_148), .Y(n_159) );
NAND3xp33_ASAP7_75t_L g160 ( .A(n_145), .B(n_97), .C(n_109), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_148), .B(n_90), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
NAND3xp33_ASAP7_75t_L g165 ( .A(n_150), .B(n_113), .C(n_115), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_129), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_150), .B(n_111), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_149), .A2(n_124), .B1(n_119), .B2(n_123), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_152), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_141), .B(n_116), .Y(n_175) );
AOI21x1_ASAP7_75t_L g176 ( .A1(n_132), .A2(n_110), .B(n_117), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_141), .B(n_107), .Y(n_177) );
NAND2xp33_ASAP7_75t_L g178 ( .A(n_138), .B(n_121), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_153), .B(n_154), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_136), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_135), .B(n_107), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_152), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_138), .B(n_152), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_138), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_138), .B(n_121), .Y(n_191) );
INVx5_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_128), .B(n_124), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_168), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_168), .B(n_155), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_181), .B(n_149), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_194), .B(n_128), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_168), .A2(n_136), .B1(n_156), .B2(n_155), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_168), .A2(n_156), .B1(n_155), .B2(n_118), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_183), .B(n_90), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_186), .A2(n_131), .B(n_142), .Y(n_204) );
BUFx12f_ASAP7_75t_L g205 ( .A(n_194), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_170), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_170), .B(n_121), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_170), .A2(n_126), .B1(n_133), .B2(n_146), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_180), .A2(n_119), .B1(n_104), .B2(n_147), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_143), .B1(n_147), .B2(n_93), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_161), .B(n_91), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_158), .B(n_91), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_167), .B(n_93), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_158), .A2(n_143), .B1(n_111), .B2(n_122), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_172), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
AND2x6_ASAP7_75t_SL g222 ( .A(n_175), .B(n_130), .Y(n_222) );
AO221x1_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_137), .B1(n_126), .B2(n_133), .C(n_139), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g224 ( .A1(n_171), .A2(n_137), .B1(n_122), .B2(n_142), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_177), .B(n_101), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_172), .B(n_121), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_175), .B(n_105), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_162), .B(n_126), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_162), .B(n_151), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
BUFx2_ASAP7_75t_R g233 ( .A(n_171), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_160), .B(n_133), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_165), .A2(n_126), .B1(n_133), .B2(n_144), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_165), .B(n_131), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_166), .B(n_126), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_166), .B(n_133), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_195), .B(n_131), .Y(n_239) );
NOR2x1p5_ASAP7_75t_L g240 ( .A(n_191), .B(n_151), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_174), .B(n_133), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
OR2x2_ASAP7_75t_SL g243 ( .A(n_191), .B(n_142), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_192), .Y(n_244) );
AND3x1_ASAP7_75t_L g245 ( .A(n_157), .B(n_12), .C(n_13), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_199), .B(n_173), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g247 ( .A(n_233), .B(n_182), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_208), .B(n_188), .Y(n_248) );
CKINVDCx8_ASAP7_75t_R g249 ( .A(n_222), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_204), .A2(n_173), .B(n_184), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_236), .A2(n_195), .B(n_188), .Y(n_251) );
AND3x4_ASAP7_75t_L g252 ( .A(n_224), .B(n_179), .C(n_185), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_242), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_223), .A2(n_151), .B1(n_146), .B2(n_139), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_239), .A2(n_184), .B(n_178), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_187), .B(n_142), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_198), .A2(n_187), .B(n_131), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_200), .B(n_182), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_200), .B(n_182), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_212), .B(n_182), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_201), .B(n_185), .Y(n_261) );
AOI33xp33_ASAP7_75t_L g262 ( .A1(n_210), .A2(n_193), .A3(n_190), .B1(n_189), .B2(n_169), .B3(n_164), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_217), .B(n_185), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_232), .A2(n_193), .B(n_190), .C(n_189), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_207), .A2(n_179), .B(n_163), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_207), .A2(n_179), .B(n_163), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_227), .A2(n_193), .B(n_157), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_163), .B(n_190), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_219), .A2(n_151), .B1(n_140), .B2(n_144), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_239), .A2(n_189), .B(n_169), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_205), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_228), .B(n_139), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_220), .A2(n_169), .B(n_164), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_221), .A2(n_151), .B(n_146), .C(n_144), .Y(n_275) );
O2A1O1Ixp5_ASAP7_75t_L g276 ( .A1(n_231), .A2(n_164), .B(n_192), .C(n_151), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_202), .B(n_139), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_197), .A2(n_146), .B1(n_144), .B2(n_140), .Y(n_278) );
OAI21xp33_ASAP7_75t_L g279 ( .A1(n_211), .A2(n_139), .B(n_140), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_197), .B(n_140), .Y(n_280) );
AOI21x1_ASAP7_75t_L g281 ( .A1(n_231), .A2(n_192), .B(n_146), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_213), .A2(n_221), .B1(n_206), .B2(n_245), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_205), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_203), .B(n_14), .Y(n_284) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_216), .B(n_14), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_213), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_213), .A2(n_146), .B1(n_144), .B2(n_140), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_223), .A2(n_144), .B(n_140), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_218), .A2(n_15), .B(n_16), .C(n_17), .Y(n_289) );
NAND2xp33_ASAP7_75t_L g290 ( .A(n_206), .B(n_192), .Y(n_290) );
O2A1O1Ixp5_ASAP7_75t_L g291 ( .A1(n_234), .A2(n_192), .B(n_52), .C(n_54), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_229), .A2(n_48), .B(n_79), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_226), .B(n_15), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_250), .A2(n_237), .B(n_241), .Y(n_295) );
AOI221x1_ASAP7_75t_L g296 ( .A1(n_282), .A2(n_196), .B1(n_214), .B2(n_234), .C(n_238), .Y(n_296) );
AO31x2_ASAP7_75t_L g297 ( .A1(n_275), .A2(n_243), .A3(n_215), .B(n_214), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_292), .A2(n_209), .B(n_240), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_SL g299 ( .A1(n_275), .A2(n_244), .B(n_230), .C(n_215), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_283), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_286), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_256), .A2(n_196), .B(n_214), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_257), .A2(n_196), .B(n_214), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_286), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_271), .A2(n_234), .B(n_235), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_248), .A2(n_243), .B1(n_244), .B2(n_230), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_251), .A2(n_244), .B(n_230), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_258), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_247), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_253), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_267), .B(n_225), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_253), .B(n_225), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_292), .A2(n_225), .B(n_51), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_246), .A2(n_225), .B1(n_18), .B2(n_20), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_265), .A2(n_47), .B(n_78), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_266), .A2(n_46), .B(n_77), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_246), .A2(n_16), .B1(n_18), .B2(n_20), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_252), .B(n_24), .Y(n_320) );
NAND3xp33_ASAP7_75t_SL g321 ( .A(n_249), .B(n_252), .C(n_289), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_26), .B(n_27), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_284), .B(n_28), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_267), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_284), .B(n_31), .C(n_34), .D(n_36), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_273), .A2(n_38), .B(n_39), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_277), .Y(n_327) );
AO31x2_ASAP7_75t_L g328 ( .A1(n_278), .A2(n_40), .A3(n_41), .B(n_42), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_288), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_274), .A2(n_45), .B(n_56), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_254), .B(n_58), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_300), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_302), .A2(n_254), .B(n_291), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_303), .A2(n_255), .B(n_280), .Y(n_334) );
OA21x2_ASAP7_75t_L g335 ( .A1(n_296), .A2(n_293), .B(n_279), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_299), .A2(n_264), .B(n_290), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_314), .A2(n_276), .B(n_269), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_323), .A2(n_268), .B(n_261), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_308), .B(n_262), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_318), .A2(n_262), .B(n_270), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_312), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_327), .B(n_306), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_295), .A2(n_287), .B(n_285), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_313), .B(n_263), .Y(n_346) );
AO31x2_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_315), .A3(n_320), .B(n_319), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_322), .A2(n_288), .B(n_260), .Y(n_348) );
INVx5_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_297), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_301), .B(n_59), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_301), .B(n_61), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_304), .B(n_62), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_305), .A2(n_63), .B(n_64), .Y(n_356) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_331), .A2(n_67), .B(n_68), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_304), .B(n_69), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
AO31x2_ASAP7_75t_L g360 ( .A1(n_330), .A2(n_85), .A3(n_71), .B(n_72), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_359), .A2(n_317), .B(n_316), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_352), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_359), .A2(n_326), .B(n_321), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_350), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_355), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_349), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_355), .B(n_312), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_341), .B(n_309), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_334), .A2(n_297), .B(n_329), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_325), .B1(n_324), .B2(n_328), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_333), .A2(n_345), .B(n_338), .Y(n_379) );
AOI21x1_ASAP7_75t_L g380 ( .A1(n_335), .A2(n_325), .B(n_328), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_347), .B(n_324), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_347), .B(n_324), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_348), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_70), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_333), .A2(n_74), .B(n_345), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_367), .B(n_347), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_372), .B(n_332), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_372), .B(n_354), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_371), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_387), .B(n_347), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_384), .B(n_354), .Y(n_395) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_376), .B(n_343), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_364), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_384), .B(n_343), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_385), .B(n_343), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_367), .B(n_347), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_387), .B(n_347), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_389), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_364), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_365), .B(n_344), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_387), .B(n_344), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_369), .B(n_351), .Y(n_418) );
INVx3_ASAP7_75t_SL g419 ( .A(n_369), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_362), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_381), .B(n_356), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_385), .B(n_343), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g425 ( .A(n_369), .B(n_349), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_357), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_366), .B(n_358), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_425), .B(n_369), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_394), .B(n_381), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_394), .B(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_397), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_405), .B(n_382), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_405), .B(n_382), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_391), .B(n_383), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_419), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_426), .B(n_368), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_409), .B(n_362), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_426), .B(n_377), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g444 ( .A(n_425), .B(n_369), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_423), .B(n_377), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_423), .B(n_377), .Y(n_448) );
NOR2x1p5_ASAP7_75t_L g449 ( .A(n_406), .B(n_383), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_414), .B(n_377), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_423), .B(n_368), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_393), .B(n_366), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_423), .B(n_368), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_390), .B(n_368), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_403), .B(n_373), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_390), .B(n_373), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_373), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_397), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_414), .A2(n_389), .B1(n_370), .B2(n_374), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_404), .B(n_373), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_412), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_411), .B(n_373), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_416), .B(n_422), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_411), .B(n_386), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_422), .B(n_386), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_413), .B(n_421), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_413), .B(n_386), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_408), .B(n_383), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_413), .B(n_386), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_417), .B(n_379), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_396), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_454), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_430), .B(n_406), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_454), .B(n_408), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_429), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_430), .B(n_417), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_430), .B(n_406), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_429), .Y(n_490) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_466), .A2(n_392), .B(n_420), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_431), .B(n_421), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_431), .B(n_436), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_436), .B(n_406), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_420), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_462), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_432), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_437), .B(n_420), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_470), .B(n_424), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_453), .B(n_421), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_432), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_440), .B(n_420), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_453), .B(n_400), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_482), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_440), .B(n_379), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_449), .B(n_370), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_433), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_439), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_434), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_459), .B(n_427), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_443), .B(n_379), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_470), .B(n_399), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_434), .B(n_395), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_441), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_427), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_451), .B(n_370), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_460), .B(n_396), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_443), .B(n_379), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_447), .B(n_418), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_446), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_445), .B(n_379), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_457), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_457), .Y(n_529) );
O2A1O1Ixp5_ASAP7_75t_L g530 ( .A1(n_447), .A2(n_374), .B(n_383), .C(n_353), .Y(n_530) );
OR2x6_ASAP7_75t_L g531 ( .A(n_481), .B(n_370), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_450), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_446), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_463), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_449), .B(n_370), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_460), .B(n_396), .Y(n_537) );
INVx3_ASAP7_75t_R g538 ( .A(n_458), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_445), .B(n_379), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_445), .B(n_363), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_467), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_468), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_529), .B(n_481), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_535), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_542), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_543), .B(n_460), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_543), .B(n_472), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_493), .B(n_448), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_487), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_531), .A2(n_481), .B1(n_457), .B2(n_439), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_468), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_491), .A2(n_452), .B1(n_455), .B2(n_448), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_525), .B(n_456), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_525), .B(n_456), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_493), .B(n_448), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_530), .A2(n_531), .B(n_528), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_R g559 ( .A1(n_538), .A2(n_456), .B(n_455), .C(n_452), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_517), .B(n_472), .Y(n_560) );
NAND2x1_ASAP7_75t_L g561 ( .A(n_528), .B(n_461), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_517), .B(n_458), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_494), .B(n_452), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_483), .B(n_467), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_496), .B(n_428), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_507), .B(n_469), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_490), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_499), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_507), .B(n_469), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_488), .B(n_471), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_494), .B(n_455), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_514), .B(n_480), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_495), .B(n_478), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_510), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_509), .B(n_475), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g578 ( .A(n_511), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_495), .B(n_478), .Y(n_579) );
INVxp33_ASAP7_75t_L g580 ( .A(n_486), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_500), .B(n_478), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_500), .B(n_478), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_484), .B(n_471), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_513), .B(n_473), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_502), .Y(n_585) );
OAI22xp33_ASAP7_75t_SL g586 ( .A1(n_531), .A2(n_444), .B1(n_428), .B2(n_389), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_514), .B(n_480), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_524), .B(n_480), .Y(n_588) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_531), .B(n_465), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_501), .A2(n_353), .B(n_358), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_485), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_484), .B(n_479), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_512), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_513), .B(n_473), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_554), .A2(n_516), .B1(n_489), .B2(n_504), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_558), .A2(n_515), .B1(n_537), .B2(n_523), .C(n_506), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_548), .B(n_566), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_550), .B(n_489), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_562), .B(n_524), .Y(n_599) );
OAI32xp33_ASAP7_75t_L g600 ( .A1(n_578), .A2(n_428), .A3(n_444), .B1(n_520), .B2(n_519), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_586), .A2(n_509), .B(n_536), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_544), .B(n_552), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_591), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_548), .B(n_522), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_566), .B(n_539), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_552), .A2(n_504), .B1(n_536), .B2(n_509), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_569), .B(n_539), .Y(n_611) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_585), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_544), .A2(n_536), .B1(n_444), .B2(n_428), .Y(n_613) );
OAI322xp33_ASAP7_75t_L g614 ( .A1(n_555), .A2(n_505), .A3(n_533), .B1(n_532), .B2(n_518), .C1(n_540), .C2(n_527), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_589), .B(n_527), .Y(n_615) );
OAI321xp33_ASAP7_75t_L g616 ( .A1(n_559), .A2(n_569), .A3(n_549), .B1(n_556), .B2(n_444), .C(n_540), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_577), .B(n_534), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_584), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g619 ( .A1(n_580), .A2(n_363), .B(n_526), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_560), .A2(n_534), .B1(n_526), .B2(n_521), .C(n_498), .Y(n_620) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_594), .A2(n_573), .B(n_588), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_583), .B(n_521), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_561), .A2(n_442), .B(n_482), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_546), .A2(n_442), .B1(n_497), .B2(n_485), .C(n_498), .Y(n_625) );
BUFx3_ASAP7_75t_L g626 ( .A(n_577), .Y(n_626) );
O2A1O1Ixp5_ASAP7_75t_L g627 ( .A1(n_547), .A2(n_593), .B(n_551), .C(n_567), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_596), .A2(n_553), .B1(n_571), .B2(n_588), .C(n_587), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_612), .A2(n_573), .B1(n_587), .B2(n_557), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_616), .A2(n_582), .B(n_581), .C(n_579), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_606), .A2(n_575), .B1(n_572), .B2(n_563), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_603), .B(n_592), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_626), .B(n_576), .Y(n_634) );
OAI321xp33_ASAP7_75t_L g635 ( .A1(n_613), .A2(n_574), .A3(n_570), .B1(n_380), .B2(n_497), .C(n_479), .Y(n_635) );
OAI32xp33_ASAP7_75t_L g636 ( .A1(n_613), .A2(n_383), .A3(n_590), .B1(n_465), .B2(n_461), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_614), .A2(n_590), .B1(n_475), .B2(n_479), .C(n_477), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_621), .A2(n_477), .B1(n_476), .B2(n_465), .C(n_461), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_595), .A2(n_363), .B1(n_476), .B2(n_461), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_608), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_601), .B(n_465), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_610), .A2(n_363), .B1(n_357), .B2(n_474), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_602), .B(n_363), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_608), .Y(n_644) );
OAI322xp33_ASAP7_75t_SL g645 ( .A1(n_597), .A2(n_474), .A3(n_464), .B1(n_375), .B2(n_378), .C1(n_346), .C2(n_380), .Y(n_645) );
OAI322xp33_ASAP7_75t_SL g646 ( .A1(n_597), .A2(n_474), .A3(n_464), .B1(n_378), .B2(n_346), .C1(n_380), .C2(n_360), .Y(n_646) );
OAI22xp33_ASAP7_75t_SL g647 ( .A1(n_604), .A2(n_349), .B1(n_464), .B2(n_336), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_605), .A2(n_357), .B1(n_356), .B2(n_349), .Y(n_648) );
AOI321xp33_ASAP7_75t_L g649 ( .A1(n_600), .A2(n_342), .A3(n_336), .B1(n_338), .B2(n_360), .C(n_357), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_627), .A2(n_342), .B1(n_356), .B2(n_361), .C(n_360), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_619), .A2(n_356), .B(n_361), .C(n_335), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_625), .A2(n_345), .B(n_361), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_620), .B(n_335), .C(n_348), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_619), .B(n_360), .C(n_388), .D(n_361), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_623), .B(n_628), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_624), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_618), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_599), .A2(n_611), .B1(n_609), .B2(n_622), .C(n_607), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_615), .B(n_388), .C(n_333), .Y(n_659) );
AOI221x1_ASAP7_75t_L g660 ( .A1(n_615), .A2(n_360), .B1(n_361), .B2(n_388), .C(n_348), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g661 ( .A1(n_656), .A2(n_631), .A3(n_633), .B1(n_637), .B2(n_644), .C1(n_640), .C2(n_657), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_635), .B(n_632), .C(n_647), .Y(n_662) );
AND4x1_ASAP7_75t_L g663 ( .A(n_638), .B(n_642), .C(n_650), .D(n_639), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_649), .B(n_629), .C(n_636), .D(n_630), .Y(n_664) );
OAI211xp5_ASAP7_75t_L g665 ( .A1(n_643), .A2(n_654), .B(n_658), .C(n_648), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_653), .B(n_655), .C(n_660), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_661), .B(n_634), .Y(n_667) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_664), .B(n_652), .C(n_641), .D(n_635), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_662), .B(n_659), .C(n_651), .D(n_646), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_665), .B(n_645), .C(n_617), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_668), .Y(n_671) );
NAND2xp33_ASAP7_75t_L g672 ( .A(n_670), .B(n_666), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_671), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_672), .B(n_667), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_674), .A2(n_669), .B1(n_617), .B2(n_663), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_675), .B(n_673), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_598), .B1(n_348), .B2(n_335), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_677), .A2(n_360), .B(n_348), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_337), .B(n_335), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_679), .A2(n_337), .B1(n_360), .B2(n_671), .Y(n_680) );
endmodule