module real_jpeg_26962_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_323, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_323;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_0),
.B(n_198),
.Y(n_203)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_52),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_52),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_43),
.B1(n_45),
.B2(n_109),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_4),
.A2(n_22),
.B1(n_26),
.B2(n_109),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_109),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_6),
.A2(n_22),
.B1(n_26),
.B2(n_58),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_58),
.Y(n_278)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_34),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_56),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_74),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_34),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_10),
.B(n_22),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_25),
.B(n_28),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_38),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_84),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_82),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_76),
.Y(n_14)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.C(n_69),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_16),
.A2(n_17),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_53),
.Y(n_17)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_18),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_18),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_18),
.A2(n_111),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_18),
.B(n_35),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_19),
.A2(n_102),
.B(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_20),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_20),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_20),
.B(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_22),
.A2(n_24),
.B(n_34),
.C(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_27),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_27),
.B(n_33),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_31),
.B(n_34),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_31),
.A2(n_169),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_34),
.A2(n_43),
.B(n_157),
.C(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_34),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_46),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_36),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_41),
.B(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_37),
.A2(n_47),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_43),
.B(n_49),
.C(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_38),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_38),
.B(n_51),
.Y(n_144)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_40),
.Y(n_157)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_42),
.B(n_48),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_45),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_43),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_45),
.B(n_61),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_48),
.B(n_115),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_48),
.A2(n_262),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_53),
.A2(n_54),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_59),
.B(n_60),
.C(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_59),
.A2(n_65),
.B(n_80),
.Y(n_286)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_63),
.B(n_107),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_65),
.B(n_80),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_67),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_67),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_67),
.A2(n_69),
.B1(n_246),
.B2(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_73),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_78),
.B(n_120),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_314),
.B(n_320),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_290),
.A3(n_309),
.B1(n_312),
.B2(n_313),
.C(n_323),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_270),
.B(n_289),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_250),
.B(n_269),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_150),
.B(n_232),
.C(n_249),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_136),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_90),
.B(n_136),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_116),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_92),
.B(n_105),
.C(n_116),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_93),
.B(n_101),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B(n_99),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_95),
.A2(n_96),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_95),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_96),
.B(n_149),
.Y(n_196)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_99),
.B(n_197),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_102),
.B(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_104),
.B(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_112),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_110),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_111),
.B(n_294),
.C(n_299),
.Y(n_308)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_118),
.B(n_123),
.C(n_126),
.Y(n_247)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_133),
.B(n_196),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_134),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_137),
.A2(n_138),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_144),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_148),
.B(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_231),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_224),
.B(n_230),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_181),
.B(n_223),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_154),
.B(n_170),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.C(n_165),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_155),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_159),
.A2(n_160),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_159),
.B(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_159),
.A2(n_160),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_160),
.A2(n_281),
.B(n_286),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_221)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_164),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_169),
.B(n_178),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_177),
.C(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_218),
.B(n_222),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_199),
.B(n_217),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_216),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_201),
.B(n_204),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_210),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_247),
.B2(n_248),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_241),
.C(n_248),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_252),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_268),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_264),
.B2(n_265),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_265),
.C(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_258),
.C(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_272),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_287),
.B2(n_288),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_280),
.C(n_288),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B(n_279),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_292),
.C(n_301),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_279),
.B(n_292),
.CI(n_301),
.CON(n_311),
.SN(n_311)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_302),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_294),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_304),
.C(n_308),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);


endmodule