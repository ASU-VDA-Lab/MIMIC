module fake_jpeg_26815_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_47),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_31),
.B1(n_21),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_78),
.B1(n_18),
.B2(n_37),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_46),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_76),
.B(n_99),
.CI(n_18),
.CON(n_120),
.SN(n_120)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_31),
.B1(n_21),
.B2(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_31),
.B1(n_21),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_100),
.B1(n_18),
.B2(n_37),
.Y(n_103)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_89),
.Y(n_118)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_92),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_47),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_12),
.C(n_16),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_61),
.B1(n_34),
.B2(n_33),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_23),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_21),
.B1(n_31),
.B2(n_29),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_24),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_76),
.B1(n_75),
.B2(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_100),
.B1(n_52),
.B2(n_58),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_62),
.B1(n_43),
.B2(n_45),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_55),
.C(n_46),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_126),
.C(n_97),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_43),
.B1(n_51),
.B2(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_112),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_33),
.B(n_34),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_27),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_23),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_46),
.C(n_41),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_49),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_88),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_48),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_91),
.C(n_79),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_114),
.C(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_138),
.Y(n_171)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_143),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_7),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_83),
.B1(n_105),
.B2(n_109),
.Y(n_174)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_156),
.Y(n_186)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_92),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_73),
.B1(n_101),
.B2(n_121),
.Y(n_177)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_123),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_159),
.Y(n_187)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_124),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_86),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_7),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_16),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_44),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_98),
.B1(n_101),
.B2(n_111),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_177),
.B1(n_157),
.B2(n_147),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_148),
.B(n_152),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_167),
.B(n_33),
.Y(n_207)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_178),
.C(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_103),
.A3(n_117),
.B1(n_35),
.B2(n_111),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_83),
.B1(n_105),
.B2(n_26),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_145),
.C(n_146),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_183),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_121),
.C(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_189),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_48),
.C(n_30),
.Y(n_224)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_44),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_194),
.A2(n_213),
.B1(n_221),
.B2(n_170),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_158),
.A3(n_138),
.B1(n_136),
.B2(n_152),
.C1(n_150),
.C2(n_133),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_201),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_159),
.B(n_136),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_200),
.B(n_209),
.C(n_28),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_157),
.B(n_147),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_142),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_214),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_17),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_48),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_210),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_172),
.B1(n_19),
.B2(n_2),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_135),
.B(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_220),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_166),
.A2(n_27),
.B1(n_26),
.B2(n_30),
.Y(n_213)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_26),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_72),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_184),
.B(n_19),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_223),
.C(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_242),
.C(n_249),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_235),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_250),
.B1(n_209),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_186),
.B1(n_187),
.B2(n_184),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_240),
.B1(n_246),
.B2(n_248),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_187),
.B1(n_180),
.B2(n_170),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_191),
.C(n_185),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_213),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_30),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_214),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_210),
.B1(n_198),
.B2(n_207),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_48),
.C(n_24),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_253),
.B1(n_257),
.B2(n_260),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_199),
.B1(n_220),
.B2(n_193),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_199),
.B1(n_200),
.B2(n_217),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_241),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_268),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_224),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_258),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_194),
.B1(n_217),
.B2(n_212),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_202),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_204),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_250),
.B1(n_240),
.B2(n_248),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_212),
.B1(n_222),
.B2(n_221),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_17),
.B1(n_28),
.B2(n_0),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_9),
.B(n_16),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_8),
.B(n_15),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_227),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_226),
.C(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_274),
.C(n_276),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_231),
.C(n_241),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_281),
.B(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_244),
.C(n_249),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_228),
.C(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_24),
.C(n_17),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_19),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_17),
.C(n_28),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_292),
.B(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_263),
.B1(n_260),
.B2(n_257),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_293),
.A2(n_265),
.B1(n_276),
.B2(n_2),
.Y(n_311)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_6),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_262),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_301),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_255),
.B(n_270),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_282),
.B(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_272),
.C(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_311),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_290),
.C(n_301),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_312),
.C(n_315),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_314),
.B(n_298),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_300),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_294),
.A2(n_5),
.B1(n_10),
.B2(n_2),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_8),
.C(n_10),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_8),
.C(n_10),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_302),
.C(n_304),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_322),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_307),
.B(n_313),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_321),
.B(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_321),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_296),
.B(n_302),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_298),
.A3(n_293),
.B1(n_3),
.B2(n_4),
.C1(n_9),
.C2(n_13),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_296),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_295),
.B(n_294),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_331),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_327),
.C(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.C(n_330),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_3),
.B1(n_13),
.B2(n_0),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_13),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_1),
.Y(n_342)
);


endmodule