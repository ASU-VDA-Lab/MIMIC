module real_jpeg_26891_n_17 (n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_1),
.A2(n_45),
.B1(n_97),
.B2(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_45),
.B1(n_156),
.B2(n_162),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_63),
.B1(n_97),
.B2(n_98),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_2),
.A2(n_63),
.B1(n_156),
.B2(n_162),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_4),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_114),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_97),
.B1(n_98),
.B2(n_114),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_114),
.B1(n_156),
.B2(n_162),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_6),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_152),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_97),
.B1(n_98),
.B2(n_152),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_6),
.A2(n_152),
.B1(n_156),
.B2(n_162),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_8),
.A2(n_56),
.B1(n_97),
.B2(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_56),
.B1(n_156),
.B2(n_162),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_9),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_9),
.A2(n_34),
.B1(n_36),
.B2(n_215),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_9),
.A2(n_97),
.B1(n_98),
.B2(n_215),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_9),
.A2(n_156),
.B1(n_162),
.B2(n_215),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_10),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_34),
.B1(n_36),
.B2(n_135),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_10),
.A2(n_97),
.B1(n_98),
.B2(n_135),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_10),
.A2(n_135),
.B1(n_156),
.B2(n_162),
.Y(n_287)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_30),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_36),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_35),
.B(n_36),
.C(n_39),
.D(n_43),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_60),
.B(n_64),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_97),
.B(n_99),
.C(n_100),
.D(n_104),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_12),
.B(n_97),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_98),
.B(n_132),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_12),
.A2(n_81),
.B1(n_156),
.B2(n_162),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_196),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_13),
.A2(n_97),
.B1(n_98),
.B2(n_196),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_13),
.A2(n_156),
.B1(n_162),
.B2(n_196),
.Y(n_319)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_324),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_311),
.B(n_323),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_275),
.A3(n_304),
.B1(n_309),
.B2(n_310),
.C(n_332),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_225),
.A3(n_264),
.B1(n_269),
.B2(n_274),
.C(n_333),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_176),
.C(n_221),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_143),
.B(n_175),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_119),
.B(n_142),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_92),
.B(n_118),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_68),
.B(n_91),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_47),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_27),
.B(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_38),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_29),
.B(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2x1_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_34),
.B(n_103),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_40),
.Y(n_41)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_36),
.A2(n_98),
.A3(n_99),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_39),
.A2(n_42),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_39),
.A2(n_42),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_39),
.A2(n_42),
.B1(n_241),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_43),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_46),
.A2(n_57),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_46),
.A2(n_139),
.B1(n_174),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_46),
.A2(n_139),
.B1(n_198),
.B2(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_46),
.A2(n_139),
.B(n_250),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_59),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_51),
.A2(n_100),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_51),
.A2(n_100),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_51),
.A2(n_100),
.B1(n_253),
.B2(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_51),
.A2(n_100),
.B(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_55),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_60),
.A2(n_76),
.B1(n_113),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_60),
.A2(n_61),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_60),
.A2(n_195),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_60),
.A2(n_76),
.B(n_214),
.Y(n_243)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_81),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_84),
.B(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g213 ( 
.A(n_67),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_78),
.B(n_90),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_77),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_76),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_73),
.A2(n_75),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_89),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_129),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_131),
.B(n_155),
.C(n_156),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_107),
.C(n_110),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_98),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_106),
.A2(n_125),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_106),
.A2(n_184),
.B1(n_210),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_106),
.A2(n_184),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_109),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_121),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_136),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_137),
.C(n_138),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.C(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_129),
.A2(n_188),
.B(n_190),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_129),
.A2(n_190),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_129),
.A2(n_232),
.B1(n_260),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_129),
.A2(n_232),
.B1(n_287),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_160),
.B1(n_189),
.B2(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_130),
.A2(n_160),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_130),
.A2(n_160),
.B1(n_319),
.B2(n_328),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_132),
.B1(n_156),
.B2(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_158),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_148),
.C(n_158),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_157),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_169),
.C(n_172),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_163),
.B(n_164),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_177),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_200),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_178),
.B(n_200),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_192),
.C(n_199),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_182),
.C(n_191),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_191),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B(n_186),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_199),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_197),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_211),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_211),
.C(n_220),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_206),
.C(n_208),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_223),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_245),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_245),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.C(n_244),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_237),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_236),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_243),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_243),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_243),
.A2(n_258),
.B(n_261),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_263),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_255),
.B1(n_256),
.B2(n_262),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_251),
.B(n_254),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_251),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_254),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_277),
.B1(n_278),
.B2(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_262),
.C(n_263),
.Y(n_305)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_270),
.B(n_273),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_292),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_289),
.C(n_290),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_286),
.B2(n_288),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_281),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_285),
.C(n_286),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_282),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_285),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_296),
.C(n_300),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_288),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_295),
.C(n_303),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_291),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_303),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_322),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_315),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_329),
.Y(n_330)
);


endmodule