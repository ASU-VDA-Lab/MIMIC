module fake_jpeg_29541_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_39),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_9),
.Y(n_81)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_37),
.B1(n_1),
.B2(n_3),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_74),
.B(n_77),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_0),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_17),
.C(n_32),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_12),
.B(n_13),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_6),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_63),
.B(n_7),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_63),
.B1(n_10),
.B2(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_88),
.B1(n_86),
.B2(n_79),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_15),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_75),
.B1(n_68),
.B2(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_89),
.C(n_84),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_18),
.C(n_20),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_92),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_98),
.B(n_80),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_23),
.C(n_24),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_34),
.B(n_25),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_26),
.Y(n_106)
);


endmodule