module fake_jpeg_10206_n_302 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_33;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_31),
.B1(n_26),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_49),
.B1(n_65),
.B2(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_70),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_21),
.B1(n_45),
.B2(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_83),
.B1(n_91),
.B2(n_34),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_0),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_34),
.A3(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_93),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_0),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_102),
.B1(n_93),
.B2(n_51),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_106),
.Y(n_123)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_54),
.B1(n_64),
.B2(n_67),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_51),
.B1(n_18),
.B2(n_28),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_59),
.B1(n_46),
.B2(n_48),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_1),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_115),
.B(n_88),
.Y(n_126)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_30),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_79),
.B1(n_91),
.B2(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_79),
.B1(n_76),
.B2(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_46),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_79),
.C(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_118),
.B1(n_72),
.B2(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_121),
.B1(n_130),
.B2(n_136),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_76),
.B1(n_75),
.B2(n_84),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_115),
.A3(n_104),
.B1(n_107),
.B2(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_129),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_144),
.B(n_101),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_93),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_84),
.B1(n_73),
.B2(n_82),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_170)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_142),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_73),
.B1(n_82),
.B2(n_72),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_78),
.B1(n_93),
.B2(n_29),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_105),
.B1(n_95),
.B2(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_22),
.B1(n_33),
.B2(n_29),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_118),
.B1(n_113),
.B2(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_51),
.B1(n_52),
.B2(n_22),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_110),
.B(n_115),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_155),
.B(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_148),
.Y(n_189)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_161),
.B(n_127),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_150),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_128),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_103),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_170),
.B1(n_144),
.B2(n_137),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_99),
.C(n_94),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_160),
.C(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_27),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_30),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_1),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_13),
.C(n_16),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_30),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_27),
.C(n_18),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_139),
.C(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_129),
.B1(n_125),
.B2(n_132),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_188),
.B1(n_9),
.B2(n_15),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_161),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_171),
.B(n_152),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_187),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_196),
.C(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_186),
.B1(n_195),
.B2(n_9),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_168),
.B1(n_167),
.B2(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_140),
.B1(n_128),
.B2(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_148),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_28),
.B(n_24),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_194),
.B1(n_170),
.B2(n_162),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_24),
.B(n_25),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_158),
.C(n_159),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_211),
.B1(n_217),
.B2(n_175),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_218),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_154),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_162),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_215),
.C(n_174),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_181),
.B1(n_195),
.B2(n_182),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_3),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_10),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_10),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_174),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_221),
.B(n_194),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_196),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_178),
.C(n_176),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_226),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_188),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_210),
.B1(n_172),
.B2(n_208),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_217),
.B1(n_211),
.B2(n_235),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_189),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_233),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_198),
.CI(n_209),
.CON(n_245),
.SN(n_245)
);

NAND2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_230),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_212),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_185),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.C(n_252),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_198),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_214),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_193),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_233),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_11),
.B(n_15),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_224),
.C(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_221),
.C(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_236),
.C(n_208),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_258),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_245),
.B1(n_247),
.B2(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_273),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_261),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_243),
.B1(n_244),
.B2(n_6),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_256),
.B(n_265),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_4),
.Y(n_277)
);

OR2x2_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_12),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_10),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_275),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_259),
.B(n_267),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_277),
.B(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_274),
.B(n_263),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_274),
.B(n_11),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_8),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_11),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_290),
.C(n_12),
.Y(n_298)
);

OAI221xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.C(n_5),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_297),
.B(n_14),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_4),
.Y(n_302)
);


endmodule