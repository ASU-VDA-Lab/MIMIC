module fake_jpeg_12607_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_27),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_9),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_86),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_66),
.Y(n_105)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_74),
.B1(n_63),
.B2(n_54),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_99),
.B1(n_100),
.B2(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_72),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_97),
.B(n_53),
.C(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_74),
.B1(n_64),
.B2(n_79),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_69),
.B1(n_57),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_64),
.B1(n_59),
.B2(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_67),
.B1(n_65),
.B2(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_115),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_60),
.B(n_58),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_11),
.B(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_116),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_118),
.B2(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_56),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_77),
.B(n_75),
.C(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_55),
.B1(n_75),
.B2(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_23),
.B1(n_50),
.B2(n_47),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_1),
.B(n_2),
.C(n_5),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_1),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_16),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_137),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_20),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_18),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_19),
.B(n_21),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_52),
.B(n_136),
.Y(n_155)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_155),
.B(n_162),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_130),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_151),
.B(n_162),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_169),
.B(n_164),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_158),
.C(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_131),
.B1(n_146),
.B2(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_166),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_177),
.C(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_159),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_175),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_146),
.Y(n_184)
);


endmodule