module fake_jpeg_26490_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_25),
.B1(n_32),
.B2(n_36),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_53),
.B1(n_40),
.B2(n_58),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_25),
.B1(n_36),
.B2(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_68),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_70),
.B(n_73),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_25),
.B1(n_41),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_93),
.B1(n_96),
.B2(n_26),
.Y(n_117)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_46),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_26),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_85),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_76),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_45),
.B1(n_34),
.B2(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_97),
.B1(n_98),
.B2(n_23),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_39),
.C(n_44),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_23),
.Y(n_133)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_22),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_87),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_37),
.B1(n_44),
.B2(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_27),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_29),
.B1(n_17),
.B2(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_45),
.B1(n_42),
.B2(n_39),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_42),
.B(n_39),
.C(n_37),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_50),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_100),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_37),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_78),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_62),
.B1(n_72),
.B2(n_83),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_98),
.B(n_93),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_94),
.B1(n_69),
.B2(n_66),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_33),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_129),
.B(n_21),
.C(n_35),
.D(n_26),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_118),
.B1(n_124),
.B2(n_119),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_R g129 ( 
.A1(n_74),
.A2(n_24),
.B(n_35),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_18),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_134),
.B(n_141),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_138),
.B(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_147),
.B1(n_148),
.B2(n_128),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_105),
.B1(n_35),
.B2(n_19),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_92),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_103),
.B1(n_63),
.B2(n_64),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_146),
.B1(n_155),
.B2(n_113),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_104),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_87),
.B1(n_102),
.B2(n_81),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_121),
.B1(n_120),
.B2(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_21),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_21),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_23),
.B(n_21),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_154),
.B(n_159),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_115),
.B(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_84),
.B1(n_26),
.B2(n_31),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_80),
.B1(n_76),
.B2(n_12),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_107),
.B1(n_113),
.B2(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_35),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_18),
.B(n_3),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_11),
.C(n_15),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_21),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_116),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_124),
.B1(n_119),
.B2(n_107),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_158),
.C(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_175),
.C(n_142),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_177),
.B1(n_136),
.B2(n_147),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_109),
.C(n_116),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_35),
.A3(n_24),
.B1(n_19),
.B2(n_18),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_1),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_1),
.B(n_2),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_190),
.B(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_24),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_187),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_23),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_19),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_159),
.Y(n_211)
);

XOR2x2_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_158),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_199),
.B(n_201),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_173),
.B1(n_171),
.B2(n_164),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_166),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_177),
.B1(n_185),
.B2(n_183),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_150),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_209),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_149),
.B(n_135),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_138),
.C(n_155),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.C(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_175),
.C(n_188),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_168),
.B1(n_167),
.B2(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_212),
.B1(n_7),
.B2(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_164),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_231),
.C(n_214),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_172),
.B(n_182),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_173),
.B1(n_171),
.B2(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_222),
.B1(n_228),
.B2(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_181),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_207),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_176),
.B1(n_182),
.B2(n_190),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_197),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_191),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_204),
.C(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_244),
.C(n_246),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_195),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_199),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_202),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_215),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_252),
.CI(n_240),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_232),
.C(n_209),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_220),
.B1(n_234),
.B2(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_233),
.B1(n_229),
.B2(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_230),
.B(n_222),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_230),
.B(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_248),
.B(n_223),
.Y(n_262)
);

OAI221xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_264),
.B1(n_238),
.B2(n_246),
.C(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_192),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_213),
.B1(n_219),
.B2(n_212),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_236),
.B(n_228),
.CI(n_232),
.CON(n_264),
.SN(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_237),
.C(n_239),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_272),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_219),
.B1(n_249),
.B2(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_256),
.C(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_263),
.Y(n_277)
);

XOR2x2_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_258),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.C(n_265),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_255),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_266),
.C(n_256),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_271),
.C(n_261),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_262),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_292),
.B(n_282),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_285),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_289),
.B(n_284),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_280),
.B(n_273),
.C(n_258),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_260),
.B(n_254),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_268),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_264),
.A3(n_7),
.B1(n_6),
.B2(n_9),
.C(n_13),
.Y(n_298)
);


endmodule