module fake_jpeg_16276_n_371 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_41),
.Y(n_118)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_45),
.B(n_52),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_59),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_6),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_62),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_5),
.C(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_68),
.Y(n_114)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_79),
.B1(n_85),
.B2(n_97),
.Y(n_126)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_80),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_42),
.B1(n_54),
.B2(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_31),
.B1(n_32),
.B2(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_9),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_40),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_32),
.B1(n_28),
.B2(n_22),
.Y(n_90)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_28),
.B1(n_18),
.B2(n_24),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_22),
.B1(n_33),
.B2(n_24),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_103),
.B1(n_118),
.B2(n_91),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_38),
.A2(n_15),
.B1(n_29),
.B2(n_33),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_43),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_106),
.B1(n_110),
.B2(n_8),
.Y(n_131)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_5),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_41),
.A2(n_23),
.B1(n_30),
.B2(n_35),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_29),
.B1(n_15),
.B2(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_74),
.B1(n_71),
.B2(n_108),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_57),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_116),
.B1(n_72),
.B2(n_91),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_48),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_37),
.B1(n_19),
.B2(n_4),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_139),
.B1(n_138),
.B2(n_123),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_37),
.B1(n_63),
.B2(n_67),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_128),
.B1(n_129),
.B2(n_155),
.Y(n_188)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_37),
.B1(n_68),
.B2(n_67),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_37),
.B1(n_68),
.B2(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_133),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_169),
.B1(n_134),
.B2(n_141),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_3),
.Y(n_133)
);

OR2x4_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_79),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_134),
.A2(n_154),
.B(n_130),
.C(n_163),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_158),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_72),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_143),
.Y(n_176)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_10),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_162),
.B1(n_164),
.B2(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_10),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_150),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_86),
.A2(n_12),
.B(n_0),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_161),
.B(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_76),
.B(n_0),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_153),
.B1(n_129),
.B2(n_128),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_93),
.B(n_113),
.CI(n_78),
.CON(n_154),
.SN(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_119),
.C(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_141),
.B1(n_161),
.B2(n_158),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_111),
.B(n_74),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_83),
.A2(n_111),
.B1(n_77),
.B2(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_83),
.A2(n_71),
.B1(n_92),
.B2(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_99),
.B(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_172),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_207),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_178),
.B(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_167),
.B1(n_126),
.B2(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_187),
.B1(n_137),
.B2(n_205),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_192),
.B1(n_165),
.B2(n_127),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_201),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_184),
.B1(n_186),
.B2(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_126),
.A2(n_132),
.B1(n_159),
.B2(n_124),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_136),
.B(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_176),
.Y(n_221)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_148),
.B1(n_133),
.B2(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_142),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_146),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_204),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_190),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_165),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_217),
.Y(n_262)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_219),
.C(n_220),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_127),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_241),
.C(n_216),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_137),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_192),
.B1(n_188),
.B2(n_185),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_220),
.B1(n_242),
.B2(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_186),
.B1(n_202),
.B2(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_221),
.B(n_224),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_175),
.B1(n_183),
.B2(n_195),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_209),
.C(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_234),
.C(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_209),
.C(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_206),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_211),
.B(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_179),
.B(n_181),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_240),
.B(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_180),
.B1(n_196),
.B2(n_175),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_208),
.B(n_171),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_247),
.A2(n_251),
.B1(n_255),
.B2(n_259),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_253),
.C(n_261),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_183),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_254),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_243),
.B1(n_223),
.B2(n_218),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_236),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_242),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_212),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_258),
.B(n_268),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_264),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_228),
.B(n_243),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_273),
.B(n_229),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_271),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_237),
.B(n_224),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_213),
.B(n_230),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_277),
.C(n_214),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_250),
.B1(n_276),
.B2(n_268),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_295),
.C(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_217),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_287),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_235),
.B1(n_221),
.B2(n_240),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_291),
.B1(n_269),
.B2(n_299),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_246),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_227),
.B1(n_247),
.B2(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_298),
.Y(n_310)
);

NAND5xp2_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_263),
.C(n_271),
.D(n_277),
.E(n_256),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_293),
.B(n_271),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_261),
.C(n_253),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_273),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_296),
.A2(n_303),
.B1(n_288),
.B2(n_285),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_251),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_302),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_248),
.B(n_250),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_307),
.C(n_311),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_265),
.C(n_252),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_288),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_265),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_303),
.B(n_296),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_269),
.C(n_258),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_320),
.C(n_286),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_260),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_318),
.B1(n_299),
.B2(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_297),
.C(n_284),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_278),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_294),
.B1(n_291),
.B2(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_327),
.B(n_332),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_315),
.B(n_297),
.C(n_296),
.D(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_328),
.B(n_338),
.Y(n_349)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_330),
.A2(n_331),
.B(n_334),
.Y(n_345)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.C(n_337),
.Y(n_340)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_294),
.B1(n_287),
.B2(n_285),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_316),
.B1(n_334),
.B2(n_331),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_301),
.C(n_300),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_303),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_320),
.C(n_307),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_344),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_326),
.C(n_304),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_309),
.Y(n_346)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_311),
.C(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_350),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_325),
.B(n_328),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_352),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_336),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_340),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_350),
.B(n_330),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_356),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_329),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_344),
.C(n_353),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_342),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_361),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_324),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_364),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_360),
.A2(n_351),
.B(n_357),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

NOR3xp33_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_362),
.C(n_348),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_366),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_345),
.A3(n_362),
.B1(n_347),
.B2(n_357),
.C1(n_349),
.C2(n_343),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);


endmodule