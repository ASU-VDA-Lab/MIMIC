module fake_netlist_1_7356_n_723 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_723);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_723;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_30), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_75), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_52), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_56), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_11), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_44), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_5), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_33), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_9), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_25), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_12), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_23), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_70), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_31), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_13), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_69), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_61), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_3), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_72), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_20), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_50), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_58), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_39), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_68), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_34), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_76), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_71), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_51), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_7), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_62), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_42), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_55), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_19), .Y(n_127) );
INVx6_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_80), .A2(n_28), .B(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_100), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_100), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_98), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_105), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_109), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_84), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_82), .B(n_29), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_88), .B(n_1), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_84), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
NOR2x1_ASAP7_75t_L g147 ( .A(n_112), .B(n_4), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_93), .B(n_6), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_82), .B(n_78), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
AOI22x1_ASAP7_75t_SL g157 ( .A1(n_97), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_107), .B(n_8), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_119), .B(n_9), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_127), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_102), .B(n_10), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_81), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_83), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_83), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_85), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_85), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_140), .A2(n_97), .B1(n_101), .B2(n_104), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_168), .B(n_126), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g175 ( .A(n_149), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_171), .B(n_99), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_129), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_170), .B(n_124), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_129), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_128), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_166), .B(n_108), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_170), .B(n_113), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_149), .B(n_123), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_171), .B(n_103), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_171), .Y(n_194) );
NAND2xp33_ASAP7_75t_R g195 ( .A(n_131), .B(n_116), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_171), .B(n_121), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_157), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_166), .B(n_117), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_168), .B(n_115), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_143), .A2(n_104), .B1(n_101), .B2(n_94), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_134), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_169), .B(n_114), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_152), .B(n_92), .C(n_90), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_169), .B(n_11), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_148), .Y(n_212) );
NAND2xp33_ASAP7_75t_SL g213 ( .A(n_170), .B(n_12), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_134), .B(n_15), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_167), .B(n_15), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_147), .B(n_18), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_150), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_165), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_170), .B(n_21), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_132), .B(n_22), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_167), .B(n_24), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_164), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_159), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_151), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_131), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_165), .B(n_26), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_131), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_151), .Y(n_235) );
AND3x1_ASAP7_75t_L g236 ( .A(n_140), .B(n_27), .C(n_32), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_159), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_175), .B(n_158), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_179), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_203), .B(n_165), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_223), .B(n_158), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g245 ( .A(n_210), .B(n_163), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_227), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_199), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_179), .A2(n_131), .B(n_142), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_203), .B(n_163), .Y(n_250) );
NOR2xp33_ASAP7_75t_R g251 ( .A(n_223), .B(n_153), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_187), .B(n_132), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_192), .A2(n_137), .B1(n_161), .B2(n_133), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_187), .B(n_133), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_230), .B(n_138), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_230), .B(n_138), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_199), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_230), .B(n_161), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_192), .B(n_134), .Y(n_259) );
BUFx12f_ASAP7_75t_SL g260 ( .A(n_220), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_176), .B(n_141), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_216), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_205), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_193), .B(n_141), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_206), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_179), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_155), .B(n_139), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_206), .B(n_159), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_183), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_232), .A2(n_139), .B(n_156), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_174), .B(n_144), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_178), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_204), .B(n_144), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_183), .A2(n_145), .B1(n_162), .B2(n_147), .Y(n_277) );
O2A1O1Ixp5_ASAP7_75t_L g278 ( .A1(n_233), .A2(n_156), .B(n_155), .C(n_146), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_208), .B(n_144), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_205), .A2(n_189), .B1(n_183), .B2(n_236), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_229), .B(n_146), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_207), .Y(n_282) );
BUFx6f_ASAP7_75t_SL g283 ( .A(n_220), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_229), .B(n_145), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_198), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_189), .A2(n_154), .B1(n_128), .B2(n_157), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_178), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_189), .B(n_225), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_236), .A2(n_154), .B1(n_128), .B2(n_151), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_197), .B(n_154), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_225), .B(n_151), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_237), .B(n_154), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_211), .A2(n_128), .B(n_37), .C(n_40), .Y(n_295) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_195), .B(n_36), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_194), .B(n_160), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_220), .B(n_160), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_237), .B(n_160), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_184), .B(n_160), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_194), .A2(n_160), .B1(n_43), .B2(n_45), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_184), .A2(n_217), .B(n_209), .C(n_173), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g305 ( .A(n_198), .B(n_41), .C(n_46), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_213), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_234), .A2(n_191), .B1(n_188), .B2(n_182), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_234), .A2(n_47), .B1(n_53), .B2(n_54), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_259), .B(n_191), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_244), .B(n_226), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_289), .A2(n_224), .B(n_231), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_243), .B(n_186), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_304), .A2(n_196), .B(n_231), .C(n_228), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_260), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_241), .B(n_60), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_250), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_263), .B(n_186), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_241), .B(n_186), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_283), .A2(n_186), .B1(n_228), .B2(n_222), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_285), .B(n_63), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_283), .A2(n_186), .B1(n_222), .B2(n_221), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_269), .B(n_65), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_280), .B(n_186), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_289), .A2(n_196), .B(n_221), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_262), .B(n_66), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_273), .A2(n_201), .B(n_172), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
BUFx2_ASAP7_75t_SL g330 ( .A(n_284), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_287), .B(n_201), .C(n_172), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_296), .B(n_235), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_262), .B(n_67), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_249), .A2(n_177), .B(n_180), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_296), .B(n_235), .Y(n_335) );
INVx5_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_272), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_270), .A2(n_177), .B(n_180), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_277), .B(n_181), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_293), .A2(n_181), .B(n_185), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_293), .A2(n_185), .B(n_190), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_248), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_299), .B(n_215), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_242), .A2(n_190), .B(n_202), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_300), .B(n_202), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_300), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_251), .B(n_215), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_252), .B(n_212), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_254), .A2(n_212), .B(n_214), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_256), .A2(n_214), .B(n_218), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_278), .A2(n_218), .B(n_215), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_258), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_276), .A2(n_215), .B(n_235), .C(n_279), .Y(n_353) );
AO32x1_ASAP7_75t_L g354 ( .A1(n_303), .A2(n_215), .A3(n_235), .B1(n_306), .B2(n_302), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_265), .A2(n_235), .B(n_274), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_253), .B(n_268), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_276), .A2(n_307), .B(n_271), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_279), .A2(n_245), .B(n_281), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_275), .B(n_288), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_248), .A2(n_257), .B(n_282), .C(n_298), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_266), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_291), .B(n_308), .C(n_295), .Y(n_362) );
NOR2x1_ASAP7_75t_SL g363 ( .A(n_336), .B(n_282), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_308), .B(n_301), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_353), .A2(n_297), .B(n_294), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_292), .B(n_290), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_257), .B(n_267), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_318), .B(n_264), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_311), .B(n_328), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_312), .B(n_286), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_333), .A2(n_292), .B(n_298), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_358), .A2(n_261), .B(n_290), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_362), .A2(n_261), .B(n_267), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_322), .A2(n_297), .B(n_240), .C(n_246), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_316), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_356), .B(n_251), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_356), .B(n_239), .Y(n_377) );
BUFx12f_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_357), .A2(n_239), .A3(n_240), .B(n_246), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_355), .A2(n_247), .B(n_305), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_314), .B(n_247), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_360), .B(n_339), .Y(n_382) );
AND2x6_ASAP7_75t_L g383 ( .A(n_317), .B(n_324), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_315), .A2(n_352), .B(n_359), .Y(n_384) );
OAI21xp33_ASAP7_75t_L g385 ( .A1(n_310), .A2(n_309), .B(n_348), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_331), .A2(n_342), .B(n_325), .C(n_361), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_330), .B(n_342), .Y(n_388) );
AO32x2_ASAP7_75t_L g389 ( .A1(n_354), .A2(n_323), .A3(n_346), .B1(n_336), .B2(n_343), .Y(n_389) );
CKINVDCx11_ASAP7_75t_R g390 ( .A(n_324), .Y(n_390) );
AOI21x1_ASAP7_75t_L g391 ( .A1(n_332), .A2(n_335), .B(n_341), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_344), .A2(n_326), .B(n_349), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_313), .A2(n_319), .B(n_347), .C(n_329), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_337), .A2(n_320), .B(n_350), .C(n_321), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_346), .B(n_345), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_346), .B(n_345), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_369), .A2(n_340), .B(n_354), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_381), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_354), .B1(n_383), .B2(n_390), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_382), .A2(n_373), .B(n_392), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_377), .B(n_376), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_391), .A2(n_382), .B(n_373), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_383), .A2(n_378), .B1(n_385), .B2(n_384), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_372), .B(n_366), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_371), .A2(n_374), .B(n_386), .Y(n_405) );
AO31x2_ASAP7_75t_L g406 ( .A1(n_379), .A2(n_365), .A3(n_389), .B(n_363), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_394), .A2(n_364), .B(n_380), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_364), .A2(n_384), .B(n_393), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_388), .B(n_396), .C(n_395), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_365), .A2(n_389), .B(n_379), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_396), .A2(n_389), .B(n_387), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_383), .A2(n_370), .B(n_375), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_383), .B(n_318), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_383), .B(n_363), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_367), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_383), .B(n_363), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_383), .B(n_363), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_384), .A2(n_280), .B(n_358), .Y(n_420) );
BUFx2_ASAP7_75t_SL g421 ( .A(n_383), .Y(n_421) );
OA21x2_ASAP7_75t_L g422 ( .A1(n_369), .A2(n_382), .B(n_373), .Y(n_422) );
BUFx2_ASAP7_75t_R g423 ( .A(n_376), .Y(n_423) );
OAI21x1_ASAP7_75t_L g424 ( .A1(n_369), .A2(n_392), .B(n_391), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_369), .A2(n_382), .B(n_373), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_398), .A2(n_401), .B1(n_403), .B2(n_421), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_407), .A2(n_397), .B(n_424), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_415), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_405), .A2(n_420), .B(n_407), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_415), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_411), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_417), .A2(n_397), .B(n_424), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_415), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_417), .Y(n_436) );
AOI21x1_ASAP7_75t_L g437 ( .A1(n_408), .A2(n_404), .B(n_400), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_408), .A2(n_410), .B(n_404), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_403), .B(n_400), .Y(n_439) );
OAI21x1_ASAP7_75t_L g440 ( .A1(n_402), .A2(n_400), .B(n_425), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_422), .B(n_425), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_400), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_422), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_415), .Y(n_446) );
AOI21x1_ASAP7_75t_L g447 ( .A1(n_402), .A2(n_425), .B(n_422), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_414), .B(n_423), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_422), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_412), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_412), .A2(n_399), .B(n_413), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_418), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_413), .A2(n_409), .B(n_410), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_421), .A2(n_416), .B1(n_418), .B2(n_419), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_425), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_406), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_410), .A2(n_419), .B(n_416), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_429), .B(n_419), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_429), .B(n_432), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_436), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_432), .B(n_434), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_441), .B(n_462), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_426), .A2(n_448), .B1(n_455), .B2(n_439), .C(n_435), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_436), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_442), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_441), .B(n_462), .Y(n_473) );
NAND2xp33_ASAP7_75t_R g474 ( .A(n_428), .B(n_446), .Y(n_474) );
OR2x2_ASAP7_75t_SL g475 ( .A(n_459), .B(n_451), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_441), .B(n_462), .Y(n_476) );
INVx8_ASAP7_75t_L g477 ( .A(n_428), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_428), .B(n_460), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_459), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_442), .B(n_431), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_444), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_428), .B(n_452), .Y(n_483) );
OR2x6_ASAP7_75t_L g484 ( .A(n_431), .B(n_435), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_444), .Y(n_486) );
NAND3xp33_ASAP7_75t_SL g487 ( .A(n_448), .B(n_455), .C(n_426), .Y(n_487) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_433), .A2(n_437), .B(n_447), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_443), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_431), .B(n_446), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_445), .B(n_457), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_457), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_428), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_453), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_446), .B(n_452), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_458), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_446), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_458), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_449), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_446), .B(n_460), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_439), .B(n_461), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_452), .B(n_460), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_433), .A2(n_440), .B(n_437), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_452), .Y(n_511) );
OR2x6_ASAP7_75t_L g512 ( .A(n_452), .B(n_460), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g513 ( .A1(n_460), .A2(n_451), .B1(n_456), .B2(n_454), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_469), .B(n_461), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_498), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_466), .B(n_461), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_469), .B(n_461), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_473), .B(n_461), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_466), .B(n_451), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_482), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_468), .B(n_451), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_482), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_486), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_473), .B(n_451), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_486), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_476), .B(n_451), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_480), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_495), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_476), .B(n_454), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_492), .B(n_454), .Y(n_531) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_490), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_492), .B(n_454), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_493), .B(n_454), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_496), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_478), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_493), .B(n_454), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_468), .B(n_430), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_496), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_484), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_464), .B(n_430), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_464), .B(n_430), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_463), .B(n_430), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_499), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_463), .B(n_430), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_472), .B(n_440), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_472), .B(n_440), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_438), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_504), .B(n_438), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_501), .B(n_438), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_481), .B(n_438), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_485), .Y(n_555) );
AND2x2_ASAP7_75t_SL g556 ( .A(n_478), .B(n_450), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_487), .B(n_450), .Y(n_557) );
INVx5_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_481), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_503), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_503), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_505), .B(n_438), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_509), .Y(n_564) );
INVxp67_ASAP7_75t_SL g565 ( .A(n_509), .Y(n_565) );
INVx4_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_427), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_520), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_522), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_559), .B(n_506), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_561), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_524), .B(n_510), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_522), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_568), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_524), .B(n_489), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_523), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_518), .B(n_475), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_527), .B(n_502), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_523), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_528), .B(n_502), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_558), .B(n_478), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_527), .B(n_508), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_514), .B(n_465), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_525), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_465), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_541), .B(n_566), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_517), .B(n_465), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_488), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_518), .B(n_475), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_516), .B(n_545), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_525), .Y(n_594) );
INVxp33_ASAP7_75t_L g595 ( .A(n_541), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_535), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_543), .B(n_478), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_565), .B(n_491), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_541), .B(n_483), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_526), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_551), .B(n_488), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_526), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_537), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_543), .B(n_513), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_558), .B(n_497), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_551), .B(n_488), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_552), .B(n_467), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_550), .B(n_479), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_547), .B(n_507), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_519), .B(n_471), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_552), .B(n_467), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_541), .B(n_484), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_515), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_544), .B(n_471), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_529), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_529), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_479), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_567), .B(n_500), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_536), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_530), .B(n_479), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_576), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_585), .B(n_538), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_591), .B(n_557), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_593), .B(n_554), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_613), .B(n_566), .Y(n_626) );
NAND2xp33_ASAP7_75t_L g627 ( .A(n_595), .B(n_558), .Y(n_627) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_602), .B(n_558), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_572), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_593), .B(n_554), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_591), .B(n_538), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_569), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_605), .B(n_470), .C(n_555), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_585), .B(n_534), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_618), .B(n_534), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_610), .B(n_533), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_589), .A2(n_566), .B1(n_556), .B2(n_558), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_610), .B(n_521), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_618), .B(n_533), .Y(n_639) );
AO221x1_ASAP7_75t_L g640 ( .A1(n_604), .A2(n_474), .B1(n_558), .B2(n_566), .C(n_562), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_601), .B(n_531), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_583), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_571), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_575), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_601), .B(n_531), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_607), .B(n_550), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_621), .B(n_556), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_578), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_607), .B(n_586), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_577), .B(n_560), .Y(n_652) );
OAI21xp33_ASAP7_75t_SL g653 ( .A1(n_573), .A2(n_556), .B(n_484), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_574), .B(n_563), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_577), .B(n_560), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_587), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_581), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_574), .B(n_563), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_635), .B(n_621), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_653), .A2(n_595), .B(n_584), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_624), .A2(n_579), .B(n_592), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_652), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_625), .B(n_579), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_633), .B(n_592), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g666 ( .A1(n_629), .A2(n_597), .A3(n_609), .B1(n_615), .B2(n_598), .C1(n_611), .C2(n_619), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_642), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_637), .A2(n_477), .B(n_619), .C(n_615), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_633), .A2(n_589), .B1(n_599), .B2(n_553), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_638), .B(n_586), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_655), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_638), .A2(n_580), .B(n_589), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_632), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_627), .A2(n_584), .B(n_599), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_643), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_622), .A2(n_599), .B1(n_553), .B2(n_479), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_644), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_623), .B(n_590), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_645), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_649), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_630), .B(n_611), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_648), .A2(n_608), .B1(n_612), .B2(n_588), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_658), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_669), .A2(n_637), .B(n_626), .C(n_647), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_665), .A2(n_640), .B1(n_623), .B2(n_627), .Y(n_685) );
NOR4xp25_ASAP7_75t_L g686 ( .A(n_666), .B(n_657), .C(n_656), .D(n_651), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_674), .A2(n_661), .B(n_668), .Y(n_687) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_662), .A2(n_631), .B1(n_646), .B2(n_641), .C(n_634), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_669), .A2(n_628), .B1(n_636), .B2(n_650), .Y(n_689) );
OA22x2_ASAP7_75t_L g690 ( .A1(n_672), .A2(n_639), .B1(n_659), .B2(n_654), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_667), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_667), .B(n_658), .C(n_539), .Y(n_692) );
OAI22xp33_ASAP7_75t_SL g693 ( .A1(n_664), .A2(n_628), .B1(n_606), .B2(n_537), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_676), .B(n_537), .C(n_483), .D(n_548), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_681), .B(n_659), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_671), .A2(n_654), .B1(n_620), .B2(n_617), .C(n_616), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_663), .B(n_580), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g698 ( .A1(n_686), .A2(n_676), .B1(n_682), .B2(n_680), .C(n_679), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_684), .B(n_677), .C(n_675), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_687), .A2(n_670), .B(n_673), .C(n_678), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_689), .B(n_683), .C(n_600), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_691), .A2(n_683), .B(n_606), .C(n_660), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_688), .A2(n_603), .B1(n_588), .B2(n_590), .C(n_612), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_696), .B(n_608), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_694), .A2(n_693), .B1(n_692), .B2(n_685), .C(n_697), .Y(n_705) );
NOR3xp33_ASAP7_75t_SL g706 ( .A(n_700), .B(n_690), .C(n_494), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_705), .A2(n_695), .B(n_477), .C(n_546), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_704), .B(n_549), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_701), .B(n_549), .C(n_546), .Y(n_709) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_699), .B(n_512), .Y(n_710) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_710), .B(n_703), .C(n_698), .D(n_702), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_708), .B(n_540), .Y(n_712) );
NOR3x1_ASAP7_75t_L g713 ( .A(n_707), .B(n_540), .C(n_542), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_706), .B1(n_709), .B2(n_542), .C(n_536), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_713), .B(n_512), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_716), .Y(n_717) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_717), .Y(n_718) );
OAI22x1_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_711), .B1(n_714), .B2(n_483), .Y(n_719) );
AOI221x1_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_564), .B1(n_562), .B2(n_614), .C(n_596), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_720), .B(n_614), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_477), .B1(n_483), .B2(n_512), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_512), .B1(n_477), .B2(n_564), .Y(n_723) );
endmodule