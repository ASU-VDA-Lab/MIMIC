module real_jpeg_16469_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_286;
wire n_215;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_1),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_1),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_1),
.B(n_369),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_3),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_3),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_3),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_4),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_4),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_4),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_4),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_4),
.B(n_476),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_4),
.B(n_506),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_6),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_6),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_7),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

AND2x4_ASAP7_75t_SL g221 ( 
.A(n_7),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_7),
.B(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_8),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx4f_ASAP7_75t_L g535 ( 
.A(n_8),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_9),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

AOI22x1_ASAP7_75t_SL g299 ( 
.A1(n_9),
.A2(n_17),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_9),
.B(n_93),
.Y(n_373)
);

AOI31xp33_ASAP7_75t_L g409 ( 
.A1(n_9),
.A2(n_299),
.A3(n_410),
.B(n_415),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_9),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_9),
.B(n_488),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_9),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_9),
.B(n_171),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_10),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_144),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_10),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_10),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_10),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_10),
.B(n_413),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_11),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_11),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_11),
.B(n_566),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_12),
.B(n_99),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_12),
.B(n_247),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_12),
.B(n_267),
.Y(n_266)
);

AND2x4_ASAP7_75t_SL g324 ( 
.A(n_12),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_12),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_12),
.B(n_422),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_12),
.B(n_370),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_14),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_14),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_14),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_14),
.B(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_14),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_14),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_14),
.B(n_533),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_15),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_15),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_17),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_17),
.B(n_258),
.Y(n_257)
);

NAND2x1_ASAP7_75t_L g261 ( 
.A(n_17),
.B(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_17),
.Y(n_411)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_18),
.Y(n_567)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_561),
.B(n_568),
.C(n_570),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_116),
.B(n_560),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_70),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_27),
.B(n_70),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_54),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_29),
.B(n_41),
.C(n_54),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_37),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_30),
.A2(n_34),
.B1(n_48),
.B2(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g563 ( 
.A(n_30),
.B(n_43),
.C(n_50),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_33),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g447 ( 
.A(n_33),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_64),
.C(n_66),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_34),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_43),
.A2(n_49),
.B1(n_565),
.B2(n_568),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_47),
.B(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_56),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_59),
.B(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2x1_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_66),
.A2(n_67),
.B1(n_107),
.B2(n_128),
.Y(n_184)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_103),
.C(n_107),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_112),
.C(n_113),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_102),
.C(n_110),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_72),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_78),
.C(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_77),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_81),
.Y(n_335)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_81),
.Y(n_418)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.C(n_96),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_166)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_100),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_110),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_103),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_124),
.C(n_129),
.Y(n_185)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_108),
.Y(n_472)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_109),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_289),
.B(n_555),
.Y(n_116)
);

NOR3x1_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_192),
.C(n_283),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_118),
.A2(n_556),
.B(n_559),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_R g118 ( 
.A(n_119),
.B(n_190),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_119),
.B(n_190),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_182),
.C(n_187),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_120),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_164),
.C(n_167),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_122),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.C(n_148),
.Y(n_122)
);

XNOR2x2_ASAP7_75t_SL g231 ( 
.A(n_123),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_129),
.A2(n_130),
.B1(n_170),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_170),
.C(n_173),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_132),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_134),
.B(n_148),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_143),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_135),
.B(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_137),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_138),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_154),
.C(n_160),
.Y(n_186)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_152),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_165),
.B(n_167),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.C(n_178),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_169),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_217),
.C(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_170),
.Y(n_230)
);

AOI22x1_ASAP7_75t_L g236 ( 
.A1(n_170),
.A2(n_221),
.B1(n_230),
.B2(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_173),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_173),
.A2(n_227),
.B1(n_312),
.B2(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_175),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_177),
.B(n_254),
.C(n_257),
.Y(n_253)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_178),
.A2(n_209),
.B1(n_212),
.B2(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_182),
.A2(n_187),
.B1(n_188),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_182),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_183),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_185),
.B(n_186),
.Y(n_278)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_273),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_193),
.B(n_273),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_231),
.C(n_233),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_195),
.B(n_231),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_213),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_197),
.B(n_200),
.C(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_209),
.C(n_212),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_208),
.Y(n_251)
);

XOR2x1_ASAP7_75t_SL g250 ( 
.A(n_204),
.B(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_211),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_226),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_214),
.B(n_216),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

BUFx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_225),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_226),
.B(n_344),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_307),
.C(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_233),
.B(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_252),
.C(n_269),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_234),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_250),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_235),
.B(n_238),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_245),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_239),
.A2(n_245),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_239),
.Y(n_386)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_242),
.B(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_245),
.B(n_444),
.C(n_448),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_245),
.A2(n_385),
.B1(n_444),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_246),
.Y(n_385)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_250),
.B(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_252),
.B(n_270),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_261),
.C(n_265),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_253),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_257),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_255),
.Y(n_506)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_256),
.Y(n_371)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_260),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_260),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_261),
.A2(n_265),
.B1(n_266),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_265),
.A2(n_266),
.B1(n_425),
.B2(n_426),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_266),
.B(n_420),
.C(n_425),
.Y(n_419)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_277),
.C(n_282),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_284),
.A2(n_557),
.B(n_558),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_285),
.B(n_288),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_394),
.B(n_552),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_387),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_347),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_292),
.B(n_347),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_340),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_293),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_315),
.C(n_336),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.C(n_306),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_296),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_298),
.A2(n_299),
.B1(n_306),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_306),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_309),
.Y(n_486)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_314),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_316),
.A2(n_336),
.B1(n_337),
.B2(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_316),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_327),
.C(n_333),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.C(n_324),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_318),
.A2(n_324),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_322),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_324),
.B(n_499),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_326),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_333),
.Y(n_382)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_331),
.Y(n_490)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.C(n_356),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_349),
.A2(n_350),
.B1(n_354),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_381),
.C(n_383),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.C(n_372),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g453 ( 
.A(n_360),
.B(n_454),
.Y(n_453)
);

XNOR2x1_ASAP7_75t_L g454 ( 
.A(n_363),
.B(n_372),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_364),
.B(n_368),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.C(n_379),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_373),
.A2(n_374),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_373),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_374),
.A2(n_441),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_374),
.B(n_518),
.C(n_522),
.Y(n_542)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_379),
.B(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_383),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_387),
.A2(n_553),
.B(n_554),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_388),
.B(n_390),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.C(n_393),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_457),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.C(n_432),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_397),
.B(n_401),
.Y(n_551)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_428),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_404),
.B(n_429),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_409),
.C(n_419),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_409),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_485),
.C(n_487),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_420),
.B(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_424),
.Y(n_470)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_421),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_421),
.A2(n_515),
.B1(n_516),
.B2(n_530),
.Y(n_529)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_455),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_455),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.C(n_453),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_434),
.B(n_549),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_437),
.B(n_453),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.C(n_451),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_480),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_452),
.Y(n_480)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

XOR2x1_ASAP7_75t_L g492 ( 
.A(n_448),
.B(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.C(n_551),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_546),
.B(n_550),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_495),
.B(n_545),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_481),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_481),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_478),
.B2(n_479),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_465),
.B(n_469),
.C(n_478),
.Y(n_547)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.C(n_473),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_471),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

AO22x1_ASAP7_75t_SL g507 ( 
.A1(n_474),
.A2(n_475),
.B1(n_477),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_477),
.Y(n_508)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_491),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_484),
.B(n_492),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_487),
.Y(n_499)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

OAI21x1_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_511),
.B(n_544),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_509),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_509),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.C(n_507),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_498),
.B(n_540),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_500),
.A2(n_501),
.B1(n_507),
.B2(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_502),
.B(n_505),
.Y(n_519)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_532),
.Y(n_531)
);

AOI21x1_ASAP7_75t_SL g511 ( 
.A1(n_512),
.A2(n_538),
.B(n_543),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_513),
.A2(n_525),
.B(n_537),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_517),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_517),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_518),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_531),
.B(n_536),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_529),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_539),
.B(n_542),
.Y(n_538)
);

NOR2x1_ASAP7_75t_SL g543 ( 
.A(n_539),
.B(n_542),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_548),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_569),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_569),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_565),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_571),
.Y(n_570)
);


endmodule