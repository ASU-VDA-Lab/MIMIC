module real_jpeg_14758_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_316, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_316;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_3),
.A2(n_46),
.B1(n_49),
.B2(n_158),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_103),
.B1(n_104),
.B2(n_158),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_3),
.A2(n_152),
.B1(n_153),
.B2(n_158),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_5),
.A2(n_48),
.B1(n_103),
.B2(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_48),
.B1(n_152),
.B2(n_153),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_6),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_40),
.B1(n_46),
.B2(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_7),
.A2(n_40),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_40),
.B1(n_152),
.B2(n_153),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_9),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_10),
.B(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_30),
.C(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_33),
.B1(n_46),
.B2(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_10),
.B(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_33),
.B1(n_103),
.B2(n_104),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_60),
.B(n_104),
.C(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_10),
.A2(n_33),
.B1(n_152),
.B2(n_153),
.Y(n_170)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_251),
.C(n_307),
.Y(n_12)
);

OA21x2_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_306),
.B(n_311),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_298),
.B(n_305),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_260),
.B(n_295),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_241),
.B(n_259),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_220),
.B(n_240),
.Y(n_17)
);

AOI321xp33_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_181),
.A3(n_213),
.B1(n_218),
.B2(n_219),
.C(n_316),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_142),
.B(n_180),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_119),
.B(n_141),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_96),
.B(n_118),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_74),
.B(n_95),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_65),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_65),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_24)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_26),
.B(n_92),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_38),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_28),
.A2(n_35),
.B(n_38),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_78),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_49),
.B(n_61),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_33),
.B(n_104),
.C(n_132),
.Y(n_151)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_35),
.A2(n_92),
.B(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_37),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_38),
.B(n_85),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_38),
.A2(n_157),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_44),
.B(n_71),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_44),
.A2(n_178),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_50),
.B(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_53),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_54),
.Y(n_178)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_62),
.C(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_58),
.B(n_109),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_58),
.A2(n_106),
.B(n_109),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_58),
.A2(n_174),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_59),
.B(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_61),
.B1(n_103),
.B2(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_73),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_88),
.B(n_94),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_82),
.B(n_87),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_86),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_110),
.C(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_104),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_107),
.B(n_136),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_107),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_179),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_111),
.B(n_123),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_113),
.A2(n_114),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_113),
.A2(n_114),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_114),
.B(n_237),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_114),
.A2(n_248),
.B(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_140),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_140),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_127),
.B1(n_128),
.B2(n_139),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_125),
.C(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_128),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.CI(n_134),
.CON(n_128),
.SN(n_128)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.C(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_131),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_133),
.B1(n_152),
.B2(n_153),
.Y(n_169)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_135),
.B(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_135),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_160),
.B2(n_161),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_147),
.B(n_148),
.C(n_160),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_156),
.B2(n_159),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_171),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_173),
.C(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_165),
.B(n_168),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_167),
.A2(n_170),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_167),
.A2(n_185),
.B(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_174),
.B(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_176),
.A2(n_177),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_176),
.A2(n_177),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_177),
.B(n_268),
.C(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_177),
.B(n_292),
.C(n_294),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_208),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_193),
.C(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_191),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_188),
.CI(n_191),
.CON(n_210),
.SN(n_210)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_185),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_230),
.Y(n_229)
);

NAND2x1_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_189),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_201),
.C(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_200),
.A2(n_252),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_200),
.B(n_230),
.Y(n_308)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_201),
.A2(n_203),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_201),
.B(n_303),
.C(n_304),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_210),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_239),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_235),
.B2(n_236),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_236),
.C(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_228),
.C(n_233),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_243),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.C(n_254),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_253),
.B2(n_254),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B(n_258),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_266),
.B1(n_267),
.B2(n_277),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_264),
.C(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_263),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_269),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_281),
.C(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_273),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_310),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);


endmodule