module fake_jpeg_1069_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_12),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_44),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_62),
.B(n_58),
.C(n_61),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_88),
.B(n_48),
.C(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_63),
.B1(n_62),
.B2(n_40),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_53),
.B1(n_55),
.B2(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_40),
.C(n_46),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_49),
.CI(n_50),
.CON(n_105),
.SN(n_105)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_56),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_47),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_22),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_56),
.B(n_70),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_49),
.B(n_2),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_100),
.B(n_4),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_52),
.B1(n_63),
.B2(n_55),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_41),
.B(n_42),
.C(n_50),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_81),
.Y(n_107)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_119),
.C(n_121),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_8),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_118),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_10),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_116),
.B1(n_99),
.B2(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_128),
.B1(n_134),
.B2(n_135),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_105),
.B1(n_23),
.B2(n_26),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_136),
.B(n_139),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_114),
.C(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_108),
.C(n_114),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_147),
.C(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_138),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_137),
.Y(n_148)
);

AOI321xp33_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_143),
.A3(n_145),
.B1(n_146),
.B2(n_144),
.C(n_14),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_133),
.B1(n_128),
.B2(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_151),
.B(n_28),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_19),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

OAI321xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_153),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_10),
.C(n_11),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_13),
.B(n_29),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_31),
.B(n_32),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_34),
.Y(n_163)
);


endmodule