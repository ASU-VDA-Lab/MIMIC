module fake_jpeg_2151_n_511 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_511);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_511;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_120)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_76),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_39),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_92),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_1),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_93),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_98),
.B(n_99),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_96),
.B(n_97),
.Y(n_162)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_23),
.B1(n_49),
.B2(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_43),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_18),
.B1(n_45),
.B2(n_27),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_104),
.B(n_111),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_107),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_101),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_18),
.B1(n_41),
.B2(n_32),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_20),
.B1(n_19),
.B2(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_114),
.A2(n_131),
.B1(n_132),
.B2(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_18),
.B1(n_41),
.B2(n_20),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_116),
.A2(n_120),
.B1(n_156),
.B2(n_2),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_47),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_54),
.A2(n_42),
.B1(n_31),
.B2(n_28),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_137),
.B1(n_156),
.B2(n_116),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_43),
.B1(n_49),
.B2(n_46),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_44),
.B1(n_32),
.B2(n_31),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_58),
.B(n_44),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_142),
.B(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_71),
.B(n_30),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_157),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_68),
.A2(n_30),
.B1(n_50),
.B2(n_26),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_50),
.B1(n_26),
.B2(n_25),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_1),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_60),
.A2(n_50),
.B1(n_26),
.B2(n_48),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_161),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_53),
.B(n_1),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_84),
.A2(n_74),
.B1(n_88),
.B2(n_66),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_166),
.B(n_174),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_100),
.C(n_52),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_170),
.C(n_206),
.Y(n_228)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_168),
.Y(n_256)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_108),
.B(n_101),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_90),
.B1(n_86),
.B2(n_83),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_172),
.A2(n_179),
.B1(n_201),
.B2(n_126),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_91),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_91),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_176),
.A2(n_216),
.B1(n_159),
.B2(n_123),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_192),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_82),
.B1(n_69),
.B2(n_65),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_100),
.C(n_73),
.Y(n_184)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_185),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_73),
.B(n_66),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_111),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_63),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

AND2x4_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_2),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_4),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_4),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_117),
.B(n_4),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_200),
.B(n_208),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_137),
.A2(n_113),
.B1(n_109),
.B2(n_130),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_140),
.B(n_5),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_141),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_6),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_6),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_16),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_209),
.C(n_9),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_106),
.B(n_109),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_105),
.B(n_16),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_106),
.B(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_211),
.B(n_9),
.Y(n_252)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_123),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_144),
.B(n_7),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_113),
.B(n_9),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_224),
.B(n_230),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_159),
.B1(n_150),
.B2(n_149),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_227),
.B1(n_239),
.B2(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_177),
.A2(n_103),
.B1(n_150),
.B2(n_149),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_141),
.B(n_154),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_229),
.A2(n_249),
.B(n_264),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_166),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_167),
.B1(n_207),
.B2(n_206),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_177),
.A2(n_103),
.B1(n_155),
.B2(n_135),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_112),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_246),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_193),
.A2(n_112),
.B(n_129),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_171),
.B(n_155),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_135),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_252),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_170),
.A2(n_126),
.B1(n_10),
.B2(n_12),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_194),
.B1(n_210),
.B2(n_213),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_259),
.B(n_261),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_199),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_12),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_163),
.A2(n_14),
.B(n_15),
.C(n_176),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_189),
.B(n_163),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_265),
.B(n_173),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_174),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_267),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_170),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_274),
.C(n_278),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_182),
.B1(n_190),
.B2(n_204),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_269),
.A2(n_304),
.B(n_245),
.Y(n_336)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_271),
.A2(n_273),
.B1(n_294),
.B2(n_229),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_272),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_190),
.B1(n_219),
.B2(n_218),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_164),
.C(n_183),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_220),
.B(n_212),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_205),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_286),
.C(n_259),
.Y(n_341)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_241),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_300),
.Y(n_317)
);

NOR2x1p5_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_188),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_224),
.Y(n_310)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_243),
.C(n_221),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_188),
.B1(n_190),
.B2(n_206),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_305),
.B1(n_230),
.B2(n_225),
.Y(n_328)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_293),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_233),
.A2(n_207),
.B1(n_209),
.B2(n_195),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_296),
.B(n_297),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_214),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_225),
.B(n_173),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_185),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_230),
.B1(n_248),
.B2(n_237),
.Y(n_308)
);

AO22x1_ASAP7_75t_L g303 ( 
.A1(n_226),
.A2(n_209),
.B1(n_168),
.B2(n_198),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_253),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_202),
.B1(n_181),
.B2(n_165),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_245),
.Y(n_306)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_310),
.A2(n_314),
.B(n_321),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_323),
.B1(n_271),
.B2(n_275),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_295),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_313),
.B(n_322),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_304),
.B(n_276),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_249),
.B(n_244),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_264),
.B1(n_225),
.B2(n_250),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_234),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_337),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_222),
.C(n_234),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_310),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_278),
.B(n_251),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_327),
.B(n_335),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_328),
.A2(n_334),
.B1(n_343),
.B2(n_282),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_330),
.A2(n_294),
.B1(n_301),
.B2(n_281),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_269),
.A2(n_222),
.B1(n_262),
.B2(n_261),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_284),
.B(n_242),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_291),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_283),
.A2(n_257),
.B(n_240),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_318),
.C(n_274),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_292),
.A2(n_263),
.B1(n_239),
.B2(n_252),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_344),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_358),
.C(n_373),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_223),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_347),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_283),
.B1(n_290),
.B2(n_288),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_290),
.B1(n_339),
.B2(n_322),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_286),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_371),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_312),
.A2(n_323),
.B1(n_330),
.B2(n_277),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_342),
.B1(n_338),
.B2(n_329),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_311),
.B(n_223),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_354),
.B(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_268),
.C(n_299),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_242),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_335),
.B(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_303),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_320),
.Y(n_380)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_257),
.Y(n_365)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_SL g366 ( 
.A(n_340),
.B(n_273),
.C(n_282),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_366),
.A2(n_227),
.B(n_303),
.Y(n_401)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_247),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_369),
.A2(n_372),
.B(n_377),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_370),
.A2(n_376),
.B1(n_330),
.B2(n_337),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_327),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_247),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_280),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_325),
.C(n_321),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_287),
.C(n_241),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_275),
.B1(n_305),
.B2(n_285),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_237),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_351),
.A2(n_336),
.B(n_350),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_378),
.A2(n_405),
.B(n_386),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_384),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_317),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_342),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_397),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_388),
.B1(n_393),
.B2(n_394),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_389),
.A2(n_402),
.B1(n_357),
.B2(n_367),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_370),
.A2(n_338),
.B1(n_329),
.B2(n_324),
.Y(n_393)
);

OAI22x1_ASAP7_75t_L g394 ( 
.A1(n_346),
.A2(n_324),
.B1(n_333),
.B2(n_332),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_333),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_376),
.A2(n_332),
.B1(n_319),
.B2(n_293),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_331),
.B1(n_319),
.B2(n_272),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_331),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_362),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_367),
.B1(n_356),
.B2(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_403),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_374),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_406),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_309),
.B(n_331),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_366),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_356),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_375),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_319),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_362),
.Y(n_416)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_383),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_417),
.A2(n_424),
.B1(n_427),
.B2(n_429),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_402),
.A2(n_346),
.B1(n_349),
.B2(n_375),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_419),
.A2(n_426),
.B1(n_394),
.B2(n_382),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_379),
.B(n_349),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_420),
.B(n_431),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_422),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_368),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_355),
.C(n_270),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_395),
.C(n_397),
.Y(n_436)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_428),
.Y(n_445)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_240),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_430),
.A2(n_378),
.B(n_386),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_405),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_L g455 ( 
.A1(n_432),
.A2(n_430),
.B(n_407),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_434),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_385),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_440),
.C(n_418),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_439),
.C(n_450),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_381),
.C(n_384),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_404),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_399),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_447),
.C(n_451),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_409),
.B(n_380),
.Y(n_447)
);

BUFx12_ASAP7_75t_L g449 ( 
.A(n_428),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_419),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_406),
.C(n_403),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_458),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_455),
.A2(n_346),
.B(n_256),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_467),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_437),
.A2(n_407),
.B1(n_427),
.B2(n_408),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_424),
.B1(n_435),
.B2(n_449),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_410),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_439),
.B(n_422),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_459),
.B(n_466),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_432),
.A2(n_446),
.B(n_450),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_445),
.B(n_443),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_416),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_255),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_412),
.B(n_421),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_462),
.A2(n_443),
.B(n_445),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_441),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_465),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_418),
.C(n_412),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_426),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_463),
.A2(n_434),
.B(n_442),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_468),
.A2(n_180),
.B(n_14),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_472),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_464),
.B(n_438),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_471),
.B(n_474),
.Y(n_490)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_449),
.C(n_346),
.Y(n_474)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_478),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_255),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_479),
.B(n_197),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_467),
.C(n_463),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_484),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_461),
.B1(n_462),
.B2(n_455),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_456),
.C(n_256),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_491),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_169),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_475),
.B(n_478),
.Y(n_493)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_493),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_480),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_494),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_477),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_498),
.B(n_489),
.Y(n_502)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_469),
.Y(n_498)
);

NAND2x1_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_489),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_500),
.A2(n_494),
.B(n_495),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_502),
.B(n_482),
.Y(n_506)
);

AO21x1_ASAP7_75t_L g507 ( 
.A1(n_504),
.A2(n_500),
.B(n_501),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_503),
.A2(n_496),
.B1(n_486),
.B2(n_487),
.Y(n_505)
);

AOI221xp5_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_506),
.B1(n_487),
.B2(n_180),
.C(n_15),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_508),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_509),
.B(n_180),
.CI(n_15),
.CON(n_510),
.SN(n_510)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_15),
.B(n_236),
.Y(n_511)
);


endmodule