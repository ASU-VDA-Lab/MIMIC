module fake_jpeg_16109_n_237 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_18),
.B1(n_28),
.B2(n_24),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_58),
.B1(n_20),
.B2(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_17),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_52),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_84),
.B(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_25),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_63),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_68),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_69),
.B1(n_73),
.B2(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_27),
.B1(n_21),
.B2(n_23),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_85),
.Y(n_119)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_58),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_32),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_88),
.C(n_67),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_26),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_32),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_33),
.B(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_52),
.B(n_33),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_31),
.B1(n_30),
.B2(n_3),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_33),
.B1(n_26),
.B2(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_80),
.B1(n_92),
.B2(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_109),
.B1(n_61),
.B2(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_120),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_86),
.CI(n_84),
.CON(n_134),
.SN(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_6),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_124),
.B1(n_108),
.B2(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_126),
.Y(n_152)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_66),
.B(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_77),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_141),
.B1(n_143),
.B2(n_101),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_84),
.B(n_86),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_140),
.B(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_65),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_82),
.B1(n_80),
.B2(n_90),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_96),
.B1(n_113),
.B2(n_95),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_110),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_89),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_75),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_74),
.B1(n_66),
.B2(n_71),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_75),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_74),
.B1(n_87),
.B2(n_9),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_116),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_153),
.C(n_166),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_128),
.B1(n_132),
.B2(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_155),
.B1(n_156),
.B2(n_164),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_115),
.B1(n_99),
.B2(n_109),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_112),
.B1(n_102),
.B2(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_95),
.B(n_107),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_163),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_107),
.B(n_33),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_161),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_26),
.B(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_26),
.B(n_10),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_150),
.B1(n_164),
.B2(n_166),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_173),
.B1(n_176),
.B2(n_181),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_133),
.A3(n_134),
.B1(n_128),
.B2(n_135),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI21x1_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_134),
.B(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_141),
.B1(n_127),
.B2(n_122),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_151),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_144),
.B1(n_137),
.B2(n_125),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_151),
.B1(n_161),
.B2(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_146),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.C(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_153),
.C(n_174),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_160),
.B(n_154),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_183),
.B(n_170),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_165),
.B1(n_152),
.B2(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_179),
.B1(n_171),
.B2(n_176),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_129),
.B1(n_116),
.B2(n_11),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_205),
.B(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_193),
.B(n_194),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_211),
.B(n_198),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_192),
.B1(n_184),
.B2(n_196),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_184),
.B1(n_185),
.B2(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_222),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_224),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_211),
.B(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_213),
.C(n_199),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_227),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_212),
.B1(n_204),
.B2(n_220),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_231),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_218),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_226),
.B(n_129),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_231),
.B(n_10),
.C(n_11),
.D(n_13),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_235),
.C(n_15),
.Y(n_236)
);

AOI321xp33_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_15),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_7),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_7),
.Y(n_237)
);


endmodule