module fake_netlist_6_1797_n_197 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_197);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_197;

wire n_52;
wire n_91;
wire n_119;
wire n_146;
wire n_163;
wire n_46;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_78;
wire n_66;
wire n_84;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_R g56 ( 
.A(n_49),
.B(n_19),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_R g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_1),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_42),
.B1(n_55),
.B2(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_62),
.B1(n_75),
.B2(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_72),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_33),
.B(n_74),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_56),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_41),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_71),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_63),
.B(n_70),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

OAI21x1_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_104),
.B(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_92),
.B(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_94),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_100),
.B1(n_106),
.B2(n_98),
.Y(n_117)
);

NOR2x1_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_102),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_106),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_106),
.C(n_113),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_119),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_114),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_119),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_118),
.B(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_87),
.B1(n_130),
.B2(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_66),
.B1(n_135),
.B2(n_87),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_132),
.B1(n_136),
.B2(n_126),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_132),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_134),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_139),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_139),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_136),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_47),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_136),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_144),
.B(n_150),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_53),
.B1(n_47),
.B2(n_46),
.C(n_43),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_53),
.B1(n_46),
.B2(n_43),
.C(n_39),
.Y(n_166)
);

NAND4xp75_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_148),
.C(n_39),
.D(n_152),
.Y(n_167)
);

OAI222xp33_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_65),
.B1(n_134),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_168)
);

NAND4xp25_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_65),
.C(n_101),
.D(n_71),
.Y(n_169)
);

OAI211xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_71),
.B(n_4),
.C(n_6),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_109),
.B(n_82),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.C(n_9),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_161),
.B(n_10),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_173),
.B1(n_170),
.B2(n_169),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_154),
.B(n_160),
.C(n_9),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_12),
.C(n_71),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_154),
.B1(n_116),
.B2(n_12),
.Y(n_178)
);

AND4x2_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_15),
.C(n_16),
.D(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_90),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_20),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_81),
.B1(n_26),
.B2(n_27),
.C(n_24),
.Y(n_182)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_116),
.Y(n_186)
);

AOI222xp33_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_84),
.B1(n_89),
.B2(n_92),
.C1(n_110),
.C2(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_177),
.B(n_182),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_191),
.B1(n_186),
.B2(n_188),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_192),
.B1(n_189),
.B2(n_187),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_194),
.B1(n_189),
.B2(n_179),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_112),
.B(n_89),
.Y(n_197)
);


endmodule