module real_jpeg_4257_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_139),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_58),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_9),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_12),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_13),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_13),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_15),
.Y(n_201)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_145),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_20),
.B(n_123),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.C(n_50),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_126),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_23),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.CI(n_31),
.CON(n_23),
.SN(n_23)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_27),
.C(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_26),
.Y(n_199)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_30),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_34),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_34),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_35),
.A2(n_36),
.B1(n_50),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.C(n_46),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_37),
.A2(n_38),
.B1(n_46),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_43),
.B(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_46),
.Y(n_216)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_55),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_76),
.B2(n_77),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_75),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_100),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.C(n_95),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_96),
.Y(n_143)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_108),
.B1(n_121),
.B2(n_122),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.Y(n_107)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_115),
.Y(n_120)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_142),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_125),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_142),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_134),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_129),
.B(n_130),
.Y(n_209)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_138),
.Y(n_188)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_218),
.B(n_222),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_204),
.B(n_217),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_185),
.B(n_203),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_165),
.B(n_184),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_162),
.B(n_164),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_154),
.Y(n_166)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_176),
.C(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_202),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_202),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.C(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_212),
.C(n_213),
.Y(n_211)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_207),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.C(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_221),
.Y(n_222)
);


endmodule