module fake_jpeg_3394_n_722 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_722);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_722;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_721;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_62),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_64),
.B(n_66),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_68),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_19),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_67),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_8),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_69),
.Y(n_224)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_75),
.B(n_79),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_21),
.B(n_8),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_83),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_9),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_84),
.B(n_87),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_85),
.Y(n_226)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_88),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_90),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_91),
.B(n_105),
.Y(n_221)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_92),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_94),
.B(n_119),
.Y(n_211)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_96),
.Y(n_217)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_100),
.Y(n_232)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_24),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_24),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_117),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx5_ASAP7_75t_SL g203 ( 
.A(n_110),
.Y(n_203)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_111),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_26),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_34),
.B(n_9),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_21),
.B(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_42),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_33),
.Y(n_151)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_43),
.Y(n_134)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_140),
.B(n_141),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_68),
.B(n_57),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_151),
.B(n_209),
.Y(n_301)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_112),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g260 ( 
.A(n_152),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_84),
.B(n_57),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_206),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_60),
.B1(n_56),
.B2(n_48),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_158),
.B(n_180),
.Y(n_287)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_159),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_163),
.B(n_166),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_80),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_172),
.A2(n_205),
.B1(n_77),
.B2(n_63),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_81),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_179),
.B(n_208),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_62),
.B(n_60),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_42),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_183),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g194 ( 
.A(n_110),
.Y(n_194)
);

BUFx4f_ASAP7_75t_SL g294 ( 
.A(n_194),
.Y(n_294)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_130),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_198),
.B(n_2),
.Y(n_296)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_124),
.A2(n_37),
.B1(n_31),
.B2(n_23),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_123),
.B(n_22),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_78),
.B(n_31),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_73),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_225),
.Y(n_270)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_74),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_99),
.A2(n_37),
.B1(n_48),
.B2(n_36),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_113),
.B1(n_115),
.B2(n_97),
.Y(n_234)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_85),
.Y(n_229)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_233),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_234),
.A2(n_274),
.B1(n_306),
.B2(n_201),
.Y(n_318)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_235),
.Y(n_379)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_236),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_0),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_237),
.B(n_259),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_240),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g351 ( 
.A1(n_241),
.A2(n_219),
.B1(n_224),
.B2(n_216),
.Y(n_351)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_242),
.Y(n_357)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_245),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_161),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_249),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_250),
.B(n_275),
.Y(n_325)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx11_ASAP7_75t_L g347 ( 
.A(n_253),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_205),
.A2(n_61),
.B1(n_89),
.B2(n_93),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_254),
.A2(n_261),
.B1(n_304),
.B2(n_169),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_192),
.A2(n_102),
.B1(n_108),
.B2(n_96),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_255),
.A2(n_169),
.B1(n_217),
.B2(n_201),
.Y(n_324)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_258),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_0),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_153),
.A2(n_106),
.B1(n_129),
.B2(n_48),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_231),
.A2(n_111),
.B1(n_92),
.B2(n_86),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

CKINVDCx12_ASAP7_75t_R g264 ( 
.A(n_147),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_182),
.Y(n_265)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_171),
.Y(n_267)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_268),
.Y(n_356)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_271),
.Y(n_330)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_200),
.A2(n_215),
.B1(n_142),
.B2(n_157),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_188),
.B(n_69),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_198),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_276),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_231),
.A2(n_106),
.B1(n_130),
.B2(n_2),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_277),
.A2(n_289),
.B1(n_295),
.B2(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_162),
.B(n_0),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_174),
.B(n_1),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_284),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_285),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_144),
.B(n_1),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_286),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_184),
.B(n_1),
.Y(n_288)
);

NAND2x1_ASAP7_75t_SL g321 ( 
.A(n_288),
.B(n_296),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_191),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_289)
);

BUFx4f_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_145),
.Y(n_292)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_178),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_297),
.B(n_16),
.Y(n_381)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_145),
.Y(n_298)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_170),
.B(n_19),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_150),
.Y(n_300)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_138),
.Y(n_302)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_144),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_158),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_304)
);

CKINVDCx12_ASAP7_75t_R g305 ( 
.A(n_147),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_305),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_222),
.A2(n_230),
.B1(n_176),
.B2(n_199),
.Y(n_306)
);

CKINVDCx12_ASAP7_75t_R g308 ( 
.A(n_160),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_181),
.B(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_310),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_193),
.Y(n_310)
);

INVx4_ASAP7_75t_SL g311 ( 
.A(n_160),
.Y(n_311)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_155),
.B(n_19),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_195),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_189),
.A2(n_165),
.B1(n_217),
.B2(n_154),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_165),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_143),
.Y(n_353)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_176),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_318),
.A2(n_331),
.B1(n_341),
.B2(n_349),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_324),
.A2(n_351),
.B1(n_353),
.B2(n_359),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_247),
.B1(n_259),
.B2(n_252),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_287),
.A2(n_158),
.B1(n_230),
.B2(n_199),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_333),
.A2(n_370),
.B1(n_373),
.B2(n_294),
.Y(n_427)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_335),
.A2(n_377),
.B1(n_253),
.B2(n_248),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_287),
.A2(n_186),
.B1(n_175),
.B2(n_193),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_338),
.A2(n_342),
.B1(n_380),
.B2(n_311),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_237),
.A2(n_212),
.B1(n_164),
.B2(n_149),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_269),
.A2(n_186),
.B1(n_175),
.B2(n_226),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_173),
.B(n_190),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_346),
.A2(n_362),
.B(n_246),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_278),
.A2(n_212),
.B1(n_164),
.B2(n_148),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_354),
.B(n_291),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_234),
.A2(n_190),
.B1(n_185),
.B2(n_195),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_271),
.A2(n_143),
.B(n_160),
.C(n_159),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_149),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_364),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_148),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_288),
.B(n_226),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_367),
.B(n_368),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_274),
.B(n_213),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_306),
.A2(n_213),
.B1(n_171),
.B2(n_136),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_312),
.A2(n_136),
.B1(n_197),
.B2(n_167),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_291),
.A2(n_185),
.B1(n_216),
.B2(n_15),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_374),
.A2(n_332),
.B1(n_273),
.B2(n_246),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_256),
.A2(n_185),
.B1(n_13),
.B2(n_15),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_243),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_381),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_387),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_333),
.A2(n_270),
.B1(n_301),
.B2(n_312),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_401),
.B1(n_406),
.B2(n_412),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_282),
.B1(n_298),
.B2(n_251),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_386),
.Y(n_443)
);

AO22x1_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_266),
.B1(n_282),
.B2(n_292),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_343),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_389),
.B(n_400),
.Y(n_436)
);

OA22x2_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_251),
.B1(n_316),
.B2(n_280),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

INVx4_ASAP7_75t_SL g391 ( 
.A(n_362),
.Y(n_391)
);

INVx13_ASAP7_75t_L g459 ( 
.A(n_391),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_284),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_392),
.A2(n_398),
.B(n_428),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_334),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_404),
.Y(n_437)
);

BUFx12f_ASAP7_75t_SL g394 ( 
.A(n_365),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_394),
.A2(n_396),
.B(n_416),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_321),
.A2(n_346),
.B(n_371),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_266),
.Y(n_398)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_399),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_260),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_352),
.A2(n_317),
.B1(n_303),
.B2(n_239),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_280),
.C(n_238),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_378),
.C(n_376),
.Y(n_449)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_325),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_364),
.B(n_367),
.Y(n_405)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_352),
.A2(n_235),
.B1(n_258),
.B2(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_407),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_343),
.B(n_314),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_411),
.B(n_413),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_363),
.A2(n_307),
.B1(n_293),
.B2(n_267),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_329),
.B(n_257),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_337),
.B(n_329),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_284),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_357),
.B(n_260),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_417),
.B(n_418),
.Y(n_458)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_419),
.B(n_420),
.Y(n_464)
);

INVx13_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_422),
.A2(n_424),
.B(n_350),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_260),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_423),
.B(n_425),
.Y(n_466)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_357),
.B(n_257),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_432),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_431),
.B1(n_330),
.B2(n_376),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_332),
.A2(n_281),
.B(n_272),
.Y(n_428)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_381),
.B(n_238),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_395),
.A2(n_370),
.B1(n_373),
.B2(n_326),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_440),
.A2(n_441),
.B1(n_463),
.B2(n_391),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_395),
.A2(n_351),
.B1(n_356),
.B2(n_327),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_327),
.C(n_356),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_449),
.C(n_460),
.Y(n_481)
);

XOR2x2_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_339),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_405),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_396),
.A2(n_330),
.B(n_328),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_461),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_339),
.B1(n_351),
.B2(n_358),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_456),
.A2(n_471),
.B1(n_422),
.B2(n_421),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_372),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_322),
.B(n_372),
.Y(n_461)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_430),
.A2(n_351),
.B1(n_336),
.B2(n_240),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_402),
.B(n_366),
.C(n_358),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_469),
.C(n_470),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_SL g469 ( 
.A(n_384),
.B(n_366),
.C(n_350),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_405),
.B(n_307),
.C(n_344),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_379),
.B1(n_336),
.B2(n_319),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_392),
.A2(n_348),
.B(n_344),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_398),
.A2(n_348),
.B(n_340),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_389),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_476),
.B(n_491),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_382),
.Y(n_477)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

CKINVDCx12_ASAP7_75t_R g478 ( 
.A(n_448),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_L g540 ( 
.A(n_478),
.B(n_487),
.C(n_506),
.Y(n_540)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_382),
.Y(n_480)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_480),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_500),
.Y(n_518)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_483),
.Y(n_543)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_484),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_464),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_488),
.A2(n_496),
.B1(n_514),
.B2(n_438),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_456),
.A2(n_405),
.B1(n_418),
.B2(n_391),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_498),
.B1(n_502),
.B2(n_455),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_404),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_413),
.Y(n_492)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_454),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_452),
.Y(n_494)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_494),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_428),
.B1(n_411),
.B2(n_432),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_457),
.B(n_412),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_507),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_444),
.A2(n_409),
.B1(n_390),
.B2(n_398),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_406),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_451),
.B(n_393),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_501),
.B(n_504),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_433),
.A2(n_390),
.B1(n_426),
.B2(n_407),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_408),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_410),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_505),
.B(n_470),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_466),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_450),
.B(n_414),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_459),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_294),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_451),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

INVx13_ASAP7_75t_L g511 ( 
.A(n_447),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_511),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_471),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_513),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_445),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_441),
.A2(n_390),
.B1(n_387),
.B2(n_416),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_475),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_387),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_454),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_530),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_500),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_525),
.A2(n_548),
.B1(n_511),
.B2(n_443),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_485),
.A2(n_448),
.B(n_435),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_527),
.A2(n_549),
.B(n_485),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_506),
.B(n_434),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_529),
.B(n_533),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_481),
.B(n_461),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_531),
.B(n_554),
.Y(n_567)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_467),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_513),
.A2(n_433),
.B1(n_458),
.B2(n_455),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_534),
.A2(n_541),
.B1(n_503),
.B2(n_442),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_450),
.Y(n_535)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_535),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_467),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_536),
.B(n_538),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_434),
.Y(n_537)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_425),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_488),
.A2(n_455),
.B1(n_435),
.B2(n_453),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_486),
.B(n_472),
.C(n_473),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_478),
.C(n_507),
.Y(n_561)
);

MAJx2_ASAP7_75t_L g545 ( 
.A(n_493),
.B(n_394),
.C(n_462),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g585 ( 
.A(n_545),
.B(n_399),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_490),
.A2(n_463),
.B1(n_440),
.B2(n_438),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_485),
.A2(n_459),
.B(n_447),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_552),
.A2(n_503),
.B1(n_508),
.B2(n_479),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_486),
.B(n_469),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_502),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_492),
.B(n_442),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_509),
.B(n_397),
.Y(n_555)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_519),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_537),
.Y(n_594)
);

XNOR2x2_ASAP7_75t_SL g593 ( 
.A(n_558),
.B(n_581),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_564),
.C(n_568),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_546),
.A2(n_495),
.B1(n_512),
.B2(n_514),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_562),
.A2(n_565),
.B1(n_573),
.B2(n_574),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_572),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_489),
.C(n_496),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_550),
.A2(n_495),
.B1(n_497),
.B2(n_510),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_386),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_566),
.B(n_589),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_517),
.B(n_489),
.C(n_498),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_519),
.Y(n_569)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_569),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_SL g603 ( 
.A(n_570),
.B(n_585),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_530),
.B(n_495),
.C(n_499),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_577),
.C(n_516),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_482),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_550),
.A2(n_515),
.B1(n_484),
.B2(n_483),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_576),
.A2(n_584),
.B1(n_588),
.B2(n_548),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_524),
.B(n_419),
.C(n_420),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_540),
.B(n_503),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_578),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_420),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_582),
.Y(n_608)
);

FAx1_ASAP7_75t_SL g581 ( 
.A(n_520),
.B(n_511),
.CI(n_399),
.CON(n_581),
.SN(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_521),
.B(n_520),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_583),
.A2(n_551),
.B1(n_544),
.B2(n_543),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_541),
.A2(n_443),
.B1(n_431),
.B2(n_347),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_535),
.B(n_294),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_551),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_534),
.A2(n_320),
.B1(n_379),
.B2(n_262),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_539),
.B(n_320),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g592 ( 
.A1(n_556),
.A2(n_526),
.B(n_525),
.Y(n_592)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_592),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_594),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_560),
.B(n_545),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_596),
.B(n_604),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_539),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_600),
.Y(n_623)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_587),
.Y(n_601)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_601),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_527),
.Y(n_604)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_607),
.Y(n_621)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_579),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_620),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_620),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_549),
.C(n_547),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_611),
.B(n_613),
.Y(n_628)
);

XNOR2x1_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_619),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_564),
.B(n_547),
.C(n_518),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_SL g614 ( 
.A(n_582),
.B(n_518),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_SL g643 ( 
.A(n_614),
.B(n_599),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_523),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_615),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_523),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_616),
.B(n_602),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_617),
.A2(n_618),
.B1(n_588),
.B2(n_543),
.Y(n_640)
);

XOR2x2_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_526),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_561),
.B(n_544),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_598),
.Y(n_626)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_626),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_613),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_611),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_632),
.Y(n_650)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_631),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_610),
.B(n_572),
.C(n_577),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_605),
.B(n_568),
.C(n_580),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_633),
.B(n_635),
.Y(n_666)
);

BUFx12_ASAP7_75t_L g634 ( 
.A(n_608),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_634),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_605),
.B(n_578),
.C(n_574),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_596),
.B(n_585),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_641),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_599),
.B(n_563),
.C(n_569),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_614),
.C(n_586),
.Y(n_654)
);

BUFx24_ASAP7_75t_SL g638 ( 
.A(n_593),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_638),
.B(n_603),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_640),
.A2(n_340),
.B1(n_345),
.B2(n_290),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_593),
.A2(n_558),
.B(n_581),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_604),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_595),
.A2(n_581),
.B(n_559),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_645),
.A2(n_612),
.B(n_532),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_647),
.B(n_663),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_648),
.B(n_623),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_633),
.B(n_619),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_651),
.B(n_653),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_629),
.B(n_608),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_654),
.B(n_658),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_656),
.A2(n_641),
.B(n_645),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_639),
.A2(n_592),
.B1(n_597),
.B2(n_528),
.Y(n_657)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_657),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_637),
.B(n_592),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_624),
.Y(n_659)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_659),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_660),
.B(n_627),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_603),
.C(n_592),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_661),
.B(n_662),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_628),
.B(n_635),
.C(n_627),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_642),
.B(n_528),
.Y(n_663)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_664),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_626),
.A2(n_290),
.B1(n_239),
.B2(n_272),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_665),
.A2(n_622),
.B1(n_623),
.B2(n_644),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_667),
.A2(n_646),
.B1(n_654),
.B2(n_647),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_668),
.B(n_679),
.Y(n_687)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_669),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_643),
.C(n_642),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_675),
.B(n_677),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_648),
.B(n_622),
.C(n_636),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_653),
.B(n_662),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g686 ( 
.A(n_678),
.B(n_651),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_655),
.B(n_639),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_680),
.B(n_661),
.Y(n_685)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_652),
.Y(n_682)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_682),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_649),
.A2(n_625),
.B(n_621),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_683),
.A2(n_665),
.B(n_663),
.Y(n_690)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_684),
.B(n_17),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_685),
.A2(n_680),
.B(n_674),
.Y(n_700)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_686),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_673),
.A2(n_666),
.B(n_625),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_688),
.B(n_691),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_690),
.A2(n_673),
.B(n_670),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_671),
.A2(n_646),
.B1(n_634),
.B2(n_403),
.Y(n_692)
);

XOR2xp5_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_677),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_667),
.A2(n_634),
.B1(n_403),
.B2(n_236),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_SL g705 ( 
.A1(n_694),
.A2(n_672),
.B1(n_696),
.B2(n_693),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g699 ( 
.A(n_695),
.B(n_697),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_678),
.B(n_233),
.Y(n_697)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_698),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_700),
.A2(n_703),
.B(n_707),
.Y(n_710)
);

MAJIxp5_ASAP7_75t_L g702 ( 
.A(n_686),
.B(n_681),
.C(n_676),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_702),
.B(n_704),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_SL g703 ( 
.A1(n_689),
.A2(n_676),
.B(n_683),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g704 ( 
.A(n_691),
.B(n_670),
.C(n_675),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_687),
.Y(n_712)
);

MAJIxp5_ASAP7_75t_L g709 ( 
.A(n_702),
.B(n_685),
.C(n_692),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_712),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_701),
.A2(n_694),
.B(n_700),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g716 ( 
.A(n_713),
.B(n_710),
.Y(n_716)
);

XOR2xp5_ASAP7_75t_L g715 ( 
.A(n_708),
.B(n_704),
.Y(n_715)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_716),
.B(n_701),
.C(n_706),
.Y(n_717)
);

MAJIxp5_ASAP7_75t_L g719 ( 
.A(n_717),
.B(n_714),
.C(n_715),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_718),
.B(n_711),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_720),
.B(n_698),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_721),
.B(n_699),
.Y(n_722)
);


endmodule