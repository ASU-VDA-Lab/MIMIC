module fake_jpeg_2844_n_125 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_38),
.B1(n_39),
.B2(n_32),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_48),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_39),
.B1(n_40),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_45),
.B1(n_56),
.B2(n_52),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_14),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_58),
.B1(n_57),
.B2(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_78),
.B1(n_37),
.B2(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_12),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_51),
.B1(n_43),
.B2(n_40),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_88),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_89),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_1),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_93),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_86),
.B1(n_85),
.B2(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_102),
.B1(n_2),
.B2(n_5),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_71),
.B(n_78),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_15),
.B(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_37),
.B1(n_34),
.B2(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_5),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_98),
.B1(n_95),
.B2(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_109),
.Y(n_116)
);

AO221x1_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_106),
.B1(n_105),
.B2(n_96),
.C(n_104),
.Y(n_110)
);

OAI322xp33_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_112),
.A3(n_30),
.B1(n_17),
.B2(n_16),
.C1(n_9),
.C2(n_10),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_13),
.B(n_26),
.C(n_25),
.D(n_20),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_117),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_108),
.B1(n_112),
.B2(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_116),
.B1(n_118),
.B2(n_115),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_119),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_6),
.B(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_7),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_11),
.Y(n_125)
);


endmodule