module fake_jpeg_15452_n_350 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_38),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_73),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_35),
.B1(n_20),
.B2(n_43),
.Y(n_86)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_18),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_31),
.B1(n_17),
.B2(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_83),
.B1(n_65),
.B2(n_81),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_31),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_100),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_23),
.B1(n_64),
.B2(n_58),
.Y(n_122)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_104),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_90),
.Y(n_115)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_44),
.B1(n_36),
.B2(n_26),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_26),
.B1(n_35),
.B2(n_20),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_29),
.B(n_34),
.C(n_32),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_35),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_59),
.B1(n_65),
.B2(n_63),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_61),
.B1(n_23),
.B2(n_21),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_25),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_120),
.B(n_121),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_122),
.B1(n_132),
.B2(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_27),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_33),
.Y(n_151)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_125),
.B1(n_128),
.B2(n_21),
.Y(n_163)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_27),
.B(n_53),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_96),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_0),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_133),
.B(n_135),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_64),
.B1(n_58),
.B2(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_101),
.B1(n_102),
.B2(n_88),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_78),
.B1(n_87),
.B2(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_53),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_27),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_93),
.B1(n_86),
.B2(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_28),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_89),
.B(n_27),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_98),
.C(n_104),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.C(n_144),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_103),
.C(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_90),
.C(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_159),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_162),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_113),
.B(n_87),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_14),
.B1(n_13),
.B2(n_90),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_123),
.B1(n_115),
.B2(n_3),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_131),
.B(n_120),
.C(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_109),
.B(n_19),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_124),
.B1(n_114),
.B2(n_125),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_133),
.B(n_122),
.C(n_121),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_171),
.B(n_175),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_182),
.B(n_152),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_121),
.B1(n_117),
.B2(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_156),
.B1(n_144),
.B2(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_185),
.B1(n_145),
.B2(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_124),
.B1(n_111),
.B2(n_116),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_139),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_176),
.C(n_183),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_134),
.B(n_107),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_143),
.C(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_115),
.B(n_136),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_132),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_115),
.B1(n_123),
.B2(n_3),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_145),
.B1(n_184),
.B2(n_181),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_21),
.B(n_2),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_159),
.B(n_151),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_192),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_201),
.B1(n_214),
.B2(n_182),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_209),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_198),
.B(n_208),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_137),
.B(n_149),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_123),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_146),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_140),
.B1(n_148),
.B2(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_170),
.B1(n_183),
.B2(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_207),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_137),
.CI(n_154),
.CON(n_209),
.SN(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_150),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_186),
.B1(n_164),
.B2(n_165),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_147),
.B(n_145),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_172),
.Y(n_215)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_25),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_164),
.C(n_176),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_217),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_174),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_222),
.C(n_233),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_227),
.B1(n_237),
.B2(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_175),
.B(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_235),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_171),
.B1(n_166),
.B2(n_165),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_197),
.B1(n_196),
.B2(n_203),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_164),
.C(n_175),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_208),
.C(n_214),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_171),
.B1(n_188),
.B2(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_188),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_234),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_247),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_256),
.B1(n_258),
.B2(n_19),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_193),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_223),
.B1(n_232),
.B2(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_205),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_259),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_226),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_205),
.B1(n_201),
.B2(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_194),
.B1(n_193),
.B2(n_199),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_230),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_211),
.C(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_264),
.C(n_228),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_206),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_215),
.C(n_199),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_231),
.B1(n_240),
.B2(n_237),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_267),
.A2(n_276),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.C(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_239),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_277),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_227),
.CI(n_238),
.CON(n_277),
.SN(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_217),
.B(n_215),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_255),
.B1(n_258),
.B2(n_244),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_19),
.C(n_2),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_19),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_1),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_19),
.C(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_256),
.B1(n_253),
.B2(n_246),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_285),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_1),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_265),
.B1(n_257),
.B2(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_265),
.B1(n_249),
.B2(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_293),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_277),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_272),
.B(n_282),
.C(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_297),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_4),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_SL g305 ( 
.A(n_300),
.B(n_276),
.C(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_278),
.C(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_297),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_308),
.B(n_298),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_277),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_283),
.B1(n_269),
.B2(n_279),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_290),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_295),
.B(n_269),
.CI(n_6),
.CON(n_310),
.SN(n_310)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_311),
.A2(n_303),
.B1(n_313),
.B2(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_298),
.C(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.C(n_299),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_5),
.C(n_6),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_317),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_321),
.B(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_290),
.C(n_301),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_321),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_6),
.C(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_306),
.B1(n_304),
.B2(n_315),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_7),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_311),
.B1(n_8),
.B2(n_10),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_328),
.B(n_11),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_330),
.A2(n_334),
.B(n_320),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_10),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_319),
.A2(n_8),
.B(n_10),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_8),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_323),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_337),
.B(n_340),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_342),
.B(n_331),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_316),
.B(n_10),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_341),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_329),
.A2(n_11),
.B(n_332),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_345),
.B(n_343),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_348),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_330),
.Y(n_350)
);


endmodule