module fake_jpeg_18072_n_51 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_51);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_51;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_28),
.B1(n_8),
.B2(n_12),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_38),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_45),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_13),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_35),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_49),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_14),
.Y(n_51)
);


endmodule