module fake_netlist_5_2578_n_108 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_108);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_108;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2x1p5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_42),
.Y(n_50)
);

NAND2x1p5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_22),
.B1(n_33),
.B2(n_7),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_9),
.B1(n_10),
.B2(n_33),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_46),
.B1(n_40),
.B2(n_44),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_53),
.B1(n_43),
.B2(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_22),
.B1(n_55),
.B2(n_54),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_54),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_46),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_61),
.C(n_45),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_62),
.B(n_63),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_57),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_63),
.B(n_57),
.C(n_40),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_63),
.B(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND4xp25_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_73),
.C(n_65),
.D(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_78),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_74),
.B(n_71),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_81),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_81),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_68),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_11),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_77),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_71),
.B(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_85),
.Y(n_94)
);

AND2x4_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_86),
.B1(n_84),
.B2(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_84),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI211xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_98),
.B(n_99),
.C(n_96),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_102),
.B1(n_96),
.B2(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_40),
.B(n_18),
.C(n_17),
.Y(n_108)
);


endmodule