module fake_jpeg_7491_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_36),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_21),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_19),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_56),
.B1(n_23),
.B2(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_32),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_18),
.B1(n_30),
.B2(n_31),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_25),
.Y(n_66)
);

AOI22x1_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_16),
.B1(n_27),
.B2(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_0),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_54),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_47),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_17),
.B(n_20),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_41),
.C(n_38),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_65),
.B(n_62),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_38),
.B1(n_35),
.B2(n_27),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_45),
.B1(n_52),
.B2(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_51),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_72),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_97),
.B1(n_102),
.B2(n_68),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_98),
.Y(n_118)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_45),
.B1(n_52),
.B2(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_108),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_48),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_86),
.C(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_85),
.B(n_82),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_120),
.B(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_133),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_128),
.B(n_134),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_26),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_91),
.B1(n_106),
.B2(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_105),
.C(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_76),
.B1(n_75),
.B2(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_126),
.B1(n_112),
.B2(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_16),
.B(n_26),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_110),
.C(n_102),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_140),
.C(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_99),
.A3(n_96),
.B1(n_111),
.B2(n_94),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_106),
.C(n_93),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_153),
.C(n_134),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_146),
.B1(n_154),
.B2(n_50),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_113),
.B1(n_127),
.B2(n_122),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_155),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_99),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_99),
.B1(n_109),
.B2(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_130),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_120),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_161),
.C(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_120),
.C(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_27),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_175),
.B1(n_164),
.B2(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_178),
.B1(n_144),
.B2(n_142),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_54),
.B1(n_46),
.B2(n_47),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_185),
.C(n_197),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_135),
.A3(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_138),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_191),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_138),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_50),
.B1(n_35),
.B2(n_4),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_26),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_196),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_184),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_200),
.C(n_205),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_171),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_206),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_178),
.B(n_165),
.C(n_190),
.D(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_179),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_162),
.C(n_166),
.Y(n_208)
);

AOI221xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_175),
.B1(n_166),
.B2(n_181),
.C(n_174),
.Y(n_209)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_5),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_167),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_1),
.B(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_26),
.B(n_6),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_8),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_5),
.B(n_6),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_7),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_7),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_205),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_231),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_229),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_199),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_213),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_220),
.B1(n_222),
.B2(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_223),
.C(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_239),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_8),
.B(n_9),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_226),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_243),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_199),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_235),
.B(n_204),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_226),
.B(n_9),
.C(n_10),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_240),
.C(n_248),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_10),
.C(n_12),
.Y(n_253)
);


endmodule