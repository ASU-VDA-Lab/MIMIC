module fake_jpeg_16624_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_35),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_19),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_49),
.B(n_23),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_20),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_31),
.B(n_30),
.C(n_28),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_36),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_64),
.Y(n_74)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_63),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_46),
.B(n_40),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_30),
.C(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_25),
.Y(n_67)
);

OAI22x1_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_46),
.B1(n_49),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_73),
.B1(n_75),
.B2(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_46),
.B1(n_39),
.B2(n_48),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_46),
.B1(n_39),
.B2(n_49),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_60),
.B(n_67),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_87),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_95),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_61),
.C(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_58),
.B1(n_48),
.B2(n_37),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_75),
.B1(n_82),
.B2(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_98),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_72),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_88),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_81),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_72),
.B1(n_73),
.B2(n_71),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_74),
.B(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_51),
.B1(n_54),
.B2(n_50),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_64),
.B1(n_50),
.B2(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_32),
.B1(n_21),
.B2(n_26),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_118),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_91),
.C(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_98),
.B1(n_96),
.B2(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_108),
.B1(n_109),
.B2(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_33),
.C(n_41),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_33),
.C(n_41),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_20),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_139),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_106),
.B(n_107),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_134),
.C(n_138),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_101),
.C(n_111),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_125),
.B1(n_126),
.B2(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_21),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_47),
.C(n_20),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_122),
.C(n_121),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_132),
.C(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_126),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_133),
.C(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_155),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_129),
.B(n_1),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_3),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_16),
.C(n_1),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_0),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_144),
.B1(n_149),
.B2(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_155),
.B1(n_151),
.B2(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_6),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_156),
.B1(n_150),
.B2(n_9),
.C(n_10),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_165),
.B(n_168),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_170),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_159),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_173),
.B(n_8),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_8),
.Y(n_175)
);


endmodule