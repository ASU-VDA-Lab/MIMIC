module real_aes_1697_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g523 ( .A(n_0), .B(n_220), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_1), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g154 ( .A(n_2), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_3), .B(n_526), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g516 ( .A(n_4), .B(n_175), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_5), .B(n_188), .Y(n_211) );
INVx1_ASAP7_75t_L g508 ( .A(n_6), .Y(n_508) );
INVx1_ASAP7_75t_L g245 ( .A(n_7), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g825 ( .A(n_8), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_9), .Y(n_262) );
AND2x2_ASAP7_75t_L g543 ( .A(n_10), .B(n_144), .Y(n_543) );
INVx2_ASAP7_75t_L g145 ( .A(n_11), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g221 ( .A(n_13), .Y(n_221) );
AOI221x1_ASAP7_75t_L g511 ( .A1(n_14), .A2(n_177), .B1(n_512), .B2(n_514), .C(n_515), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g797 ( .A1(n_14), .A2(n_59), .B1(n_798), .B2(n_799), .Y(n_797) );
INVxp67_ASAP7_75t_L g799 ( .A(n_14), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_15), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_16), .B(n_526), .Y(n_579) );
INVx1_ASAP7_75t_L g119 ( .A(n_17), .Y(n_119) );
INVx1_ASAP7_75t_L g218 ( .A(n_18), .Y(n_218) );
INVx1_ASAP7_75t_SL g166 ( .A(n_19), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_20), .B(n_169), .Y(n_191) );
AOI33xp33_ASAP7_75t_L g236 ( .A1(n_21), .A2(n_49), .A3(n_151), .B1(n_162), .B2(n_237), .B3(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_22), .A2(n_514), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_23), .B(n_220), .Y(n_548) );
AOI221xp5_ASAP7_75t_SL g588 ( .A1(n_24), .A2(n_40), .B1(n_514), .B2(n_526), .C(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g255 ( .A(n_25), .Y(n_255) );
OR2x2_ASAP7_75t_L g146 ( .A(n_26), .B(n_93), .Y(n_146) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_26), .A2(n_93), .B(n_145), .Y(n_179) );
INVxp67_ASAP7_75t_L g510 ( .A(n_27), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_28), .B(n_223), .Y(n_583) );
AND2x2_ASAP7_75t_L g537 ( .A(n_29), .B(n_143), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_30), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_31), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_32), .A2(n_514), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_33), .B(n_223), .Y(n_590) );
AND2x2_ASAP7_75t_L g156 ( .A(n_34), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g161 ( .A(n_34), .Y(n_161) );
AND2x2_ASAP7_75t_L g175 ( .A(n_34), .B(n_154), .Y(n_175) );
OR2x6_ASAP7_75t_L g117 ( .A(n_35), .B(n_118), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g823 ( .A(n_35), .B(n_824), .C(n_826), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_36), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_37), .B(n_149), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_38), .A2(n_178), .B1(n_184), .B2(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_39), .B(n_193), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_41), .A2(n_85), .B1(n_159), .B2(n_514), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_42), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_43), .B(n_220), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_44), .B(n_195), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_45), .B(n_169), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_46), .Y(n_187) );
AND2x2_ASAP7_75t_L g527 ( .A(n_47), .B(n_143), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_48), .B(n_143), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_50), .B(n_169), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_51), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_51), .A2(n_64), .B1(n_434), .B2(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_52), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g152 ( .A(n_53), .Y(n_152) );
INVx1_ASAP7_75t_L g171 ( .A(n_53), .Y(n_171) );
AOI22x1_ASAP7_75t_L g124 ( .A1(n_54), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_54), .Y(n_125) );
AND2x2_ASAP7_75t_L g287 ( .A(n_55), .B(n_143), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_56), .A2(n_78), .B1(n_149), .B2(n_159), .C(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_57), .B(n_149), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_58), .B(n_526), .Y(n_536) );
INVx1_ASAP7_75t_L g798 ( .A(n_59), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_60), .B(n_178), .Y(n_264) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_61), .A2(n_159), .B(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g564 ( .A(n_62), .B(n_143), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_63), .B(n_223), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_64), .Y(n_810) );
INVx1_ASAP7_75t_L g214 ( .A(n_65), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_66), .B(n_220), .Y(n_562) );
AND2x2_ASAP7_75t_SL g584 ( .A(n_67), .B(n_144), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_68), .A2(n_514), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g285 ( .A(n_69), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_70), .B(n_223), .Y(n_549) );
AND2x2_ASAP7_75t_SL g556 ( .A(n_71), .B(n_195), .Y(n_556) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_72), .B(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_73), .A2(n_104), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_73), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_74), .A2(n_159), .B(n_284), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_75), .A2(n_808), .B1(n_809), .B2(n_811), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_75), .Y(n_808) );
INVx1_ASAP7_75t_L g157 ( .A(n_76), .Y(n_157) );
INVx1_ASAP7_75t_L g173 ( .A(n_76), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_77), .B(n_149), .Y(n_239) );
AND2x2_ASAP7_75t_L g176 ( .A(n_79), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g215 ( .A(n_80), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_81), .A2(n_159), .B(n_165), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_82), .A2(n_159), .B(n_190), .C(n_194), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_83), .A2(n_88), .B1(n_149), .B2(n_526), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_84), .B(n_526), .Y(n_563) );
INVx1_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_86), .B(n_119), .Y(n_827) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_87), .B(n_177), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_89), .A2(n_159), .B1(n_234), .B2(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_90), .B(n_220), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_91), .B(n_220), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_92), .A2(n_514), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g202 ( .A(n_94), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_95), .B(n_223), .Y(n_561) );
AND2x2_ASAP7_75t_L g240 ( .A(n_96), .B(n_177), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_97), .A2(n_253), .B(n_254), .C(n_256), .Y(n_252) );
INVxp67_ASAP7_75t_L g513 ( .A(n_98), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_99), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_100), .B(n_223), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_101), .A2(n_514), .B(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g111 ( .A(n_102), .Y(n_111) );
INVx1_ASAP7_75t_SL g795 ( .A(n_102), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_103), .B(n_169), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_104), .Y(n_129) );
AOI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_820), .B(n_828), .Y(n_105) );
AO21x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B(n_793), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_121), .Y(n_112) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x6_ASAP7_75t_SL g498 ( .A(n_116), .B(n_117), .Y(n_498) );
OR2x6_ASAP7_75t_SL g789 ( .A(n_116), .B(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_116), .B(n_790), .Y(n_816) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_116), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_117), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_130), .B2(n_791), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_497), .B1(n_499), .B2(n_787), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_132), .A2(n_497), .B1(n_500), .B2(n_792), .Y(n_791) );
AND3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_491), .C(n_494), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_391), .C(n_421), .D(n_435), .E(n_461), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_135), .A2(n_434), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g804 ( .A(n_135), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_340), .Y(n_135) );
NOR3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_288), .C(n_322), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_205), .B(n_227), .C(n_266), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_180), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_140), .B(n_278), .Y(n_343) );
AND2x2_ASAP7_75t_L g430 ( .A(n_140), .B(n_208), .Y(n_430) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g226 ( .A(n_141), .B(n_197), .Y(n_226) );
INVx1_ASAP7_75t_L g268 ( .A(n_141), .Y(n_268) );
INVx2_ASAP7_75t_L g273 ( .A(n_141), .Y(n_273) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_141), .Y(n_301) );
INVx1_ASAP7_75t_L g315 ( .A(n_141), .Y(n_315) );
AND2x2_ASAP7_75t_L g319 ( .A(n_141), .B(n_210), .Y(n_319) );
AND2x2_ASAP7_75t_L g400 ( .A(n_141), .B(n_209), .Y(n_400) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_176), .Y(n_141) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_142), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_142), .A2(n_558), .B(n_564), .Y(n_557) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_142), .A2(n_531), .B(n_537), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_143), .A2(n_588), .B(n_592), .Y(n_587) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g188 ( .A(n_145), .B(n_146), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_158), .Y(n_147) );
INVx1_ASAP7_75t_L g265 ( .A(n_149), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_149), .A2(n_159), .B1(n_507), .B2(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_155), .Y(n_149) );
INVx1_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
OR2x6_ASAP7_75t_L g167 ( .A(n_151), .B(n_163), .Y(n_167) );
INVxp33_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g164 ( .A(n_152), .B(n_154), .Y(n_164) );
AND2x4_ASAP7_75t_L g223 ( .A(n_152), .B(n_172), .Y(n_223) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g514 ( .A(n_156), .B(n_164), .Y(n_514) );
INVx2_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
AND2x6_ASAP7_75t_L g220 ( .A(n_157), .B(n_170), .Y(n_220) );
INVxp67_ASAP7_75t_L g263 ( .A(n_159), .Y(n_263) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
NOR2x1p5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx1_ASAP7_75t_L g238 ( .A(n_162), .Y(n_238) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_174), .Y(n_165) );
INVx2_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_174), .B(n_202), .C(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_167), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_167), .A2(n_174), .B(n_245), .C(n_246), .Y(n_244) );
INVxp67_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_167), .A2(n_174), .B(n_285), .C(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
AND2x4_ASAP7_75t_L g526 ( .A(n_169), .B(n_175), .Y(n_526) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_172), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_174), .A2(n_191), .B(n_192), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_174), .B(n_188), .Y(n_224) );
INVx1_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_174), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_174), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_174), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_174), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_174), .A2(n_582), .B(n_583), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_174), .A2(n_590), .B(n_591), .Y(n_589) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_177), .A2(n_252), .B1(n_257), .B2(n_258), .Y(n_251) );
INVx3_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_178), .B(n_261), .Y(n_260) );
AOI21x1_ASAP7_75t_L g519 ( .A1(n_178), .A2(n_520), .B(n_527), .Y(n_519) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_179), .Y(n_195) );
AND2x4_ASAP7_75t_SL g180 ( .A(n_181), .B(n_196), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g225 ( .A(n_182), .Y(n_225) );
AND2x2_ASAP7_75t_L g269 ( .A(n_182), .B(n_210), .Y(n_269) );
AND2x2_ASAP7_75t_L g290 ( .A(n_182), .B(n_197), .Y(n_290) );
INVx1_ASAP7_75t_L g313 ( .A(n_182), .Y(n_313) );
AND2x4_ASAP7_75t_L g380 ( .A(n_182), .B(n_209), .Y(n_380) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_189), .Y(n_182) );
NOR3xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .C(n_187), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_188), .A2(n_200), .B(n_204), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_188), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_188), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_188), .B(n_513), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_188), .B(n_216), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_188), .A2(n_545), .B(n_546), .Y(n_544) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_194), .A2(n_232), .B(n_240), .Y(n_231) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_194), .A2(n_232), .B(n_240), .Y(n_295) );
AOI21x1_ASAP7_75t_L g552 ( .A1(n_194), .A2(n_553), .B(n_556), .Y(n_552) );
INVx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_195), .A2(n_243), .B(n_247), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_195), .A2(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g396 ( .A(n_196), .B(n_313), .Y(n_396) );
OR2x2_ASAP7_75t_L g437 ( .A(n_196), .B(n_438), .Y(n_437) );
NOR2xp67_ASAP7_75t_SL g456 ( .A(n_196), .B(n_329), .Y(n_456) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_196), .B(n_388), .Y(n_474) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2x1_ASAP7_75t_SL g274 ( .A(n_197), .B(n_210), .Y(n_274) );
AND2x4_ASAP7_75t_L g312 ( .A(n_197), .B(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_197), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_197), .B(n_272), .Y(n_350) );
INVx2_ASAP7_75t_L g364 ( .A(n_197), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_197), .B(n_316), .Y(n_386) );
AND2x2_ASAP7_75t_L g478 ( .A(n_197), .B(n_336), .Y(n_478) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2x1_ASAP7_75t_L g206 ( .A(n_207), .B(n_226), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_208), .B(n_315), .Y(n_329) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_208), .B(n_318), .Y(n_338) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_225), .Y(n_208) );
INVx1_ASAP7_75t_L g316 ( .A(n_209), .Y(n_316) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g336 ( .A(n_210), .Y(n_336) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_217), .B(n_224), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_216), .B(n_255), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B1(n_221), .B2(n_222), .Y(n_217) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVxp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g369 ( .A(n_225), .Y(n_369) );
INVx2_ASAP7_75t_SL g414 ( .A(n_226), .Y(n_414) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_248), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_229), .B(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_L g360 ( .A(n_229), .Y(n_360) );
AND2x2_ASAP7_75t_L g484 ( .A(n_229), .B(n_309), .Y(n_484) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_241), .Y(n_229) );
AND2x4_ASAP7_75t_L g297 ( .A(n_230), .B(n_279), .Y(n_297) );
INVx1_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
AND2x2_ASAP7_75t_L g339 ( .A(n_230), .B(n_294), .Y(n_339) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_231), .B(n_242), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_231), .B(n_280), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_233), .B(n_239), .Y(n_232) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVxp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g277 ( .A(n_242), .Y(n_277) );
AND2x4_ASAP7_75t_L g345 ( .A(n_242), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g357 ( .A(n_242), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_242), .Y(n_399) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_242), .Y(n_411) );
AND2x2_ASAP7_75t_L g427 ( .A(n_242), .B(n_250), .Y(n_427) );
BUFx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g374 ( .A(n_249), .B(n_332), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_249), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_249), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g276 ( .A(n_250), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
INVx2_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_250), .B(n_280), .Y(n_325) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_258), .A2(n_281), .B(n_287), .Y(n_280) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_281), .B(n_287), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B1(n_264), .B2(n_265), .Y(n_259) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_275), .Y(n_266) );
INVx1_ASAP7_75t_L g406 ( .A(n_267), .Y(n_406) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g326 ( .A(n_269), .Y(n_326) );
AND2x2_ASAP7_75t_L g382 ( .A(n_269), .B(n_318), .Y(n_382) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx1_ASAP7_75t_L g296 ( .A(n_271), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_271), .B(n_312), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_271), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g403 ( .A(n_271), .B(n_396), .Y(n_403) );
AND2x2_ASAP7_75t_L g477 ( .A(n_271), .B(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_272), .Y(n_465) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_273), .Y(n_385) );
AND2x2_ASAP7_75t_L g298 ( .A(n_274), .B(n_299), .Y(n_298) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_274), .A2(n_487), .B(n_489), .Y(n_486) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx3_ASAP7_75t_L g372 ( .A(n_276), .Y(n_372) );
NAND2x1_ASAP7_75t_SL g416 ( .A(n_276), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g419 ( .A(n_276), .B(n_297), .Y(n_419) );
AND2x2_ASAP7_75t_L g331 ( .A(n_278), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g468 ( .A(n_278), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g479 ( .A(n_278), .B(n_427), .Y(n_479) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_279), .B(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g410 ( .A(n_280), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_302), .B(n_305), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_297), .B2(n_298), .Y(n_289) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
AND2x2_ASAP7_75t_L g320 ( .A(n_292), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g426 ( .A(n_292), .B(n_427), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_292), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_292), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_294), .B(n_310), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_294), .B(n_310), .Y(n_390) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_294), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g346 ( .A(n_295), .Y(n_346) );
AND2x2_ASAP7_75t_L g354 ( .A(n_295), .B(n_310), .Y(n_354) );
INVx1_ASAP7_75t_L g417 ( .A(n_295), .Y(n_417) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_300), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g447 ( .A(n_303), .B(n_332), .Y(n_447) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
AND2x2_ASAP7_75t_L g344 ( .A(n_304), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g432 ( .A(n_304), .B(n_339), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_311), .B1(n_317), .B2(n_320), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g440 ( .A(n_307), .B(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g470 ( .A(n_310), .B(n_357), .Y(n_470) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g337 ( .A(n_312), .Y(n_337) );
OAI21xp33_ASAP7_75t_SL g483 ( .A1(n_312), .A2(n_484), .B(n_485), .Y(n_483) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_315), .Y(n_473) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_SL g415 ( .A1(n_318), .A2(n_416), .B(n_418), .C(n_420), .Y(n_415) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_319), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g420 ( .A(n_319), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_319), .B(n_396), .Y(n_460) );
INVx1_ASAP7_75t_SL g327 ( .A(n_320), .Y(n_327) );
AND2x2_ASAP7_75t_L g408 ( .A(n_321), .B(n_345), .Y(n_408) );
INVx1_ASAP7_75t_L g453 ( .A(n_321), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B1(n_327), .B2(n_328), .C(n_330), .Y(n_322) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_323), .Y(n_442) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g490 ( .A(n_325), .B(n_333), .Y(n_490) );
OR2x2_ASAP7_75t_L g349 ( .A(n_326), .B(n_350), .Y(n_349) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_326), .B(n_363), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_326), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g488 ( .A(n_326), .B(n_385), .Y(n_488) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI32xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .A3(n_337), .B1(n_338), .B2(n_339), .Y(n_330) );
INVx1_ASAP7_75t_L g351 ( .A(n_332), .Y(n_351) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_334), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g446 ( .A(n_335), .Y(n_446) );
OAI22xp33_ASAP7_75t_SL g428 ( .A1(n_337), .A2(n_429), .B1(n_431), .B2(n_433), .Y(n_428) );
INVx1_ASAP7_75t_L g459 ( .A(n_338), .Y(n_459) );
AOI211x1_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B(n_348), .C(n_365), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_342), .B(n_427), .Y(n_433) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g389 ( .A(n_345), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g455 ( .A(n_345), .Y(n_455) );
OAI222xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_352), .B2(n_358), .C1(n_359), .C2(n_361), .Y(n_348) );
INVxp67_ASAP7_75t_L g445 ( .A(n_349), .Y(n_445) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_353), .B(n_438), .Y(n_485) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g401 ( .A(n_354), .B(n_398), .Y(n_401) );
INVx3_ASAP7_75t_L g441 ( .A(n_356), .Y(n_441) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_364), .B(n_380), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B1(n_373), .B2(n_378), .C(n_381), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_367), .A2(n_424), .B(n_426), .Y(n_423) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g377 ( .A(n_371), .Y(n_377) );
OR2x2_ASAP7_75t_L g481 ( .A(n_372), .B(n_417), .Y(n_481) );
NOR2xp67_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_375), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_378), .A2(n_407), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_379), .A2(n_451), .B(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g388 ( .A(n_380), .Y(n_388) );
OAI31xp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_383), .A3(n_387), .B(n_389), .Y(n_381) );
INVx1_ASAP7_75t_L g439 ( .A(n_383), .Y(n_439) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_404), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_392), .B(n_404), .C(n_423), .D(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_402), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B1(n_400), .B2(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g464 ( .A(n_396), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_397), .B(n_417), .Y(n_425) );
INVx1_ASAP7_75t_SL g438 ( .A(n_400), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_415), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_409), .B2(n_412), .Y(n_405) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_414), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_476) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_428), .C(n_434), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g493 ( .A(n_428), .Y(n_493) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_434), .A2(n_495), .B(n_496), .Y(n_494) );
INVxp33_ASAP7_75t_L g495 ( .A(n_435), .Y(n_495) );
AND2x2_ASAP7_75t_L g803 ( .A(n_435), .B(n_461), .Y(n_803) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_436), .B(n_443), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_440), .A2(n_463), .B(n_466), .Y(n_462) );
INVx2_ASAP7_75t_L g450 ( .A(n_441), .Y(n_450) );
NAND3xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_448), .C(n_457), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B1(n_454), .B2(n_456), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVxp33_ASAP7_75t_SL g496 ( .A(n_461), .Y(n_496) );
NOR3x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_475), .C(n_482), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_483), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g805 ( .A(n_492), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_664), .Y(n_500) );
NOR4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_607), .C(n_646), .D(n_653), .Y(n_501) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_528), .B1(n_565), .B2(n_574), .C(n_593), .Y(n_502) );
OR2x2_ASAP7_75t_L g737 ( .A(n_503), .B(n_599), .Y(n_737) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g652 ( .A(n_504), .B(n_577), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_504), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_504), .B(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_517), .Y(n_504) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_505), .B(n_577), .Y(n_576) );
INVx3_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
AND2x2_ASAP7_75t_L g633 ( .A(n_505), .B(n_606), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_505), .B(n_518), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_505), .B(n_600), .Y(n_685) );
OR2x2_ASAP7_75t_L g763 ( .A(n_505), .B(n_577), .Y(n_763) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_518), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g611 ( .A(n_518), .Y(n_611) );
OR2x2_ASAP7_75t_L g616 ( .A(n_518), .B(n_600), .Y(n_616) );
AND2x2_ASAP7_75t_L g629 ( .A(n_518), .B(n_587), .Y(n_629) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_518), .Y(n_632) );
INVx1_ASAP7_75t_L g644 ( .A(n_518), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_518), .B(n_598), .Y(n_709) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_538), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g573 ( .A(n_530), .B(n_557), .Y(n_573) );
AND2x4_ASAP7_75t_L g603 ( .A(n_530), .B(n_542), .Y(n_603) );
INVx2_ASAP7_75t_L g637 ( .A(n_530), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_530), .B(n_557), .Y(n_695) );
AND2x2_ASAP7_75t_L g742 ( .A(n_530), .B(n_571), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_538), .A2(n_602), .B1(n_645), .B2(n_705), .C1(n_731), .C2(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_550), .Y(n_539) );
AND2x2_ASAP7_75t_L g649 ( .A(n_540), .B(n_569), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_540), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g778 ( .A(n_540), .B(n_618), .Y(n_778) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_541), .A2(n_609), .B(n_613), .Y(n_608) );
AND2x2_ASAP7_75t_L g689 ( .A(n_541), .B(n_572), .Y(n_689) );
OR2x2_ASAP7_75t_L g714 ( .A(n_541), .B(n_573), .Y(n_714) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx5_ASAP7_75t_L g568 ( .A(n_542), .Y(n_568) );
AND2x2_ASAP7_75t_L g655 ( .A(n_542), .B(n_637), .Y(n_655) );
AND2x2_ASAP7_75t_L g681 ( .A(n_542), .B(n_557), .Y(n_681) );
OR2x2_ASAP7_75t_L g684 ( .A(n_542), .B(n_571), .Y(n_684) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_542), .Y(n_702) );
AND2x4_ASAP7_75t_SL g759 ( .A(n_542), .B(n_636), .Y(n_759) );
OR2x2_ASAP7_75t_L g768 ( .A(n_542), .B(n_595), .Y(n_768) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
AOI221xp5_ASAP7_75t_SL g719 ( .A1(n_550), .A2(n_603), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_719) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
OR2x2_ASAP7_75t_L g658 ( .A(n_551), .B(n_628), .Y(n_658) );
OR2x2_ASAP7_75t_L g668 ( .A(n_551), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g694 ( .A(n_551), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g700 ( .A(n_551), .B(n_619), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_551), .B(n_683), .Y(n_712) );
INVx2_ASAP7_75t_L g725 ( .A(n_551), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_551), .B(n_603), .Y(n_746) );
AND2x2_ASAP7_75t_L g750 ( .A(n_551), .B(n_572), .Y(n_750) );
AND2x2_ASAP7_75t_L g758 ( .A(n_551), .B(n_759), .Y(n_758) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_557), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g602 ( .A(n_557), .B(n_571), .Y(n_602) );
INVx2_ASAP7_75t_L g619 ( .A(n_557), .Y(n_619) );
AND2x4_ASAP7_75t_L g636 ( .A(n_557), .B(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_557), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g748 ( .A(n_567), .B(n_570), .Y(n_748) );
AND2x4_ASAP7_75t_L g594 ( .A(n_568), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g635 ( .A(n_568), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g662 ( .A(n_568), .B(n_602), .Y(n_662) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g766 ( .A(n_570), .B(n_767), .Y(n_766) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g618 ( .A(n_571), .B(n_619), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_572), .A2(n_639), .B(n_645), .Y(n_638) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_585), .Y(n_575) );
INVx1_ASAP7_75t_SL g692 ( .A(n_576), .Y(n_692) );
AND2x2_ASAP7_75t_L g722 ( .A(n_576), .B(n_632), .Y(n_722) );
AND2x4_ASAP7_75t_L g733 ( .A(n_576), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g599 ( .A(n_577), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g606 ( .A(n_577), .Y(n_606) );
AND2x4_ASAP7_75t_L g612 ( .A(n_577), .B(n_598), .Y(n_612) );
INVx2_ASAP7_75t_L g623 ( .A(n_577), .Y(n_623) );
INVx1_ASAP7_75t_L g672 ( .A(n_577), .Y(n_672) );
OR2x2_ASAP7_75t_L g693 ( .A(n_577), .B(n_677), .Y(n_693) );
OR2x2_ASAP7_75t_L g707 ( .A(n_577), .B(n_587), .Y(n_707) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_577), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_577), .B(n_629), .Y(n_779) );
OR2x6_ASAP7_75t_L g577 ( .A(n_578), .B(n_584), .Y(n_577) );
INVx1_ASAP7_75t_L g624 ( .A(n_585), .Y(n_624) );
AND2x2_ASAP7_75t_L g757 ( .A(n_585), .B(n_623), .Y(n_757) );
AND2x2_ASAP7_75t_L g782 ( .A(n_585), .B(n_612), .Y(n_782) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g600 ( .A(n_587), .Y(n_600) );
BUFx3_ASAP7_75t_L g642 ( .A(n_587), .Y(n_642) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
INVx1_ASAP7_75t_L g678 ( .A(n_587), .Y(n_678) );
AOI33xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .A3(n_601), .B1(n_602), .B2(n_603), .B3(n_604), .Y(n_593) );
AOI21x1_ASAP7_75t_SL g696 ( .A1(n_594), .A2(n_618), .B(n_680), .Y(n_696) );
INVx2_ASAP7_75t_L g726 ( .A(n_594), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_594), .B(n_725), .Y(n_732) );
AND2x2_ASAP7_75t_L g680 ( .A(n_595), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g643 ( .A(n_598), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g744 ( .A(n_599), .Y(n_744) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_600), .Y(n_734) );
OAI32xp33_ASAP7_75t_L g783 ( .A1(n_601), .A2(n_603), .A3(n_779), .B1(n_784), .B2(n_786), .Y(n_783) );
AND2x2_ASAP7_75t_L g701 ( .A(n_602), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g691 ( .A(n_603), .Y(n_691) );
AND2x2_ASAP7_75t_L g756 ( .A(n_603), .B(n_700), .Y(n_756) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_617), .B1(n_620), .B2(n_634), .C(n_638), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_611), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_612), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_612), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_612), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g661 ( .A(n_616), .Y(n_661) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .C(n_630), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_622), .A2(n_684), .B1(n_724), .B2(n_727), .Y(n_723) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g627 ( .A(n_623), .Y(n_627) );
NOR2x1p5_ASAP7_75t_L g641 ( .A(n_623), .B(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_623), .Y(n_663) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g690 ( .A1(n_626), .A2(n_668), .A3(n_691), .B1(n_692), .B2(n_693), .C1(n_694), .C2(n_696), .Y(n_690) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_628), .A2(n_647), .B(n_648), .C(n_650), .Y(n_646) );
OR2x2_ASAP7_75t_L g738 ( .A(n_628), .B(n_692), .Y(n_738) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g645 ( .A(n_629), .B(n_633), .Y(n_645) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g651 ( .A(n_635), .B(n_652), .Y(n_651) );
INVx3_ASAP7_75t_SL g683 ( .A(n_636), .Y(n_683) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_640), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_SL g687 ( .A(n_643), .Y(n_687) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_644), .Y(n_729) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_647), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g774 ( .A1(n_652), .A2(n_775), .B(n_776), .C(n_783), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_659), .C(n_663), .Y(n_653) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_654), .A2(n_666), .B(n_673), .C(n_697), .Y(n_665) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_710), .C(n_754), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_669), .Y(n_761) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g716 ( .A(n_672), .Y(n_716) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_686), .C(n_690), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B1(n_682), .B2(n_685), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g718 ( .A(n_678), .Y(n_718) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_678), .Y(n_785) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_SL g771 ( .A(n_684), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OR2x2_ASAP7_75t_L g721 ( .A(n_687), .B(n_707), .Y(n_721) );
OR2x2_ASAP7_75t_L g772 ( .A(n_687), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g770 ( .A(n_695), .Y(n_770) );
OR2x2_ASAP7_75t_L g786 ( .A(n_695), .B(n_725), .Y(n_786) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B(n_703), .Y(n_697) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_698), .A2(n_712), .A3(n_713), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g743 ( .A(n_708), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND4xp25_ASAP7_75t_SL g710 ( .A(n_711), .B(n_719), .C(n_730), .D(n_735), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_718), .Y(n_753) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_739), .B1(n_743), .B2(n_745), .C(n_747), .Y(n_735) );
NAND2xp33_ASAP7_75t_SL g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g780 ( .A(n_739), .Y(n_780) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g775 ( .A(n_749), .Y(n_775) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_755), .B(n_774), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_758), .B2(n_760), .C(n_764), .Y(n_755) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
AOI21xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_769), .B(n_772), .Y(n_764) );
INVxp33_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_788), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_796), .B(n_817), .Y(n_793) );
INVx2_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_800), .B(n_812), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_797), .A2(n_813), .B(n_814), .Y(n_812) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g813 ( .A(n_801), .Y(n_813) );
XNOR2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_806), .Y(n_801) );
NAND3x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .C(n_805), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g811 ( .A(n_809), .Y(n_811) );
CKINVDCx11_ASAP7_75t_R g819 ( .A(n_814), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
BUFx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
BUFx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
BUFx4f_ASAP7_75t_SL g831 ( .A(n_822), .Y(n_831) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_823), .B(n_827), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
endmodule