module fake_jpeg_12202_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_78),
.Y(n_91)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_76),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_103),
.B(n_55),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_85),
.B1(n_84),
.B2(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_100),
.B1(n_102),
.B2(n_72),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_69),
.B1(n_62),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_69),
.B1(n_64),
.B2(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_65),
.B1(n_63),
.B2(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_125),
.Y(n_144)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_53),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_67),
.B1(n_52),
.B2(n_58),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_122),
.B1(n_118),
.B2(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_3),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_0),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_138),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_136),
.B1(n_11),
.B2(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_1),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_26),
.C(n_50),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_9),
.C(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_4),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_130),
.B(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_157),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_142),
.B1(n_19),
.B2(n_20),
.C(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_154),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_7),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_9),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_10),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_17),
.B1(n_29),
.B2(n_32),
.Y(n_178)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_142),
.B1(n_24),
.B2(n_27),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_15),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_139),
.C(n_132),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_154),
.C(n_160),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_164),
.C(n_35),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_158),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.C(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_185),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_162),
.C(n_40),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_34),
.C(n_42),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_187),
.C(n_186),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_177),
.B(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_172),
.C(n_182),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_195),
.B(n_174),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_168),
.Y(n_197)
);


endmodule