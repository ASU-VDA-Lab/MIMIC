module real_aes_7872_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_734, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_734;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g481 ( .A1(n_0), .A2(n_186), .B(n_482), .C(n_485), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_1), .A2(n_105), .B1(n_435), .B2(n_444), .C(n_447), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_1), .A2(n_108), .B1(n_109), .B2(n_424), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_1), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_1), .B(n_476), .Y(n_486) );
INVx1_ASAP7_75t_L g430 ( .A(n_2), .Y(n_430) );
INVx1_ASAP7_75t_L g221 ( .A(n_3), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_4), .B(n_138), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_471), .B(n_559), .Y(n_558) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_6), .A2(n_161), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_7), .A2(n_37), .B1(n_131), .B2(n_155), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_8), .B(n_161), .Y(n_233) );
AND2x6_ASAP7_75t_L g146 ( .A(n_9), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_10), .A2(n_146), .B(n_462), .C(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_11), .B(n_38), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g110 ( .A1(n_12), .A2(n_76), .B1(n_111), .B2(n_112), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_14), .B(n_136), .Y(n_169) );
INVx1_ASAP7_75t_L g213 ( .A(n_15), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_16), .B(n_138), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_17), .B(n_162), .Y(n_200) );
AO32x2_ASAP7_75t_L g183 ( .A1(n_18), .A2(n_160), .A3(n_161), .B1(n_184), .B2(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_19), .B(n_131), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_20), .B(n_162), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_21), .A2(n_56), .B1(n_131), .B2(n_155), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g158 ( .A1(n_22), .A2(n_82), .B1(n_131), .B2(n_136), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_23), .B(n_131), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_24), .A2(n_160), .B(n_462), .C(n_509), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_25), .A2(n_160), .B(n_462), .C(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_27), .B(n_123), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_28), .A2(n_94), .B1(n_719), .B2(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_28), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_29), .A2(n_717), .B1(n_718), .B2(n_721), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_29), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_30), .A2(n_471), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_31), .B(n_123), .Y(n_148) );
INVx2_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_33), .A2(n_468), .B(n_494), .C(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_34), .B(n_131), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_35), .B(n_123), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_36), .B(n_171), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_39), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_40), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_41), .A2(n_93), .B1(n_136), .B2(n_137), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_42), .B(n_138), .Y(n_547) );
OAI22xp5_ASAP7_75t_SL g420 ( .A1(n_43), .A2(n_103), .B1(n_421), .B2(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_43), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_43), .A2(n_114), .B1(n_422), .B2(n_423), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_44), .B(n_471), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_45), .B(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_46), .A2(n_468), .B(n_494), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_47), .B(n_131), .Y(n_228) );
INVx1_ASAP7_75t_L g483 ( .A(n_48), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_49), .A2(n_91), .B1(n_155), .B2(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g546 ( .A(n_50), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_51), .B(n_131), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_131), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_53), .A2(n_715), .B1(n_716), .B2(n_722), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_53), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_54), .B(n_471), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_55), .B(n_219), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_57), .A2(n_61), .B1(n_131), .B2(n_136), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_58), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_59), .B(n_131), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_60), .B(n_131), .Y(n_241) );
INVx1_ASAP7_75t_L g147 ( .A(n_62), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_63), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_64), .B(n_476), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_65), .A2(n_216), .B(n_219), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_66), .B(n_131), .Y(n_222) );
INVx1_ASAP7_75t_L g126 ( .A(n_67), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_68), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_69), .B(n_138), .Y(n_499) );
AO32x2_ASAP7_75t_L g152 ( .A1(n_70), .A2(n_153), .A3(n_159), .B1(n_160), .B2(n_161), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_71), .B(n_139), .Y(n_536) );
INVx1_ASAP7_75t_L g240 ( .A(n_72), .Y(n_240) );
INVx1_ASAP7_75t_L g134 ( .A(n_73), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_74), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_75), .B(n_498), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_77), .A2(n_462), .B(n_464), .C(n_468), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_78), .B(n_136), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_79), .Y(n_560) );
INVx1_ASAP7_75t_L g443 ( .A(n_80), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_81), .B(n_497), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_83), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_84), .B(n_155), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_85), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_86), .B(n_136), .Y(n_143) );
INVx2_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_88), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_89), .B(n_157), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_90), .B(n_136), .Y(n_229) );
OR2x2_ASAP7_75t_L g427 ( .A(n_92), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g452 ( .A(n_92), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_94), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_95), .B(n_471), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_96), .Y(n_496) );
INVxp67_ASAP7_75t_L g563 ( .A(n_97), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_98), .B(n_136), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_99), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g465 ( .A(n_100), .Y(n_465) );
INVx1_ASAP7_75t_L g532 ( .A(n_101), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_102), .B(n_123), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_103), .Y(n_421) );
OAI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_425), .B(n_432), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
XNOR2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_113), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_419), .B1(n_420), .B2(n_423), .Y(n_113) );
INVx1_ASAP7_75t_L g423 ( .A(n_114), .Y(n_423) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_340), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_289), .C(n_331), .Y(n_115) );
AOI211xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_194), .B(n_243), .C(n_265), .Y(n_116) );
OAI211xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_149), .B(n_177), .C(n_189), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_119), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g352 ( .A(n_119), .B(n_269), .Y(n_352) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g254 ( .A(n_120), .B(n_180), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_120), .B(n_165), .Y(n_371) );
INVx1_ASAP7_75t_L g389 ( .A(n_120), .Y(n_389) );
AND2x2_ASAP7_75t_L g398 ( .A(n_120), .B(n_286), .Y(n_398) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g281 ( .A(n_121), .B(n_165), .Y(n_281) );
AND2x2_ASAP7_75t_L g339 ( .A(n_121), .B(n_286), .Y(n_339) );
INVx1_ASAP7_75t_L g383 ( .A(n_121), .Y(n_383) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g260 ( .A(n_122), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g268 ( .A(n_122), .Y(n_268) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_122), .Y(n_308) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_148), .Y(n_122) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_123), .A2(n_166), .B(n_176), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_123), .A2(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g515 ( .A(n_123), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_123), .A2(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_L g162 ( .A(n_124), .B(n_125), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_141), .B(n_146), .Y(n_128) );
O2A1O1Ixp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_134), .B(n_135), .C(n_138), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_131), .Y(n_467) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_132), .Y(n_156) );
AND2x6_ASAP7_75t_L g462 ( .A(n_132), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_133), .Y(n_137) );
INVx1_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
INVx2_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_138), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_138), .A2(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_138), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_139), .A2(n_154), .B1(n_157), .B2(n_158), .Y(n_153) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
INVx1_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g463 ( .A(n_140), .Y(n_463) );
AND2x2_ASAP7_75t_L g472 ( .A(n_140), .B(n_220), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g498 ( .A(n_145), .Y(n_498) );
BUFx3_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_146), .A2(n_167), .B(n_172), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_146), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_146), .A2(n_227), .B(n_230), .Y(n_226) );
INVx4_ASAP7_75t_SL g469 ( .A(n_146), .Y(n_469) );
AND2x4_ASAP7_75t_L g471 ( .A(n_146), .B(n_472), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_146), .B(n_472), .Y(n_533) );
INVxp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_163), .Y(n_150) );
AND2x2_ASAP7_75t_L g247 ( .A(n_151), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g280 ( .A(n_151), .Y(n_280) );
OR2x2_ASAP7_75t_L g406 ( .A(n_151), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_151), .B(n_165), .Y(n_410) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
AND2x2_ASAP7_75t_L g269 ( .A(n_152), .B(n_182), .Y(n_269) );
AND2x2_ASAP7_75t_L g309 ( .A(n_152), .B(n_183), .Y(n_309) );
INVx2_ASAP7_75t_L g485 ( .A(n_156), .Y(n_485) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_156), .Y(n_500) );
INVx2_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_157), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_157), .A2(n_186), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx4_ASAP7_75t_L g484 ( .A(n_157), .Y(n_484) );
INVx1_ASAP7_75t_L g512 ( .A(n_159), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_160), .B(n_202), .C(n_205), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_160), .A2(n_236), .B(n_239), .Y(n_235) );
INVx4_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_161), .A2(n_226), .B(n_233), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_161), .A2(n_522), .B(n_523), .Y(n_521) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_161), .Y(n_557) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVxp67_ASAP7_75t_L g351 ( .A(n_163), .Y(n_351) );
AND2x4_ASAP7_75t_L g376 ( .A(n_163), .B(n_269), .Y(n_376) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_164), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g181 ( .A(n_165), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g255 ( .A(n_165), .B(n_183), .Y(n_255) );
INVx1_ASAP7_75t_L g261 ( .A(n_165), .Y(n_261) );
INVx2_ASAP7_75t_L g287 ( .A(n_165), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_165), .B(n_304), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_175), .A2(n_218), .B(n_240), .C(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_178), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
AND2x2_ASAP7_75t_L g366 ( .A(n_180), .B(n_182), .Y(n_366) );
AND2x2_ASAP7_75t_L g283 ( .A(n_181), .B(n_268), .Y(n_283) );
AND2x2_ASAP7_75t_L g382 ( .A(n_181), .B(n_383), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_182), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g407 ( .A(n_182), .B(n_268), .Y(n_407) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g193 ( .A(n_183), .Y(n_193) );
AND2x2_ASAP7_75t_L g286 ( .A(n_183), .B(n_287), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_218), .B(n_221), .C(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_186), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g210 ( .A(n_188), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_188), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
AND2x2_ASAP7_75t_L g332 ( .A(n_191), .B(n_267), .Y(n_332) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_192), .B(n_268), .Y(n_317) );
INVx2_ASAP7_75t_L g316 ( .A(n_193), .Y(n_316) );
OAI222xp33_ASAP7_75t_L g320 ( .A1(n_193), .A2(n_260), .B1(n_321), .B2(n_323), .C1(n_324), .C2(n_327), .Y(n_320) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
OR2x2_ASAP7_75t_L g356 ( .A(n_198), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g278 ( .A(n_199), .Y(n_278) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_199), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g335 ( .A(n_199), .B(n_249), .Y(n_335) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
AO21x1_ASAP7_75t_L g295 ( .A1(n_202), .A2(n_205), .B(n_296), .Y(n_295) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_205), .A2(n_460), .B(n_473), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_205), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g476 ( .A(n_205), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_205), .B(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_205), .A2(n_531), .B(n_538), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_206), .A2(n_299), .B1(n_338), .B2(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_224), .Y(n_206) );
INVx3_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
OR2x2_ASAP7_75t_L g404 ( .A(n_207), .B(n_280), .Y(n_404) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g277 ( .A(n_208), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g293 ( .A(n_208), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_208), .B(n_249), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_208), .B(n_225), .Y(n_357) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g252 ( .A(n_209), .B(n_225), .Y(n_252) );
AND2x2_ASAP7_75t_L g328 ( .A(n_209), .B(n_275), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_209), .B(n_234), .Y(n_368) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_223), .Y(n_209) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_210), .A2(n_235), .B(n_242), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .C(n_216), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_214), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_214), .A2(n_536), .B(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_216), .A2(n_465), .B(n_466), .C(n_467), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_218), .A2(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_224), .B(n_245), .Y(n_284) );
AND2x2_ASAP7_75t_L g288 ( .A(n_224), .B(n_278), .Y(n_288) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
INVx3_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_225), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g409 ( .A(n_225), .B(n_392), .Y(n_409) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
INVx2_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
AND2x2_ASAP7_75t_L g319 ( .A(n_234), .B(n_295), .Y(n_319) );
INVx1_ASAP7_75t_L g362 ( .A(n_234), .Y(n_362) );
OR2x2_ASAP7_75t_L g393 ( .A(n_234), .B(n_295), .Y(n_393) );
AND2x2_ASAP7_75t_L g413 ( .A(n_234), .B(n_249), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g251 ( .A(n_245), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_245), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g370 ( .A(n_247), .Y(n_370) );
INVx2_ASAP7_75t_SL g264 ( .A(n_248), .Y(n_264) );
AND2x2_ASAP7_75t_L g384 ( .A(n_248), .B(n_278), .Y(n_384) );
INVx2_ASAP7_75t_L g330 ( .A(n_249), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_249), .B(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B1(n_256), .B2(n_262), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_252), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g418 ( .A(n_252), .Y(n_418) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g343 ( .A(n_254), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_254), .B(n_286), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_255), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_308), .Y(n_359) );
INVx2_ASAP7_75t_L g415 ( .A(n_255), .Y(n_415) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g285 ( .A(n_258), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_258), .B(n_303), .Y(n_336) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_260), .B(n_280), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g347 ( .A1(n_264), .A2(n_348), .B(n_350), .C(n_353), .Y(n_347) );
OR2x2_ASAP7_75t_L g374 ( .A(n_264), .B(n_278), .Y(n_374) );
OAI221xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_270), .B1(n_272), .B2(n_279), .C(n_282), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_267), .B(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_267), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g401 ( .A(n_267), .Y(n_401) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g379 ( .A(n_271), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_271), .B(n_319), .Y(n_395) );
INVx2_ASAP7_75t_L g381 ( .A(n_272), .Y(n_381) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_293), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_274), .A2(n_290), .B(n_332), .C(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_295), .Y(n_300) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_279), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g348 ( .A(n_280), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_285), .B2(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
INVx1_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
INVx1_ASAP7_75t_L g400 ( .A(n_288), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_297), .C(n_320), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g363 ( .A(n_293), .Y(n_363) );
AND2x2_ASAP7_75t_L g412 ( .A(n_293), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B(n_310), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g326 ( .A(n_300), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_300), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g394 ( .A(n_301), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_301), .A2(n_353), .A3(n_360), .B1(n_401), .B2(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_SL g373 ( .A(n_303), .Y(n_373) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g313 ( .A(n_309), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_312), .A2(n_360), .B1(n_386), .B2(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_316), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_339), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_385), .Y(n_380) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_364), .C(n_380), .D(n_390), .E(n_408), .Y(n_340) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_347), .C(n_354), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g411 ( .A(n_348), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_SL g387 ( .A(n_357), .Y(n_387) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g369 ( .A1(n_360), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_373), .C1(n_374), .C2(n_375), .Y(n_369) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_362), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_362), .B(n_387), .Y(n_386) );
AOI211xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_367), .B(n_369), .C(n_377), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_373), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_398), .B1(n_399), .B2(n_403), .C(n_405), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_395), .C(n_396), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g417 ( .A(n_393), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_408) );
AOI21xp33_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_417), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_427), .Y(n_434) );
BUFx2_ASAP7_75t_L g446 ( .A(n_427), .Y(n_446) );
INVx1_ASAP7_75t_SL g732 ( .A(n_427), .Y(n_732) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_428), .B(n_452), .Y(n_728) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_429), .A2(n_450), .B1(n_451), .B2(n_714), .C(n_723), .Y(n_449) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_440), .A2(n_441), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g730 ( .A(n_440), .B(n_442), .Y(n_730) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_724), .B(n_729), .Y(n_447) );
INVxp33_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
AO22x2_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_453), .B1(n_454), .B2(n_713), .Y(n_451) );
INVx1_ASAP7_75t_L g713 ( .A(n_452), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_455), .B(n_656), .Y(n_454) );
AND4x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_596), .C(n_611), .D(n_636), .Y(n_455) );
NOR2xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_569), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_487), .B(n_549), .Y(n_457) );
AND2x2_ASAP7_75t_L g599 ( .A(n_458), .B(n_504), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_458), .B(n_503), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_458), .B(n_488), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_458), .Y(n_666) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_475), .Y(n_458) );
INVx2_ASAP7_75t_L g583 ( .A(n_459), .Y(n_583) );
BUFx2_ASAP7_75t_L g610 ( .A(n_459), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_470), .Y(n_460) );
INVx5_ASAP7_75t_L g480 ( .A(n_462), .Y(n_480) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_469), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_469), .A2(n_480), .B(n_560), .C(n_561), .Y(n_559) );
BUFx2_ASAP7_75t_L g507 ( .A(n_471), .Y(n_507) );
AND2x2_ASAP7_75t_L g550 ( .A(n_475), .B(n_504), .Y(n_550) );
INVx2_ASAP7_75t_L g566 ( .A(n_475), .Y(n_566) );
AND2x2_ASAP7_75t_L g575 ( .A(n_475), .B(n_503), .Y(n_575) );
AND2x2_ASAP7_75t_L g654 ( .A(n_475), .B(n_583), .Y(n_654) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_486), .Y(n_475) );
INVx2_ASAP7_75t_L g494 ( .A(n_480), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_516), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_488), .B(n_581), .Y(n_619) );
INVx1_ASAP7_75t_L g707 ( .A(n_488), .Y(n_707) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_503), .Y(n_488) );
AND2x2_ASAP7_75t_L g565 ( .A(n_489), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g579 ( .A(n_489), .B(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_489), .Y(n_608) );
OR2x2_ASAP7_75t_L g640 ( .A(n_489), .B(n_582), .Y(n_640) );
AND2x2_ASAP7_75t_L g648 ( .A(n_489), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g681 ( .A(n_489), .B(n_650), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_489), .B(n_550), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_489), .B(n_610), .Y(n_706) );
AND2x2_ASAP7_75t_L g712 ( .A(n_489), .B(n_599), .Y(n_712) );
INVx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g572 ( .A(n_490), .Y(n_572) );
AND2x2_ASAP7_75t_L g602 ( .A(n_490), .B(n_582), .Y(n_602) );
AND2x2_ASAP7_75t_L g635 ( .A(n_490), .B(n_595), .Y(n_635) );
AND2x2_ASAP7_75t_L g655 ( .A(n_490), .B(n_504), .Y(n_655) );
AND2x2_ASAP7_75t_L g689 ( .A(n_490), .B(n_555), .Y(n_689) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_499), .C(n_500), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_497), .A2(n_500), .B(n_546), .C(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g595 ( .A(n_503), .B(n_566), .Y(n_595) );
AND2x2_ASAP7_75t_L g606 ( .A(n_503), .B(n_602), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_503), .B(n_582), .Y(n_645) );
INVx2_ASAP7_75t_L g660 ( .A(n_503), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_503), .B(n_594), .Y(n_683) );
AND2x2_ASAP7_75t_L g702 ( .A(n_503), .B(n_654), .Y(n_702) );
INVx5_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_504), .Y(n_601) );
AND2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g650 ( .A(n_504), .B(n_566), .Y(n_650) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
AOI21xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_508), .B(n_512), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
AND2x2_ASAP7_75t_L g573 ( .A(n_518), .B(n_556), .Y(n_573) );
INVx1_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_519), .B(n_530), .Y(n_553) );
OR2x2_ASAP7_75t_L g586 ( .A(n_519), .B(n_556), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_519), .B(n_556), .Y(n_591) );
AND2x2_ASAP7_75t_L g618 ( .A(n_519), .B(n_555), .Y(n_618) );
AND2x2_ASAP7_75t_L g670 ( .A(n_519), .B(n_529), .Y(n_670) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_520), .B(n_540), .Y(n_578) );
AND2x2_ASAP7_75t_L g614 ( .A(n_520), .B(n_530), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_527), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g604 ( .A(n_528), .B(n_586), .Y(n_604) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
OAI322xp33_ASAP7_75t_L g569 ( .A1(n_529), .A2(n_570), .A3(n_574), .B1(n_576), .B2(n_579), .C1(n_584), .C2(n_592), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_529), .B(n_555), .Y(n_577) );
OR2x2_ASAP7_75t_L g587 ( .A(n_529), .B(n_541), .Y(n_587) );
AND2x2_ASAP7_75t_L g589 ( .A(n_529), .B(n_541), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_529), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_529), .B(n_556), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_529), .B(n_685), .Y(n_684) );
INVx5_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_530), .B(n_573), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_540), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g567 ( .A(n_540), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_540), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g629 ( .A(n_540), .B(n_556), .Y(n_629) );
AOI211xp5_ASAP7_75t_SL g657 ( .A1(n_540), .A2(n_658), .B(n_661), .C(n_673), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_540), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g695 ( .A(n_540), .B(n_670), .Y(n_695) );
INVx5_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g623 ( .A(n_541), .B(n_556), .Y(n_623) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_541), .Y(n_632) );
AND2x2_ASAP7_75t_L g672 ( .A(n_541), .B(n_670), .Y(n_672) );
AND2x2_ASAP7_75t_SL g703 ( .A(n_541), .B(n_573), .Y(n_703) );
AND2x2_ASAP7_75t_L g710 ( .A(n_541), .B(n_669), .Y(n_710) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_565), .B2(n_567), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_550), .B(n_572), .Y(n_620) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g568 ( .A(n_553), .Y(n_568) );
OR2x2_ASAP7_75t_L g628 ( .A(n_553), .B(n_629), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_553), .A2(n_677), .B1(n_679), .B2(n_680), .C(n_682), .Y(n_676) );
INVx2_ASAP7_75t_L g615 ( .A(n_554), .Y(n_615) );
AND2x2_ASAP7_75t_L g588 ( .A(n_555), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g678 ( .A(n_555), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_555), .B(n_670), .Y(n_691) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVxp67_ASAP7_75t_L g633 ( .A(n_556), .Y(n_633) );
AND2x2_ASAP7_75t_L g669 ( .A(n_556), .B(n_670), .Y(n_669) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_564), .Y(n_556) );
AND2x2_ASAP7_75t_L g671 ( .A(n_565), .B(n_610), .Y(n_671) );
AND2x2_ASAP7_75t_L g581 ( .A(n_566), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_566), .B(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g652 ( .A(n_568), .B(n_615), .Y(n_652) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g658 ( .A(n_571), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OR2x2_ASAP7_75t_L g644 ( .A(n_572), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g709 ( .A(n_572), .B(n_654), .Y(n_709) );
INVx2_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
NAND4xp25_ASAP7_75t_SL g705 ( .A(n_574), .B(n_706), .C(n_707), .D(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_575), .B(n_639), .Y(n_674) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g711 ( .A(n_578), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_SL g673 ( .A1(n_579), .A2(n_642), .B(n_646), .C(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g668 ( .A(n_581), .B(n_660), .Y(n_668) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_582), .Y(n_594) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B(n_588), .C(n_590), .Y(n_584) );
AND2x2_ASAP7_75t_L g605 ( .A(n_585), .B(n_589), .Y(n_605) );
OAI322xp33_ASAP7_75t_SL g643 ( .A1(n_585), .A2(n_644), .A3(n_646), .B1(n_647), .B2(n_651), .C1(n_652), .C2(n_653), .Y(n_643) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g665 ( .A(n_587), .B(n_591), .Y(n_665) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
INVx1_ASAP7_75t_SL g664 ( .A(n_591), .Y(n_664) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_603), .B1(n_605), .B2(n_606), .C1(n_607), .C2(n_734), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
OAI322xp33_ASAP7_75t_L g686 ( .A1(n_598), .A2(n_660), .A3(n_665), .B1(n_687), .B2(n_688), .C1(n_690), .C2(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_599), .A2(n_613), .B1(n_637), .B2(n_641), .C(n_643), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OAI222xp33_ASAP7_75t_L g616 ( .A1(n_604), .A2(n_617), .B1(n_619), .B2(n_620), .C1(n_621), .C2(n_624), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_606), .A2(n_613), .B1(n_683), .B2(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_616), .C(n_627), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_613), .A2(n_650), .B(n_693), .C(n_696), .Y(n_692) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g622 ( .A(n_614), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g685 ( .A(n_618), .Y(n_685) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_625), .B(n_650), .Y(n_679) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_634), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g696 ( .A1(n_628), .A2(n_697), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_696) );
INVxp33_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_632), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_639), .B(n_650), .Y(n_690) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
AND2x2_ASAP7_75t_L g701 ( .A(n_654), .B(n_660), .Y(n_701) );
AND4x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_675), .C(n_692), .D(n_704), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI221xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g697 ( .A(n_668), .Y(n_697) );
INVx1_ASAP7_75t_SL g687 ( .A(n_672), .Y(n_687) );
NOR2xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_686), .Y(n_675) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_688), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_695), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g723 ( .A(n_714), .Y(n_723) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
INVxp33_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx3_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NAND2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
endmodule