module fake_jpeg_19818_n_263 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_23),
.B1(n_13),
.B2(n_17),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_22),
.B1(n_29),
.B2(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_56),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_25),
.A3(n_27),
.B1(n_24),
.B2(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_39),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_53),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_73),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_56),
.Y(n_88)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_57),
.B(n_47),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_85),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_86),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_56),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_35),
.C(n_52),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_26),
.C(n_28),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_35),
.B1(n_56),
.B2(n_41),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_92),
.B1(n_60),
.B2(n_28),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_46),
.B1(n_45),
.B2(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_73),
.B1(n_69),
.B2(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_78),
.B1(n_82),
.B2(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_63),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_90),
.B(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_103),
.B1(n_94),
.B2(n_95),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_26),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_76),
.B1(n_63),
.B2(n_51),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_76),
.B(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_109),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_62),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_83),
.B1(n_79),
.B2(n_88),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_28),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_116),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_78),
.B(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_134),
.B(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_133),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_131),
.B(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_140),
.B1(n_55),
.B2(n_37),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_92),
.B1(n_87),
.B2(n_86),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_72),
.B1(n_26),
.B2(n_64),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_59),
.B(n_77),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_59),
.B(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_66),
.B(n_1),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_102),
.C(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_72),
.C(n_43),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_20),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_22),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_111),
.B1(n_110),
.B2(n_72),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_21),
.B(n_20),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_64),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_147),
.C(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_136),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_165),
.Y(n_168)
);

INVxp33_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_70),
.B1(n_66),
.B2(n_58),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_133),
.B1(n_119),
.B2(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_139),
.B1(n_134),
.B2(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_166),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_70),
.B1(n_66),
.B2(n_58),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_70),
.B1(n_32),
.B2(n_31),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_16),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_22),
.B1(n_12),
.B2(n_18),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_32),
.C(n_31),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_125),
.B(n_120),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_175),
.B(n_12),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_128),
.B(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_174),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_117),
.B(n_15),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_15),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_156),
.B1(n_151),
.B2(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_164),
.B1(n_158),
.B2(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_186),
.B1(n_179),
.B2(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_159),
.B1(n_163),
.B2(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_166),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_172),
.Y(n_211)
);

OAI21x1_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_176),
.B(n_182),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_31),
.C(n_30),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_32),
.C(n_30),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_191),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_210),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_171),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_212),
.C(n_173),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_216),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_169),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_173),
.C(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_177),
.C(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_190),
.B1(n_189),
.B2(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_183),
.C(n_173),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_174),
.C(n_30),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_227),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_16),
.C(n_1),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_16),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_5),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_207),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_205),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_5),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_235),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_6),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_7),
.B(n_2),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_4),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_228),
.B(n_1),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_240),
.A2(n_244),
.B(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_7),
.B(n_2),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_7),
.C(n_2),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_3),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_3),
.C(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_3),
.B(n_4),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_242),
.B(n_241),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_255),
.B(n_10),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_4),
.B(n_7),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_248),
.B(n_8),
.C(n_9),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_9),
.B1(n_10),
.B2(n_0),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_9),
.C(n_0),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_261),
.B(n_9),
.CI(n_0),
.CON(n_262),
.SN(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);


endmodule