module real_jpeg_15238_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_104),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_0),
.A2(n_104),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_0),
.A2(n_104),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_1),
.A2(n_101),
.B1(n_304),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_1),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_1),
.A2(n_307),
.B1(n_436),
.B2(n_439),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_1),
.A2(n_307),
.B1(n_497),
.B2(n_499),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_89),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_2),
.A2(n_89),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_2),
.A2(n_89),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_545),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_3),
.B(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

OAI22x1_ASAP7_75t_L g266 ( 
.A1(n_6),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_6),
.A2(n_270),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

OAI22x1_ASAP7_75t_SL g467 ( 
.A1(n_6),
.A2(n_270),
.B1(n_468),
.B2(n_470),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_6),
.A2(n_270),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_7),
.A2(n_36),
.B1(n_122),
.B2(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_7),
.A2(n_125),
.B1(n_283),
.B2(n_287),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_7),
.A2(n_125),
.B1(n_423),
.B2(n_425),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_7),
.A2(n_125),
.B1(n_381),
.B2(n_503),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_9),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_10),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_10),
.Y(n_438)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_11),
.B(n_87),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_11),
.A2(n_45),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_11),
.A2(n_241),
.A3(n_246),
.B1(n_247),
.B2(n_250),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_11),
.B(n_293),
.Y(n_292)
);

OAI32xp33_ASAP7_75t_L g340 ( 
.A1(n_11),
.A2(n_341),
.A3(n_345),
.B1(n_350),
.B2(n_354),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_11),
.A2(n_45),
.B1(n_373),
.B2(n_376),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_L g429 ( 
.A1(n_11),
.A2(n_341),
.A3(n_345),
.B1(n_350),
.B2(n_354),
.Y(n_429)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_12),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_12),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_12),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_13),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_14),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_14),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_130),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_14),
.A2(n_130),
.B1(n_311),
.B2(n_317),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_14),
.A2(n_130),
.B1(n_356),
.B2(n_415),
.Y(n_414)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_16),
.A2(n_331),
.B1(n_335),
.B2(n_339),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_16),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_16),
.A2(n_339),
.B1(n_452),
.B2(n_454),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_16),
.A2(n_339),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_17),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_17),
.Y(n_357)
);

BUFx8_ASAP7_75t_L g382 ( 
.A(n_17),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_17),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_514),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_481),
.B(n_511),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_404),
.B(n_478),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_321),
.B(n_403),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_274),
.B(n_320),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_196),
.B(n_273),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_145),
.B(n_195),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_97),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_29),
.B(n_97),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_60),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_30),
.A2(n_60),
.B1(n_61),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_30),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.A3(n_40),
.B1(n_44),
.B2(n_50),
.Y(n_30)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_39),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_45),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_45),
.A2(n_108),
.B1(n_166),
.B2(n_171),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_45),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_45),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_87),
.B2(n_88),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_87),
.B1(n_88),
.B2(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_67),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_67),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_67),
.B(n_396),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_70),
.Y(n_286)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_70),
.Y(n_442)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_70),
.Y(n_453)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_71),
.Y(n_399)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_78),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_78),
.B(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_78),
.A2(n_201),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_80),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_80),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_84),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_87),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_87),
.B(n_435),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_95),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_126),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_98),
.B(n_127),
.C(n_133),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_108),
.B(n_115),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_108),
.A2(n_149),
.B1(n_171),
.B2(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_108),
.B(n_266),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_108),
.A2(n_121),
.B(n_488),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_111),
.Y(n_488)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_116),
.B(n_308),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_121),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_134),
.B(n_467),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_134),
.A2(n_419),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

AO22x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_134)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_135),
.Y(n_454)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_141),
.Y(n_222)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_163),
.B(n_194),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_161),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_161),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_154),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_154),
.A2(n_157),
.B1(n_303),
.B2(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_154),
.A2(n_261),
.B(n_330),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_187),
.B(n_193),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_179),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_175),
.Y(n_269)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_175),
.Y(n_334)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_197),
.B(n_198),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_239),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_211),
.C(n_239),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_201),
.A2(n_282),
.B(n_395),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_201),
.A2(n_395),
.B(n_451),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_227),
.B1(n_233),
.B2(n_238),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_212),
.A2(n_233),
.B1(n_238),
.B2(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_212),
.A2(n_238),
.B1(n_310),
.B2(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_212),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_212),
.A2(n_422),
.B(n_466),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_212),
.A2(n_238),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_222),
.B2(n_223),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_218),
.Y(n_527)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_220),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_221),
.Y(n_316)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_226),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_226),
.Y(n_469)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_228),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_230),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g421 ( 
.A(n_238),
.B(n_422),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_259),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_259),
.Y(n_278)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_244),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_245),
.Y(n_393)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_254),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_255),
.Y(n_344)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_275),
.B(n_276),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_288),
.B1(n_289),
.B2(n_319),
.Y(n_276)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

XOR2x1_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_279),
.C(n_288),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_281),
.B(n_529),
.Y(n_528)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_309),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_299),
.B2(n_300),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_300),
.C(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OR2x6_ASAP7_75t_L g363 ( 
.A(n_293),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_293),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_293),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_293),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_293),
.B(n_536),
.Y(n_535)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g366 ( 
.A(n_295),
.Y(n_366)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_296),
.Y(n_427)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_318),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_323),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_361),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_326),
.B(n_327),
.C(n_361),
.Y(n_475)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_340),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_329),
.B(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_356),
.A2(n_365),
.B1(n_367),
.B2(n_369),
.Y(n_364)
);

INVx8_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_357),
.Y(n_539)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_384),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_385),
.C(n_394),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_372),
.B1(n_379),
.B2(n_383),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_363),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_363),
.A2(n_383),
.B1(n_414),
.B2(n_460),
.Y(n_459)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_363),
.A2(n_460),
.B(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_363),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_378),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

BUFx12f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_394),
.Y(n_384)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_474),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_444),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_407),
.B(n_444),
.C(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_430),
.C(n_431),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_408),
.B(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_428),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_418),
.C(n_428),
.Y(n_445)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B(n_421),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_431),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_433),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_443),
.Y(n_433)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_455),
.C(n_473),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_455),
.B1(n_456),
.B2(n_473),
.Y(n_446)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_449),
.Y(n_505)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_456),
.Y(n_455)
);

XOR2x2_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_508),
.C(n_509),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_465),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_459),
.Y(n_508)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_476),
.Y(n_480)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_484),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_485),
.A2(n_506),
.B1(n_507),
.B2(n_510),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_485),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_492),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_486),
.B(n_492),
.C(n_506),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_487),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_487),
.A2(n_491),
.B1(n_533),
.B2(n_540),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_490),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_505),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_500),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_494),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_519),
.C(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_544),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_517),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_531),
.B1(n_542),
.B2(n_543),
.Y(n_521)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_522),
.Y(n_543)
);

OAI21xp33_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_528),
.B(n_530),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_528),
.Y(n_530)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_541),
.Y(n_531)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);


endmodule