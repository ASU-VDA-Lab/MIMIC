module fake_jpeg_2251_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_52),
.Y(n_95)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_48),
.B(n_49),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_51),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_2),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_58),
.C(n_76),
.Y(n_129)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g136 ( 
.A(n_57),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_2),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_62),
.Y(n_103)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_3),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_4),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_5),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_31),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_82),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_35),
.B(n_5),
.Y(n_82)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_33),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_31),
.B1(n_24),
.B2(n_38),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_91),
.A2(n_102),
.B1(n_117),
.B2(n_108),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_96),
.B(n_98),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_37),
.B1(n_22),
.B2(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_104),
.B1(n_117),
.B2(n_119),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_28),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_31),
.B1(n_24),
.B2(n_38),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_64),
.B1(n_66),
.B2(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_113),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_28),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_98),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_52),
.B(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_116),
.B(n_132),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_22),
.B1(n_36),
.B2(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_28),
.B1(n_35),
.B2(n_33),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_124),
.B1(n_109),
.B2(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_39),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_9),
.C(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_73),
.B(n_87),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_10),
.B(n_129),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_169),
.B(n_175),
.C(n_92),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_89),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_147),
.B(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_94),
.A2(n_104),
.B1(n_120),
.B2(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_161),
.B1(n_170),
.B2(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_131),
.Y(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_166),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_103),
.B(n_90),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_160),
.Y(n_188)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_120),
.B1(n_100),
.B2(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_163),
.Y(n_189)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_114),
.B(n_96),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_118),
.B(n_88),
.C(n_107),
.Y(n_169)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_173),
.Y(n_204)
);

BUFx4f_ASAP7_75t_SL g173 ( 
.A(n_88),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_173),
.Y(n_197)
);

OR2x4_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_109),
.Y(n_175)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_179),
.Y(n_207)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_192),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_92),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_92),
.B1(n_175),
.B2(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_180),
.B1(n_181),
.B2(n_188),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_143),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_160),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_150),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_205),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_177),
.B1(n_179),
.B2(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_172),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_218),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_169),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_221),
.C(n_227),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_158),
.B(n_176),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_186),
.B(n_195),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_153),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_195),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_235),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_192),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_189),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_189),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_198),
.B1(n_194),
.B2(n_207),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_226),
.B1(n_236),
.B2(n_253),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_206),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_249),
.C(n_231),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_182),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_196),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_251),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_196),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_223),
.C(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_235),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_221),
.C(n_223),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_263),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_215),
.B1(n_224),
.B2(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_219),
.C(n_217),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_214),
.Y(n_264)
);

BUFx12f_ASAP7_75t_SL g279 ( 
.A(n_264),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_265),
.A2(n_244),
.B1(n_236),
.B2(n_248),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_220),
.B(n_218),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_241),
.B(n_252),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_245),
.B(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_272),
.B1(n_278),
.B2(n_256),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_262),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_280),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_258),
.C(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_224),
.B1(n_216),
.B2(n_182),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_211),
.B(n_200),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_282),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_274),
.C(n_276),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_271),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_266),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_270),
.B1(n_272),
.B2(n_278),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_262),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_268),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_279),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.C(n_294),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_296),
.B(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_292),
.C(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_269),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_301),
.C(n_280),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_305),
.B(n_259),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_211),
.Y(n_308)
);


endmodule