module real_jpeg_33369_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g383 ( 
.A(n_0),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_83),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_83),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_1),
.A2(n_36),
.B1(n_83),
.B2(n_257),
.Y(n_256)
);

CKINVDCx11_ASAP7_75t_R g472 ( 
.A(n_2),
.Y(n_472)
);

CKINVDCx11_ASAP7_75t_R g482 ( 
.A(n_2),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_3),
.B(n_472),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_6),
.Y(n_196)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_48),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_48),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_7),
.A2(n_48),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_7),
.B(n_306),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_7),
.A2(n_322),
.A3(n_324),
.B1(n_326),
.B2(n_332),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_7),
.B(n_94),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_7),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_7),
.B(n_160),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_8),
.Y(n_337)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_11),
.A2(n_108),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_108),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_11),
.A2(n_108),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_36),
.B1(n_39),
.B2(n_43),
.Y(n_35)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_13),
.A2(n_43),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_13),
.A2(n_43),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_470),
.B(n_481),
.Y(n_14)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_15),
.A2(n_471),
.B(n_474),
.C(n_482),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_259),
.B(n_464),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_236),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_203),
.Y(n_17)
);

OAI21x1_ASAP7_75t_SL g465 ( 
.A1(n_18),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_145),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_19),
.B(n_145),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_20),
.B(n_21),
.C(n_127),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.C(n_91),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_21),
.A2(n_22),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_22),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_24),
.B(n_210),
.C(n_266),
.Y(n_428)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g420 ( 
.A1(n_25),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_25),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_44),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_26),
.A2(n_35),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_26),
.B(n_132),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_244),
.B(n_250),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_26),
.A2(n_132),
.B1(n_244),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_52),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_27),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_43),
.A2(n_142),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_43),
.B(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_44),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_45),
.B(n_202),
.Y(n_201)
);

OAI21x1_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_48),
.B(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_48),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_48),
.B(n_370),
.Y(n_369)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_49),
.A2(n_245),
.A3(n_273),
.B1(n_277),
.B2(n_280),
.Y(n_272)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_56),
.Y(n_282)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_59),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_60),
.A2(n_61),
.B1(n_91),
.B2(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_61),
.B(n_129),
.C(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_82),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_62),
.B(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_74),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_74),
.Y(n_63)
);

NAND2x1p5_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_74),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_66),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_66),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_66),
.Y(n_373)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_69),
.Y(n_368)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_74),
.B(n_226),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_76),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_79),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_80),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_82),
.A2(n_152),
.B1(n_158),
.B2(n_160),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_85),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_96),
.B1(n_99),
.B2(n_103),
.Y(n_95)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_89),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_105),
.B(n_112),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_105),
.B1(n_136),
.B2(n_144),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_93),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_R g242 ( 
.A(n_93),
.B(n_144),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_93),
.A2(n_144),
.B(n_162),
.Y(n_422)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_94),
.B(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_113),
.B(n_117),
.Y(n_212)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_123),
.Y(n_331)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_125),
.Y(n_284)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_129),
.B(n_210),
.C(n_213),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_129),
.B(n_161),
.C(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g426 ( 
.A1(n_130),
.A2(n_131),
.B1(n_161),
.B2(n_303),
.Y(n_426)
);

AOI22x1_ASAP7_75t_L g445 ( 
.A1(n_130),
.A2(n_131),
.B1(n_210),
.B2(n_267),
.Y(n_445)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_139),
.Y(n_323)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_168),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_150),
.A2(n_151),
.B(n_161),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_160),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_160),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_161),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_161),
.A2(n_303),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_205),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_179),
.B(n_200),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_234),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_178),
.B(n_179),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_170),
.B(n_178),
.Y(n_442)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_172),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_200),
.B1(n_201),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_179),
.A2(n_235),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_187),
.Y(n_288)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_188),
.B(n_295),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_190),
.A2(n_286),
.B1(n_292),
.B2(n_295),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_190),
.B(n_295),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_194),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_202),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_204),
.B(n_207),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_231),
.C(n_232),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_209),
.B(n_231),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_210),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_265)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_210),
.A2(n_267),
.B1(n_345),
.B2(n_347),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_213),
.B(n_445),
.Y(n_444)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g413 ( 
.A1(n_214),
.A2(n_319),
.B1(n_398),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_214),
.Y(n_414)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_218),
.A2(n_312),
.B(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_223),
.B(n_350),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_223),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_233),
.B(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_253),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_237),
.A2(n_253),
.B(n_465),
.C(n_468),
.D(n_469),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_238),
.B(n_239),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_239),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.CI(n_251),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_243),
.C(n_251),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_R g469 ( 
.A(n_254),
.B(n_258),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_254),
.B(n_476),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_254),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_256),
.B(n_478),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_456),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_405),
.B(n_455),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_339),
.B(n_404),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_313),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_263),
.B(n_313),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_264),
.B(n_271),
.C(n_302),
.Y(n_430)
);

XNOR2x1_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_267),
.B(n_392),
.C(n_402),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_269),
.B(n_437),
.C(n_438),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_269),
.B(n_437),
.C(n_438),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_302),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_285),
.B1(n_300),
.B2(n_301),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_272),
.B(n_301),
.Y(n_411)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_285),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_285),
.B(n_385),
.Y(n_386)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx4f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_301),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.C(n_307),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_354),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_307),
.B(n_354),
.Y(n_387)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_308),
.B(n_379),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_311),
.B(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_318),
.C(n_320),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_314),
.A2(n_315),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_349),
.C(n_350),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_319),
.A2(n_320),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_338),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_321),
.B(n_338),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx4f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_395),
.B(n_403),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_351),
.B(n_394),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_348),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_348),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_355),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_417),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_345),
.B(n_417),
.Y(n_427)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_388),
.B(n_393),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_377),
.B(n_387),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_361),
.B1(n_369),
.B2(n_374),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_374),
.B(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_384),
.B(n_386),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_391),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_401),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_397),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_433),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_429),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_424),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_424),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_453),
.C(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_420),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_427),
.C(n_428),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_428),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_431),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_448),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_434),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_446),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_446),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_439),
.C(n_443),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_444),
.Y(n_451)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_452),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_463),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B(n_461),
.C(n_462),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_480),
.Y(n_479)
);


endmodule