module fake_jpeg_4604_n_214 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_6),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_6),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_59),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_73),
.B1(n_81),
.B2(n_84),
.Y(n_105)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_62),
.Y(n_98)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_71),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_25),
.B(n_24),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_14),
.B1(n_27),
.B2(n_4),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_14),
.B1(n_31),
.B2(n_16),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_24),
.B(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_19),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_85),
.Y(n_87)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_60),
.Y(n_99)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_95),
.B(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_11),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_25),
.B(n_14),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_58),
.B(n_53),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_37),
.B1(n_14),
.B2(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_102),
.B1(n_62),
.B2(n_49),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_2),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_49),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_8),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_11),
.C(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_113),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_89),
.B(n_109),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_131),
.B1(n_102),
.B2(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_93),
.B1(n_94),
.B2(n_91),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_132),
.B1(n_104),
.B2(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_87),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_54),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_64),
.B1(n_50),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_87),
.B(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_13),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_123),
.B1(n_126),
.B2(n_116),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_90),
.B1(n_95),
.B2(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_140),
.B1(n_153),
.B2(n_141),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_149),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_136),
.B(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_157),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_154),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_107),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_122),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_93),
.B1(n_103),
.B2(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_164),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_114),
.B1(n_125),
.B2(n_121),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_165),
.B1(n_170),
.B2(n_93),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_121),
.B(n_113),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_127),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_114),
.B1(n_118),
.B2(n_132),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_138),
.C(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_119),
.B(n_136),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_171),
.B(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_137),
.B(n_154),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_137),
.B1(n_152),
.B2(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_167),
.C(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_146),
.B1(n_145),
.B2(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_174),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_188),
.B1(n_169),
.B2(n_182),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_165),
.B1(n_161),
.B2(n_170),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_166),
.B(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_199),
.B(n_189),
.Y(n_204)
);

OAI211xp5_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_194),
.B(n_188),
.C(n_166),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_181),
.B1(n_179),
.B2(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_173),
.B(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_186),
.C(n_190),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_179),
.B(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_103),
.C(n_106),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_202),
.B(n_106),
.C(n_108),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_193),
.B1(n_189),
.B2(n_143),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_163),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_124),
.B(n_88),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.C(n_203),
.Y(n_209)
);

AOI31xp33_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_210),
.A3(n_108),
.B(n_13),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_91),
.C(n_96),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_96),
.B(n_108),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);


endmodule