module fake_jpeg_22849_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_21),
.B(n_34),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_18),
.B(n_31),
.C(n_30),
.Y(n_76)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_26),
.B1(n_34),
.B2(n_19),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_67),
.B(n_76),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_70),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_34),
.B1(n_38),
.B2(n_20),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_45),
.B1(n_41),
.B2(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_34),
.B1(n_38),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_38),
.B1(n_20),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_32),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_87),
.B1(n_88),
.B2(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_44),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_24),
.B1(n_37),
.B2(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_37),
.B1(n_31),
.B2(n_30),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_92),
.B(n_116),
.Y(n_135)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_94),
.A2(n_84),
.B1(n_52),
.B2(n_51),
.Y(n_140)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_105),
.B1(n_93),
.B2(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_49),
.C(n_44),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_50),
.B(n_83),
.Y(n_128)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_28),
.B1(n_30),
.B2(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_43),
.Y(n_152)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_60),
.B(n_1),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_82),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_150),
.B1(n_69),
.B2(n_73),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_68),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_146),
.C(n_109),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_138),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_117),
.B(n_103),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_142),
.B(n_143),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_88),
.C(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_51),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_153),
.B1(n_108),
.B2(n_73),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_49),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_18),
.C(n_73),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_50),
.B(n_52),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_49),
.B(n_18),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_44),
.B(n_43),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_119),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_43),
.B1(n_41),
.B2(n_57),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_111),
.B1(n_108),
.B2(n_118),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_97),
.A2(n_43),
.B1(n_69),
.B2(n_57),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_116),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_166),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_91),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_128),
.B(n_137),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_91),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_176),
.B(n_178),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_164),
.B1(n_139),
.B2(n_123),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_184),
.B1(n_151),
.B2(n_148),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_170),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_177),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_120),
.C(n_101),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_182),
.C(n_129),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_101),
.B(n_95),
.C(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_95),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_18),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_170),
.B1(n_136),
.B2(n_122),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_69),
.B1(n_119),
.B2(n_17),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_187),
.B(n_194),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_198),
.C(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_136),
.A3(n_16),
.B1(n_126),
.B2(n_134),
.C1(n_7),
.C2(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_126),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_148),
.B1(n_151),
.B2(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_164),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_194),
.B(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_217),
.B1(n_226),
.B2(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_227),
.B1(n_228),
.B2(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_167),
.Y(n_219)
);

FAx1_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_154),
.CI(n_157),
.CON(n_236),
.SN(n_236)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_179),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_220),
.Y(n_234)
);

OAI321xp33_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_170),
.A3(n_186),
.B1(n_206),
.B2(n_196),
.C(n_183),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_162),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_177),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_188),
.C(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_157),
.C(n_187),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_155),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_166),
.B(n_161),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_239),
.C(n_240),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_156),
.B1(n_185),
.B2(n_181),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_237),
.B1(n_242),
.B2(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_225),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_211),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_219),
.B(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_200),
.B1(n_176),
.B2(n_204),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_238),
.B(n_219),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_203),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_202),
.B1(n_208),
.B2(n_159),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_159),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_215),
.C(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_231),
.B1(n_236),
.B2(n_241),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_228),
.B(n_221),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_6),
.B(n_9),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_225),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_257),
.B1(n_258),
.B2(n_6),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_256),
.C(n_240),
.Y(n_259)
);

XOR2x1_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_209),
.C(n_226),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_209),
.B1(n_224),
.B2(n_16),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_267),
.B1(n_268),
.B2(n_6),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_234),
.C(n_7),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_257),
.Y(n_270)
);

OAI21x1_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_10),
.B(n_11),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_248),
.B1(n_246),
.B2(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_259),
.B1(n_247),
.B2(n_266),
.Y(n_276)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_255),
.B1(n_249),
.B2(n_247),
.C(n_250),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_10),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_10),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.C(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_266),
.C(n_262),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_275),
.B(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_270),
.Y(n_286)
);

OAI321xp33_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_287),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_285),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_279),
.B(n_271),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_13),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_14),
.Y(n_290)
);


endmodule