module fake_jpeg_7103_n_80 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_2),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_55),
.B1(n_45),
.B2(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_4),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_61),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_39),
.B(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_57),
.C(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_35),
.B1(n_38),
.B2(n_8),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_70),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B(n_7),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_44),
.C(n_12),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_72),
.B1(n_62),
.B2(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_13),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_16),
.B(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_33),
.B1(n_22),
.B2(n_23),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_27),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_28),
.Y(n_80)
);


endmodule