module fake_jpeg_28890_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx8_ASAP7_75t_SL g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_17),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_57),
.C(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_45),
.B1(n_58),
.B2(n_3),
.Y(n_69)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_65),
.Y(n_68)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_75),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_44),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_52),
.B1(n_46),
.B2(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_52),
.B1(n_53),
.B2(n_48),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_50),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_0),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_8),
.C(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_99)
);

OAI211xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_23),
.B(n_43),
.C(n_42),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_79),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_50),
.B(n_19),
.C(n_20),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_13),
.B(n_30),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_89),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_4),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_110),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_6),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_8),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_24),
.B1(n_40),
.B2(n_39),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_15),
.B(n_38),
.Y(n_114)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_120),
.B(n_122),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_14),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_107),
.C(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_123),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_16),
.B(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_127),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_112),
.A2(n_101),
.B1(n_111),
.B2(n_105),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_98),
.C(n_33),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_9),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_122),
.B(n_115),
.C(n_117),
.D(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_134),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_126),
.B1(n_117),
.B2(n_125),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_128),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_135),
.B(n_136),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_132),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_41),
.B(n_10),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_10),
.Y(n_142)
);


endmodule