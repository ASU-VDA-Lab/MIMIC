module fake_jpeg_2578_n_613 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_613);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_58),
.B(n_88),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_11),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_61),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_66),
.Y(n_160)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_33),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_76),
.B(n_78),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_10),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_79),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_10),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_93),
.Y(n_171)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_29),
.B(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_10),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_96),
.Y(n_209)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_113),
.Y(n_186)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_35),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx12f_ASAP7_75t_SL g200 ( 
.A(n_126),
.Y(n_200)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_57),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_131),
.A2(n_185),
.B(n_187),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_56),
.B(n_52),
.C(n_53),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_134),
.B(n_177),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_90),
.B(n_56),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_140),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_82),
.B1(n_120),
.B2(n_83),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_139),
.A2(n_154),
.B1(n_170),
.B2(n_137),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_69),
.B(n_85),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_30),
.B1(n_46),
.B2(n_45),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_142),
.A2(n_166),
.B1(n_192),
.B2(n_214),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_150),
.B(n_158),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_63),
.A2(n_57),
.B1(n_53),
.B2(n_51),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_152),
.A2(n_181),
.B1(n_49),
.B2(n_32),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_59),
.A2(n_57),
.B1(n_53),
.B2(n_51),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_86),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_43),
.B1(n_38),
.B2(n_46),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_106),
.A2(n_51),
.B1(n_50),
.B2(n_45),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_71),
.B(n_44),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_50),
.B1(n_44),
.B2(n_43),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_96),
.A2(n_29),
.B1(n_39),
.B2(n_38),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_103),
.B(n_50),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_77),
.B(n_39),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_210),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_79),
.A2(n_35),
.B1(n_49),
.B2(n_32),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_111),
.B(n_114),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_0),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_80),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_116),
.B(n_15),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_87),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_95),
.A2(n_35),
.B1(n_49),
.B2(n_32),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_119),
.B(n_15),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_136),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

BUFx2_ASAP7_75t_SL g315 ( 
.A(n_222),
.Y(n_315)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_170),
.B1(n_201),
.B2(n_206),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_128),
.B1(n_124),
.B2(n_35),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_225),
.A2(n_214),
.B1(n_210),
.B2(n_130),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_227),
.B(n_228),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_186),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_136),
.A2(n_171),
.B(n_169),
.C(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_229),
.B(n_231),
.Y(n_310)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_233),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_163),
.A2(n_35),
.B1(n_49),
.B2(n_32),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_234),
.A2(n_258),
.B1(n_271),
.B2(n_285),
.Y(n_319)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_236),
.A2(n_241),
.B1(n_249),
.B2(n_289),
.Y(n_327)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_137),
.Y(n_237)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_238),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_246),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_171),
.A2(n_49),
.B1(n_32),
.B2(n_26),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_161),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_244),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_12),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_247),
.Y(n_336)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_181),
.A2(n_26),
.B1(n_13),
.B2(n_4),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_252),
.Y(n_351)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_148),
.Y(n_253)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_255),
.B(n_265),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_161),
.Y(n_256)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_7),
.B1(n_17),
.B2(n_4),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_132),
.Y(n_259)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_259),
.Y(n_324)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_146),
.Y(n_261)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_267),
.Y(n_317)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_143),
.B(n_7),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_270),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_140),
.Y(n_270)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_272),
.B(n_275),
.Y(n_335)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_174),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_273),
.B(n_274),
.Y(n_353)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_149),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_165),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_167),
.B(n_198),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_279),
.Y(n_340)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_277),
.B(n_278),
.Y(n_357)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_146),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_280),
.Y(n_326)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_282),
.Y(n_337)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_283),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_7),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_293),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_147),
.A2(n_7),
.B1(n_17),
.B2(n_4),
.Y(n_285)
);

INVx3_ASAP7_75t_SL g286 ( 
.A(n_129),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_286),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_153),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_332)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_180),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_15),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_300),
.B1(n_204),
.B2(n_213),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_133),
.B(n_5),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_184),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_296),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_154),
.A2(n_5),
.B1(n_6),
.B2(n_16),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_295),
.A2(n_151),
.B1(n_162),
.B2(n_203),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_159),
.Y(n_296)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_196),
.Y(n_338)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_162),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_226),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_316),
.C(n_333),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_313),
.A2(n_338),
.B1(n_337),
.B2(n_344),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_135),
.B1(n_141),
.B2(n_194),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_314),
.A2(n_322),
.B1(n_343),
.B2(n_261),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_193),
.C(n_195),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_223),
.A2(n_212),
.B1(n_179),
.B2(n_144),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

OAI22x1_ASAP7_75t_L g328 ( 
.A1(n_224),
.A2(n_191),
.B1(n_188),
.B2(n_205),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_328),
.A2(n_292),
.B1(n_290),
.B2(n_256),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_243),
.B(n_272),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_338),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_255),
.B(n_212),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_286),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_225),
.A2(n_179),
.B1(n_144),
.B2(n_213),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_268),
.A2(n_151),
.B(n_16),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_354),
.B(n_237),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_352),
.A2(n_356),
.B1(n_323),
.B2(n_327),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_230),
.A2(n_16),
.B(n_17),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_289),
.A2(n_262),
.B1(n_203),
.B2(n_232),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_327),
.A2(n_234),
.B1(n_291),
.B2(n_285),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_359),
.A2(n_388),
.B1(n_392),
.B2(n_325),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_341),
.A2(n_252),
.B1(n_299),
.B2(n_248),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_360),
.A2(n_377),
.B1(n_378),
.B2(n_387),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_298),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_361),
.B(n_362),
.C(n_380),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_245),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_310),
.A2(n_258),
.B(n_239),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_364),
.A2(n_373),
.B(n_376),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_306),
.B(n_296),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_366),
.B(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_372),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_265),
.A3(n_274),
.B1(n_278),
.B2(n_277),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_322),
.A2(n_250),
.B1(n_244),
.B2(n_238),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_280),
.B1(n_300),
.B2(n_264),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_267),
.C(n_253),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_303),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_335),
.B(n_288),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_386),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_311),
.A2(n_257),
.B1(n_271),
.B2(n_235),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_308),
.B1(n_341),
.B2(n_314),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_340),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

BUFx24_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx13_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_325),
.Y(n_391)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_311),
.A2(n_17),
.B1(n_18),
.B2(n_0),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_308),
.B(n_0),
.C(n_18),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_401),
.Y(n_414)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_308),
.A2(n_328),
.B(n_319),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_358),
.B(n_351),
.Y(n_422)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_396),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_305),
.Y(n_397)
);

INVx3_ASAP7_75t_SL g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_318),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_399),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_326),
.B(n_354),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_302),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_302),
.B(n_350),
.Y(n_403)
);

OAI32xp33_ASAP7_75t_L g440 ( 
.A1(n_403),
.A2(n_346),
.A3(n_331),
.B1(n_329),
.B2(n_304),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_343),
.B1(n_332),
.B2(n_345),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_413),
.A2(n_419),
.B1(n_423),
.B2(n_431),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_364),
.A2(n_357),
.B(n_339),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_416),
.A2(n_422),
.B(n_402),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_430),
.B1(n_437),
.B2(n_373),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_385),
.A2(n_345),
.B1(n_358),
.B2(n_301),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_395),
.A2(n_301),
.B1(n_355),
.B2(n_330),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_357),
.B(n_330),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_368),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_SL g429 ( 
.A1(n_393),
.A2(n_357),
.B(n_317),
.C(n_355),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_331),
.B(n_390),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_359),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_379),
.A2(n_348),
.B1(n_317),
.B2(n_305),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_374),
.B(n_329),
.CI(n_317),
.CON(n_434),
.SN(n_434)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_382),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_381),
.A2(n_346),
.B1(n_315),
.B2(n_304),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_372),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_438),
.B(n_362),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_441),
.B(n_442),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_431),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_370),
.B1(n_402),
.B2(n_376),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_444),
.A2(n_450),
.B1(n_455),
.B2(n_460),
.Y(n_484)
);

OAI22x1_ASAP7_75t_SL g445 ( 
.A1(n_430),
.A2(n_425),
.B1(n_411),
.B2(n_412),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_445),
.A2(n_417),
.B1(n_435),
.B2(n_433),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_374),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_449),
.C(n_451),
.Y(n_477)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_447),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_361),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_461),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_380),
.C(n_401),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_398),
.C(n_384),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_452),
.A2(n_456),
.B(n_468),
.Y(n_488)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_394),
.C(n_396),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_465),
.C(n_466),
.Y(n_492)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_438),
.B(n_439),
.Y(n_479)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_426),
.A2(n_399),
.B1(n_367),
.B2(n_403),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_371),
.Y(n_461)
);

XOR2x2_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_375),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_421),
.Y(n_494)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_437),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_464),
.B(n_440),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_369),
.C(n_363),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_411),
.B(n_391),
.C(n_320),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_307),
.C(n_320),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_471),
.Y(n_480)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_469),
.Y(n_500)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_307),
.C(n_390),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_474),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_390),
.B1(n_397),
.B2(n_425),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_420),
.B1(n_422),
.B2(n_404),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_479),
.A2(n_481),
.B1(n_491),
.B2(n_495),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_415),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_502),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_462),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_487),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_452),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_417),
.B1(n_420),
.B2(n_413),
.Y(n_491)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_504),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_444),
.A2(n_420),
.B1(n_432),
.B2(n_435),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_433),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_471),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_468),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_497),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_450),
.A2(n_423),
.B1(n_419),
.B2(n_432),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_498),
.A2(n_503),
.B1(n_443),
.B2(n_452),
.Y(n_509)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_472),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_473),
.A2(n_443),
.B1(n_474),
.B2(n_460),
.Y(n_503)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_429),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_427),
.Y(n_505)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_506),
.A2(n_512),
.B(n_515),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_477),
.B(n_449),
.C(n_448),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_511),
.C(n_513),
.Y(n_533)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_503),
.A2(n_465),
.B1(n_456),
.B2(n_429),
.Y(n_510)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_496),
.C(n_476),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_497),
.A2(n_429),
.B(n_447),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_451),
.C(n_461),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_488),
.A2(n_429),
.B(n_409),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_522),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_504),
.B(n_424),
.Y(n_518)
);

XNOR2x1_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_500),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_498),
.A2(n_409),
.B1(n_406),
.B2(n_424),
.Y(n_519)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_409),
.C(n_427),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_521),
.C(n_526),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_480),
.C(n_494),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_480),
.B(n_478),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_488),
.A2(n_478),
.B(n_495),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_523),
.A2(n_500),
.B(n_501),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_485),
.C(n_484),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_475),
.Y(n_527)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_491),
.C(n_489),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_483),
.C(n_482),
.Y(n_541)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_475),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_502),
.Y(n_535)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_535),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_528),
.Y(n_536)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_536),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_483),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_538),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_483),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_482),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_539),
.B(n_544),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_541),
.B(n_542),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_490),
.C(n_493),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_490),
.C(n_493),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_543),
.B(n_531),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_549),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g548 ( 
.A1(n_507),
.A2(n_525),
.B(n_517),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_548),
.B(n_510),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_526),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_536),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_555),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_542),
.B(n_520),
.C(n_522),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_524),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_558),
.B(n_562),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_532),
.A2(n_545),
.B1(n_547),
.B2(n_509),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_559),
.A2(n_565),
.B1(n_545),
.B2(n_547),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_561),
.A2(n_515),
.B(n_537),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_539),
.B(n_513),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_521),
.C(n_516),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_566),
.C(n_533),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_532),
.A2(n_524),
.B1(n_529),
.B2(n_523),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_514),
.C(n_518),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_567),
.B(n_546),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_554),
.Y(n_568)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_569),
.B(n_570),
.Y(n_587)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_560),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_577),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_541),
.Y(n_573)
);

MAJx2_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_579),
.C(n_569),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_555),
.B(n_533),
.C(n_551),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_563),
.C(n_551),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_576),
.A2(n_553),
.B1(n_506),
.B2(n_564),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_538),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_534),
.B(n_512),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_578),
.A2(n_581),
.B(n_564),
.Y(n_585)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_560),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_535),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_554),
.A2(n_534),
.B(n_544),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_588),
.Y(n_593)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_583),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_585),
.A2(n_578),
.B(n_581),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_576),
.A2(n_565),
.B1(n_553),
.B2(n_559),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_590),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_550),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_591),
.B(n_585),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_506),
.C(n_519),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_592),
.B(n_573),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_597),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_586),
.A2(n_572),
.B(n_568),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_596),
.B(n_584),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_599),
.B(n_592),
.Y(n_604)
);

NOR2x1_ASAP7_75t_L g600 ( 
.A(n_598),
.B(n_583),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_600),
.B(n_601),
.C(n_604),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_593),
.B(n_582),
.C(n_571),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_602),
.B(n_594),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_606),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_595),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_607),
.A2(n_603),
.B(n_587),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_609),
.A2(n_605),
.B1(n_588),
.B2(n_589),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_608),
.C(n_550),
.Y(n_611)
);

FAx1_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_527),
.CI(n_501),
.CON(n_612),
.SN(n_612)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_514),
.Y(n_613)
);


endmodule