module fake_jpeg_12942_n_98 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_24),
.B(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_2),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_28),
.B1(n_38),
.B2(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_26),
.B1(n_39),
.B2(n_43),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_55),
.Y(n_67)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_32),
.B1(n_38),
.B2(n_37),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_3),
.C(n_4),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_29),
.B1(n_31),
.B2(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_27),
.Y(n_55)
);

AOI31xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.A3(n_50),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_45),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_31),
.B(n_29),
.C(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_52),
.B(n_6),
.Y(n_77)
);

AOI22x1_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_82),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_83),
.B1(n_5),
.B2(n_9),
.Y(n_87)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_70),
.B1(n_78),
.B2(n_10),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_88),
.B1(n_85),
.B2(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_9),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_10),
.C(n_11),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_83),
.C(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_89),
.C(n_84),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_11),
.B(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_13),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_13),
.Y(n_98)
);


endmodule