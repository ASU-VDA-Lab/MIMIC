module fake_jpeg_29254_n_487 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_54),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_0),
.C(n_2),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_61),
.B(n_62),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_68),
.Y(n_108)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_3),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_73),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_31),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_23),
.B1(n_43),
.B2(n_39),
.Y(n_153)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_91),
.Y(n_165)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_17),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_26),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_29),
.B(n_4),
.C(n_9),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_49),
.C(n_43),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_147),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_56),
.A2(n_51),
.B1(n_34),
.B2(n_36),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_114),
.A2(n_116),
.B1(n_139),
.B2(n_141),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_51),
.B1(n_34),
.B2(n_36),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_34),
.B1(n_51),
.B2(n_41),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_153),
.B1(n_162),
.B2(n_164),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_42),
.B1(n_52),
.B2(n_24),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_42),
.B1(n_52),
.B2(n_24),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_73),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_95),
.A2(n_49),
.B1(n_35),
.B2(n_28),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_104),
.A2(n_19),
.B1(n_20),
.B2(n_32),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_106),
.B1(n_83),
.B2(n_82),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_207),
.B1(n_211),
.B2(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_61),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_169),
.Y(n_238)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_68),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_160),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_174),
.B(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_28),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_178),
.B(n_188),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_107),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_165),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_74),
.B1(n_57),
.B2(n_55),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_192),
.B1(n_141),
.B2(n_163),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_63),
.B1(n_72),
.B2(n_67),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_23),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_194),
.B(n_199),
.Y(n_243)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_91),
.B(n_88),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_197),
.A2(n_138),
.B(n_25),
.Y(n_250)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_200),
.B(n_206),
.Y(n_248)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_35),
.Y(n_203)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_116),
.A2(n_65),
.B1(n_18),
.B2(n_27),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_26),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_91),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_123),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_25),
.B1(n_18),
.B2(n_19),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_123),
.Y(n_235)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_216),
.A2(n_211),
.B1(n_205),
.B2(n_186),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_113),
.B1(n_138),
.B2(n_134),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_210),
.B(n_197),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_122),
.B1(n_131),
.B2(n_159),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_232),
.B1(n_234),
.B2(n_167),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_181),
.A2(n_159),
.B1(n_119),
.B2(n_148),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_181),
.A2(n_119),
.B1(n_157),
.B2(n_148),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_191),
.B1(n_192),
.B2(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_132),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_210),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_145),
.A3(n_155),
.B1(n_133),
.B2(n_120),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_177),
.B(n_146),
.C(n_212),
.D(n_174),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_255),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_259),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_168),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_210),
.B1(n_132),
.B2(n_157),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_265),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_196),
.C(n_195),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_282),
.C(n_234),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_213),
.B1(n_180),
.B2(n_184),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_216),
.A2(n_201),
.B1(n_198),
.B2(n_202),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_279),
.B1(n_247),
.B2(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_221),
.B(n_171),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_281),
.B(n_262),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_SL g273 ( 
.A1(n_226),
.A2(n_190),
.B(n_170),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_247),
.Y(n_274)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_221),
.A2(n_143),
.B1(n_185),
.B2(n_179),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_220),
.B1(n_218),
.B2(n_224),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_240),
.B(n_19),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_19),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_217),
.A2(n_204),
.B1(n_182),
.B2(n_179),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_219),
.B(n_227),
.C(n_231),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_182),
.C(n_204),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_287),
.B1(n_296),
.B2(n_261),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_243),
.B(n_231),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_286),
.A2(n_307),
.B(n_309),
.C(n_272),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_246),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_299),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_282),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_246),
.B(n_238),
.C(n_222),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_260),
.B(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_290),
.B1(n_311),
.B2(n_282),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_267),
.A2(n_238),
.B1(n_249),
.B2(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_218),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_301),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_251),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_220),
.C(n_230),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_310),
.C(n_239),
.Y(n_332)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_311),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_236),
.B(n_230),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_281),
.A2(n_236),
.B(n_223),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_233),
.C(n_223),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_239),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_303),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_304),
.B(n_286),
.C(n_308),
.D(n_309),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_308),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_315),
.A2(n_316),
.B1(n_295),
.B2(n_303),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_263),
.B1(n_273),
.B2(n_253),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_332),
.C(n_310),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_318),
.A2(n_327),
.B(n_339),
.Y(n_363)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_275),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_329),
.B1(n_334),
.B2(n_297),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_325),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_293),
.A2(n_255),
.B1(n_267),
.B2(n_269),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_330),
.B1(n_331),
.B2(n_283),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_272),
.B(n_279),
.C(n_274),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_265),
.B(n_264),
.C(n_268),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_296),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_242),
.B1(n_245),
.B2(n_251),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_291),
.B1(n_303),
.B2(n_298),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_302),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_333),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_233),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_228),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_228),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_336),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_288),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_294),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_338),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_340),
.Y(n_368)
);

XOR2x2_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_344),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_305),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_318),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_345),
.B(n_318),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_326),
.B1(n_318),
.B2(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_285),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_324),
.Y(n_351)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_332),
.C(n_323),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_358),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_359),
.B1(n_367),
.B2(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_361),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_292),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_325),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_315),
.B(n_316),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_361),
.A2(n_330),
.B(n_313),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_357),
.B1(n_346),
.B2(n_363),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_382),
.C(n_386),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_380),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_389),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_388),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_327),
.B(n_325),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_385),
.A2(n_358),
.B(n_341),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_292),
.C(n_288),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_306),
.C(n_301),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_362),
.C(n_348),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_327),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_340),
.Y(n_389)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_294),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_366),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_285),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_349),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_377),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_405),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_387),
.B(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_400),
.B(n_401),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_376),
.B(n_343),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_369),
.B1(n_379),
.B2(n_371),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_363),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_386),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_407),
.C(n_409),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_351),
.C(n_350),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_353),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_343),
.C(n_341),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_384),
.Y(n_411)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_379),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_368),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_413),
.A2(n_402),
.B(n_410),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_418),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_420),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_393),
.B1(n_372),
.B2(n_373),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_392),
.C(n_388),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_32),
.C(n_10),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_384),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_409),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_383),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_402),
.A2(n_385),
.B(n_373),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_427),
.A2(n_416),
.B(n_429),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_430),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_380),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_410),
.A2(n_369),
.B1(n_383),
.B2(n_347),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_4),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_394),
.C(n_396),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_436),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_442),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_419),
.C(n_421),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_438),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_407),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_443),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_440),
.A2(n_444),
.B(n_445),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_395),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_405),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_406),
.C(n_414),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_414),
.C(n_19),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_446),
.A2(n_429),
.B1(n_422),
.B2(n_430),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_431),
.C(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_448),
.B(n_452),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_437),
.B(n_425),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_459),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_432),
.B(n_428),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_457),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_435),
.B(n_9),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_32),
.C(n_10),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_450),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_446),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_11),
.B(n_13),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_460),
.A2(n_11),
.B(n_14),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_465),
.Y(n_475)
);

AO21x1_ASAP7_75t_L g476 ( 
.A1(n_462),
.A2(n_468),
.B(n_470),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_456),
.A2(n_442),
.B(n_441),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_463),
.A2(n_448),
.B(n_458),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_441),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_447),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_459),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_449),
.A2(n_14),
.B(n_15),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_14),
.C(n_15),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_451),
.Y(n_471)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_464),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_472),
.A2(n_477),
.B(n_469),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_474),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_32),
.C(n_14),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_470),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_479),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_475),
.C(n_476),
.Y(n_483)
);

NAND2x1_ASAP7_75t_SL g484 ( 
.A(n_483),
.B(n_478),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_484),
.A2(n_482),
.B(n_480),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g486 ( 
.A(n_485),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_486),
.A2(n_15),
.B(n_32),
.Y(n_487)
);


endmodule