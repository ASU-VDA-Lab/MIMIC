module fake_ariane_1451_n_3437 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_913, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_943, n_678, n_651, n_936, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_878, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_908, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_906, n_416, n_283, n_919, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_924, n_927, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_864, n_952, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_940, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_897, n_32, n_949, n_956, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_891, n_737, n_137, n_885, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_917, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_870, n_87, n_714, n_279, n_905, n_702, n_945, n_958, n_207, n_790, n_857, n_898, n_363, n_720, n_354, n_41, n_813, n_926, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_900, n_154, n_883, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_871, n_315, n_903, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_879, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_855, n_158, n_69, n_259, n_835, n_95, n_808, n_953, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_858, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_928, n_3, n_271, n_465, n_486, n_507, n_901, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_894, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_868, n_326, n_681, n_778, n_227, n_48, n_874, n_188, n_323, n_550, n_635, n_707, n_330, n_914, n_400, n_689, n_694, n_884, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_921, n_620, n_228, n_325, n_276, n_93, n_688, n_859, n_636, n_427, n_108, n_587, n_497, n_693, n_863, n_303, n_671, n_442, n_777, n_929, n_168, n_81, n_1, n_206, n_352, n_538, n_899, n_920, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_887, n_661, n_488, n_775, n_667, n_300, n_533, n_904, n_505, n_14, n_163, n_88, n_869, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_957, n_512, n_715, n_889, n_935, n_579, n_844, n_459, n_685, n_221, n_321, n_911, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_861, n_175, n_950, n_711, n_877, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_942, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_907, n_235, n_881, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_941, n_700, n_910, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_939, n_371, n_845, n_888, n_199, n_918, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_865, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_948, n_582, n_94, n_284, n_922, n_4, n_448, n_593, n_755, n_710, n_860, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_890, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_896, n_409, n_171, n_947, n_930, n_519, n_902, n_384, n_468, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_872, n_933, n_13, n_27, n_916, n_254, n_596, n_954, n_912, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_915, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_955, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_951, n_213, n_938, n_862, n_110, n_304, n_895, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_946, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_875, n_669, n_785, n_827, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_937, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_880, n_793, n_852, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_873, n_51, n_496, n_739, n_76, n_342, n_866, n_26, n_246, n_517, n_925, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_892, n_608, n_959, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_923, n_250, n_932, n_773, n_165, n_144, n_882, n_317, n_867, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_944, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_856, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_876, n_618, n_411, n_484, n_712, n_849, n_909, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_893, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_854, n_471, n_351, n_886, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_934, n_783, n_675, n_3437);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_913;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_943;
input n_678;
input n_651;
input n_936;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_878;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_908;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_906;
input n_416;
input n_283;
input n_919;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_924;
input n_927;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_864;
input n_952;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_940;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_897;
input n_32;
input n_949;
input n_956;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_891;
input n_737;
input n_137;
input n_885;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_917;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_870;
input n_87;
input n_714;
input n_279;
input n_905;
input n_702;
input n_945;
input n_958;
input n_207;
input n_790;
input n_857;
input n_898;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_926;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_900;
input n_154;
input n_883;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_871;
input n_315;
input n_903;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_879;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_855;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_953;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_858;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_928;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_901;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_894;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_868;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_874;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_914;
input n_400;
input n_689;
input n_694;
input n_884;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_921;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_859;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_863;
input n_303;
input n_671;
input n_442;
input n_777;
input n_929;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_899;
input n_920;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_887;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_904;
input n_505;
input n_14;
input n_163;
input n_88;
input n_869;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_957;
input n_512;
input n_715;
input n_889;
input n_935;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_911;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_861;
input n_175;
input n_950;
input n_711;
input n_877;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_942;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_907;
input n_235;
input n_881;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_941;
input n_700;
input n_910;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_939;
input n_371;
input n_845;
input n_888;
input n_199;
input n_918;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_865;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_948;
input n_582;
input n_94;
input n_284;
input n_922;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_860;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_890;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_896;
input n_409;
input n_171;
input n_947;
input n_930;
input n_519;
input n_902;
input n_384;
input n_468;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_872;
input n_933;
input n_13;
input n_27;
input n_916;
input n_254;
input n_596;
input n_954;
input n_912;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_915;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_955;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_951;
input n_213;
input n_938;
input n_862;
input n_110;
input n_304;
input n_895;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_875;
input n_669;
input n_785;
input n_827;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_937;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_880;
input n_793;
input n_852;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_873;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_866;
input n_26;
input n_246;
input n_517;
input n_925;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_892;
input n_608;
input n_959;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_923;
input n_250;
input n_932;
input n_773;
input n_165;
input n_144;
input n_882;
input n_317;
input n_867;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_944;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_856;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_876;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_909;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_893;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_854;
input n_471;
input n_351;
input n_886;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_934;
input n_783;
input n_675;

output n_3437;

wire n_2752;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_3416;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3063;
wire n_3281;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_3270;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_2370;
wire n_1944;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_1254;
wire n_3207;
wire n_2433;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1790;
wire n_1354;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_3126;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3119;
wire n_1108;
wire n_1590;
wire n_1351;
wire n_3234;
wire n_3280;
wire n_3413;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_2134;
wire n_1260;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_2791;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3159;
wire n_992;
wire n_966;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_1292;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3372;
wire n_1623;
wire n_990;
wire n_1903;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3179;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_2718;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3286;
wire n_3370;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2496;
wire n_1614;
wire n_1162;
wire n_1377;
wire n_2418;
wire n_2031;
wire n_3260;
wire n_3349;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_3290;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_1242;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_2949;
wire n_2300;
wire n_2894;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3423;
wire n_1975;
wire n_1373;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3333;
wire n_1860;
wire n_1734;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_3024;
wire n_2772;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3097;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2723;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_1657;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_2546;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2890;
wire n_3381;
wire n_3313;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_3345;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1603;
wire n_1370;
wire n_2935;
wire n_2401;
wire n_3255;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_2886;
wire n_2478;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_3396;
wire n_1210;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_1968;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_3363;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_1653;
wire n_3409;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3241;
wire n_1584;
wire n_1157;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_3106;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3402;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3410;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3269;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3248;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3431;
wire n_2176;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_2012;
wire n_1937;
wire n_3182;
wire n_2967;
wire n_1064;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3232;
wire n_3001;
wire n_3188;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1684;
wire n_1588;
wire n_1409;
wire n_1148;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_3366;
wire n_2430;
wire n_2504;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_2017;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3293;
wire n_3361;
wire n_1683;
wire n_1229;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_1891;
wire n_1328;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_2047;
wire n_3058;
wire n_2792;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3075;
wire n_3030;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3308;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g960 ( 
.A(n_189),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_71),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_318),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_193),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_662),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_567),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_390),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

CKINVDCx16_ASAP7_75t_R g968 ( 
.A(n_893),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_167),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_792),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_345),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_747),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_820),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_24),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_889),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_753),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_777),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_916),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_256),
.B(n_911),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_122),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_913),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_785),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_386),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_885),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_819),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_746),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_496),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_257),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_894),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_457),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_349),
.Y(n_991)
);

CKINVDCx16_ASAP7_75t_R g992 ( 
.A(n_518),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_565),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_784),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_29),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_794),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_732),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_15),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_813),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_601),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_545),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_748),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_625),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_896),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_695),
.Y(n_1005)
);

CKINVDCx16_ASAP7_75t_R g1006 ( 
.A(n_73),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_426),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_55),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_918),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_40),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_253),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_807),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_898),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_186),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_31),
.B(n_703),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_760),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_947),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_252),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_625),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_206),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_773),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_589),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_880),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_884),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_248),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_829),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_689),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_445),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_192),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_225),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_864),
.Y(n_1031)
);

CKINVDCx14_ASAP7_75t_R g1032 ( 
.A(n_942),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_795),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_917),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_646),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_241),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_862),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_206),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_526),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_487),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_834),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_192),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_111),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_152),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_369),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_853),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_51),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_325),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_66),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_299),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_331),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_59),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_354),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_546),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_338),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_846),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_865),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_827),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_596),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_821),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_261),
.Y(n_1061)
);

BUFx8_ASAP7_75t_SL g1062 ( 
.A(n_342),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_630),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_957),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_327),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_706),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_941),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_27),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_729),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_676),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_522),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_830),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_728),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_892),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_84),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_163),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_342),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_848),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_905),
.Y(n_1079)
);

BUFx5_ASAP7_75t_L g1080 ( 
.A(n_783),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_423),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_655),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_713),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_39),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_286),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_808),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_512),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_796),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_737),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_798),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_936),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_126),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_247),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_389),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_10),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_851),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_492),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_226),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_602),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_809),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_197),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_453),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_445),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_543),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_750),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_682),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_882),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_540),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_513),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_298),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_940),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_850),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_845),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_595),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_408),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_719),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_65),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_900),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_912),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_915),
.Y(n_1120)
);

BUFx5_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_92),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_142),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_550),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_788),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_888),
.Y(n_1126)
);

BUFx8_ASAP7_75t_SL g1127 ( 
.A(n_498),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_401),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_642),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_125),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_477),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_841),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_297),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_847),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_455),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_685),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_300),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_887),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_34),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_875),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_860),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_805),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_480),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_636),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_537),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_211),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_519),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_831),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_786),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_800),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_62),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_654),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_549),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_473),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_42),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_326),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_L g1157 ( 
.A(n_815),
.B(n_361),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_162),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_495),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_344),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_424),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_790),
.Y(n_1162)
);

CKINVDCx14_ASAP7_75t_R g1163 ( 
.A(n_929),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_491),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_367),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_171),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_239),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_870),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_811),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_842),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_874),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_31),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_930),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_932),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_623),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_338),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_233),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_171),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_450),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_26),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_791),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_836),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_824),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_277),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_946),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_5),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_382),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_327),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_569),
.B(n_260),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_793),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_802),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_602),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_700),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_392),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_787),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_496),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_804),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_55),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_838),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_153),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_468),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_903),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_876),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_111),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_243),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_814),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_514),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_596),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_16),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_473),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_944),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_277),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_505),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_844),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_46),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_414),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_512),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_545),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_161),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_126),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_895),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_883),
.Y(n_1222)
);

CKINVDCx14_ASAP7_75t_R g1223 ( 
.A(n_878),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_183),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_482),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_858),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_949),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_16),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_525),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_593),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_856),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_897),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_7),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_928),
.Y(n_1234)
);

BUFx8_ASAP7_75t_SL g1235 ( 
.A(n_180),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_938),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_34),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_891),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_268),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_27),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_245),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_852),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_610),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_613),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_859),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_13),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_779),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_477),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_494),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_843),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_461),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_101),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_294),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_43),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_197),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_855),
.Y(n_1256)
);

CKINVDCx16_ASAP7_75t_R g1257 ( 
.A(n_137),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_202),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_872),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_24),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_910),
.B(n_677),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_347),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_835),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_863),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_931),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_364),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_467),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_475),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_909),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_630),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_945),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_610),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_248),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_142),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_209),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_879),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_837),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_344),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_839),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_516),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_881),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_765),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_414),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_948),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_854),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_914),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_561),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_866),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_840),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_70),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_451),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_871),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_207),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_816),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_203),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_449),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_313),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_538),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_511),
.Y(n_1299)
);

BUFx5_ASAP7_75t_L g1300 ( 
.A(n_253),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_828),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_257),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_907),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_22),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_886),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_923),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_833),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_803),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_517),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_6),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_518),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_935),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_184),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_812),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_801),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_857),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_483),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_925),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_116),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_255),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_459),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_183),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_424),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_202),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_135),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_175),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_458),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_141),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_937),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_733),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_823),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_201),
.Y(n_1332)
);

BUFx8_ASAP7_75t_SL g1333 ( 
.A(n_659),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_902),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_906),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_922),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_825),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_340),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_301),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_593),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_223),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_687),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_956),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_899),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_797),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_959),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_265),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_49),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_213),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_52),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_585),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_954),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_921),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_601),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_868),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_411),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_530),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_806),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_901),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_658),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_335),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_642),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_849),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_220),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_4),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_587),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_423),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_771),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_403),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_867),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_446),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_920),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_64),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_904),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_869),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_205),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_908),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_407),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_365),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_117),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_933),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_799),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_555),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_861),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_832),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_454),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_873),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_567),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_557),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_609),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_684),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_163),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_232),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_943),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_822),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_552),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_114),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_640),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_810),
.B(n_694),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_926),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_924),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_919),
.B(n_939),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_193),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_877),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_675),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_141),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_215),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_525),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_399),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_65),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_167),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_817),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_890),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_353),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_156),
.B(n_349),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_789),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_818),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_504),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_621),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_927),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_316),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_952),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_934),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_708),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_826),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_275),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_589),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_51),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_367),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_R g1430 ( 
.A(n_1032),
.B(n_649),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1300),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1055),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1004),
.A2(n_1005),
.B1(n_1060),
.B2(n_1027),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_965),
.B(n_0),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1066),
.B(n_0),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_1062),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1203),
.B(n_1),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1043),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1016),
.A2(n_651),
.B(n_650),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1300),
.Y(n_1440)
);

BUFx8_ASAP7_75t_SL g1441 ( 
.A(n_1127),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1160),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1194),
.Y(n_1443)
);

INVx5_ASAP7_75t_L g1444 ( 
.A(n_1120),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1300),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1180),
.B(n_1),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1311),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1392),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1259),
.B(n_3),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1055),
.Y(n_1450)
);

BUFx8_ASAP7_75t_SL g1451 ( 
.A(n_1235),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1247),
.B(n_2),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1053),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1055),
.Y(n_1454)
);

AOI22x1_ASAP7_75t_SL g1455 ( 
.A1(n_974),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1300),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1120),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1053),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1343),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1098),
.B(n_1099),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_992),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1006),
.B(n_5),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1112),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1300),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1147),
.B(n_6),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1343),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1097),
.Y(n_1467)
);

BUFx8_ASAP7_75t_SL g1468 ( 
.A(n_995),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1359),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1359),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1097),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1333),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1028),
.B(n_7),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1257),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1097),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1204),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_960),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1164),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1164),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1340),
.Y(n_1480)
);

BUFx8_ASAP7_75t_L g1481 ( 
.A(n_1035),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1367),
.B(n_8),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_SL g1483 ( 
.A(n_968),
.B(n_652),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1413),
.B(n_9),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1021),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1274),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1204),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_964),
.B(n_8),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1280),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_962),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1191),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_967),
.B(n_9),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1164),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1165),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1280),
.B(n_10),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_963),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1165),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1313),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1165),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1418),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1199),
.Y(n_1501)
);

INVx5_ASAP7_75t_L g1502 ( 
.A(n_1207),
.Y(n_1502)
);

BUFx12f_ASAP7_75t_L g1503 ( 
.A(n_1313),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1317),
.Y(n_1504)
);

AND2x6_ASAP7_75t_L g1505 ( 
.A(n_1088),
.B(n_653),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_966),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1207),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1207),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1218),
.B(n_11),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1225),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1000),
.B(n_11),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1317),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1225),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1007),
.B(n_12),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1328),
.B(n_12),
.Y(n_1515)
);

OAI22x1_ASAP7_75t_SL g1516 ( 
.A1(n_1001),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_978),
.A2(n_994),
.B(n_981),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1010),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1236),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1014),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1019),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1225),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1029),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1030),
.B(n_14),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1320),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1320),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_999),
.B(n_17),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1034),
.B(n_17),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1039),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1320),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1324),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_969),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1324),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1324),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1328),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1411),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1042),
.B(n_18),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1054),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1061),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1076),
.B(n_18),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1081),
.B(n_19),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1357),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1357),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1411),
.B(n_19),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1357),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1084),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1250),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1373),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1100),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_971),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_980),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1087),
.B(n_20),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1092),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1093),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1373),
.Y(n_1555)
);

AND2x6_ASAP7_75t_L g1556 ( 
.A(n_1106),
.B(n_656),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1152),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1094),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1102),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1373),
.Y(n_1560)
);

BUFx2_ASAP7_75t_SL g1561 ( 
.A(n_1472),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1432),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1491),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1501),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1463),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1519),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1431),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1436),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_R g1569 ( 
.A(n_1483),
.B(n_1163),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1445),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1500),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1450),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1441),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1451),
.Y(n_1574)
);

XNOR2xp5_ASAP7_75t_L g1575 ( 
.A(n_1433),
.B(n_1124),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1454),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1468),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1489),
.Y(n_1578)
);

BUFx10_ASAP7_75t_L g1579 ( 
.A(n_1449),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1472),
.B(n_1423),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1480),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_R g1582 ( 
.A(n_1458),
.B(n_1223),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1457),
.Y(n_1583)
);

CKINVDCx6p67_ASAP7_75t_R g1584 ( 
.A(n_1503),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1504),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1456),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1440),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1439),
.A2(n_1402),
.B(n_1058),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1464),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1467),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1535),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1459),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1477),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1471),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1466),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1490),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1551),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1496),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1485),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1557),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1461),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1444),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1444),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1518),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1474),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1506),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_R g1607 ( 
.A(n_1476),
.B(n_1335),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1475),
.Y(n_1608)
);

BUFx10_ASAP7_75t_L g1609 ( 
.A(n_1484),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_1462),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1469),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1469),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_R g1613 ( 
.A(n_1487),
.B(n_1346),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1520),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1523),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1513),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1470),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1513),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_R g1619 ( 
.A(n_1512),
.B(n_1360),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1479),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1529),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1470),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1538),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1539),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1532),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1546),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1550),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1536),
.B(n_961),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1481),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1493),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1486),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1494),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1553),
.Y(n_1633)
);

AOI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1517),
.A2(n_1067),
.B(n_1057),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1554),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1430),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1460),
.B(n_1003),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1558),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1559),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1549),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_R g1641 ( 
.A(n_1453),
.B(n_1417),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_R g1642 ( 
.A(n_1498),
.B(n_1119),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1438),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1442),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1497),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1581),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1588),
.A2(n_1492),
.B(n_1488),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1567),
.B(n_1505),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1587),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1636),
.B(n_1473),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1631),
.B(n_1447),
.Y(n_1651)
);

AO221x1_ASAP7_75t_L g1652 ( 
.A1(n_1644),
.A2(n_1426),
.B1(n_1270),
.B2(n_1184),
.C(n_1521),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1596),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1598),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1599),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1570),
.B(n_1586),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1589),
.B(n_1604),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1505),
.Y(n_1659)
);

NAND2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1569),
.B(n_1482),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1592),
.B(n_1435),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1637),
.A2(n_1515),
.B1(n_1544),
.B2(n_1495),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1579),
.A2(n_1437),
.B1(n_1446),
.B2(n_1434),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1615),
.B(n_1556),
.Y(n_1665)
);

BUFx5_ASAP7_75t_L g1666 ( 
.A(n_1621),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1571),
.B(n_1452),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1623),
.B(n_1556),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1626),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1633),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1595),
.B(n_1509),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1638),
.B(n_1555),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1600),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1642),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1597),
.B(n_1443),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1634),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1555),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1609),
.B(n_1527),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1582),
.B(n_1511),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1628),
.B(n_1514),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1609),
.B(n_1528),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1610),
.B(n_1258),
.C(n_1249),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1579),
.B(n_1465),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1562),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1625),
.Y(n_1688)
);

NOR2xp67_ASAP7_75t_L g1689 ( 
.A(n_1583),
.B(n_1502),
.Y(n_1689)
);

BUFx2_ASAP7_75t_R g1690 ( 
.A(n_1568),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1641),
.B(n_1524),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1607),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1628),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1637),
.B(n_1537),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1572),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1576),
.Y(n_1696)
);

BUFx5_ASAP7_75t_L g1697 ( 
.A(n_1618),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1602),
.B(n_1540),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1613),
.B(n_1541),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1619),
.B(n_1552),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1601),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_L g1702 ( 
.A(n_1563),
.B(n_1015),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1608),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_SL g1704 ( 
.A(n_1564),
.B(n_1044),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1605),
.B(n_1448),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_L g1706 ( 
.A(n_1566),
.B(n_1547),
.C(n_1244),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1585),
.B(n_1289),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1603),
.B(n_1478),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1643),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_L g1710 ( 
.A(n_1611),
.B(n_1189),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1620),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1630),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1612),
.B(n_983),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1632),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_L g1715 ( 
.A(n_1573),
.B(n_1321),
.C(n_1036),
.Y(n_1715)
);

XOR2xp5_ASAP7_75t_L g1716 ( 
.A(n_1565),
.B(n_1455),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1645),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1590),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1617),
.B(n_1510),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1606),
.B(n_1522),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1590),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1622),
.B(n_1499),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1561),
.B(n_1580),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1627),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1590),
.B(n_1525),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1594),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1584),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1594),
.B(n_1507),
.Y(n_1728)
);

NOR2xp67_ASAP7_75t_L g1729 ( 
.A(n_1591),
.B(n_1574),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1594),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1629),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1575),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1578),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1681),
.A2(n_1415),
.B1(n_987),
.B2(n_990),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1690),
.B(n_1577),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1667),
.B(n_988),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1649),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1653),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1646),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1663),
.A2(n_1085),
.B1(n_1135),
.B2(n_1052),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1669),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1716),
.A2(n_1212),
.B1(n_1278),
.B2(n_1210),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1656),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1684),
.B(n_996),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1677),
.B(n_991),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1675),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1666),
.B(n_997),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1664),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1654),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1666),
.B(n_1107),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1664),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1666),
.B(n_1222),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1720),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1670),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1692),
.B(n_1362),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1702),
.A2(n_1298),
.B1(n_1326),
.B2(n_1287),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_SL g1758 ( 
.A(n_1686),
.B(n_998),
.C(n_993),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1688),
.B(n_1364),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1701),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1682),
.B(n_1008),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_SL g1762 ( 
.A(n_1704),
.B(n_1341),
.C(n_1327),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1666),
.B(n_1011),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1655),
.B(n_1370),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1671),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1676),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1673),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1724),
.B(n_1516),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1727),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1709),
.B(n_1376),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1687),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1658),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1651),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1695),
.Y(n_1774)
);

INVx5_ASAP7_75t_L g1775 ( 
.A(n_1678),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1705),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1657),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1662),
.B(n_1018),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1659),
.B(n_1022),
.Y(n_1779)
);

NAND2x1p5_ASAP7_75t_L g1780 ( 
.A(n_1729),
.B(n_1530),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1718),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1706),
.A2(n_1403),
.B1(n_1410),
.B2(n_1406),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1665),
.B(n_1025),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1721),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1696),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1726),
.Y(n_1786)
);

AND2x6_ASAP7_75t_L g1787 ( 
.A(n_1668),
.B(n_1070),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1648),
.B(n_1073),
.Y(n_1788)
);

AND3x2_ASAP7_75t_SL g1789 ( 
.A(n_1712),
.B(n_1101),
.C(n_1020),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1647),
.A2(n_1157),
.B(n_979),
.C(n_1109),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1661),
.B(n_1366),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1694),
.B(n_1038),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1660),
.B(n_1040),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1731),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1703),
.Y(n_1795)
);

INVx5_ASAP7_75t_L g1796 ( 
.A(n_1689),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1707),
.B(n_1693),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_SL g1798 ( 
.A(n_1715),
.B(n_1047),
.C(n_1045),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1710),
.A2(n_1318),
.B1(n_1111),
.B2(n_1125),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1650),
.B(n_1048),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1728),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1730),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1683),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1711),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1691),
.B(n_1049),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1685),
.A2(n_1126),
.B1(n_1134),
.B2(n_1086),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1697),
.B(n_1700),
.Y(n_1807)
);

AND3x1_ASAP7_75t_L g1808 ( 
.A(n_1698),
.B(n_1128),
.C(n_1104),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1719),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1699),
.B(n_1427),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1697),
.B(n_1050),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1697),
.B(n_1680),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1697),
.B(n_1051),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1672),
.A2(n_1150),
.B1(n_1162),
.B2(n_1149),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1652),
.A2(n_1192),
.B1(n_1201),
.B2(n_1133),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1714),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1708),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1717),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1674),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1722),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1679),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1713),
.B(n_1723),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1725),
.B(n_1059),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1732),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1681),
.B(n_1063),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1667),
.B(n_1065),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1646),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1656),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1678),
.B(n_1508),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1656),
.B(n_1144),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1653),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1656),
.B(n_1145),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_SL g1833 ( 
.A(n_1663),
.B(n_1071),
.C(n_1068),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1653),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1649),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1653),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1667),
.B(n_1075),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1649),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1647),
.A2(n_1170),
.B(n_1168),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1656),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1653),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1667),
.B(n_1077),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1681),
.B(n_1095),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1649),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1646),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1653),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1649),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1656),
.Y(n_1848)
);

NAND2x2_ASAP7_75t_L g1849 ( 
.A(n_1733),
.B(n_1103),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1656),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1667),
.B(n_1108),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1656),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1656),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1664),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1667),
.B(n_1110),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1667),
.B(n_1114),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1667),
.B(n_1115),
.Y(n_1857)
);

INVx6_ASAP7_75t_L g1858 ( 
.A(n_1720),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1656),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1667),
.B(n_1117),
.Y(n_1860)
);

INVxp67_ASAP7_75t_SL g1861 ( 
.A(n_1646),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1649),
.Y(n_1862)
);

AND2x6_ASAP7_75t_SL g1863 ( 
.A(n_1678),
.B(n_1179),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1656),
.B(n_1175),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1646),
.Y(n_1865)
);

AND2x6_ASAP7_75t_L g1866 ( 
.A(n_1656),
.B(n_1173),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1653),
.Y(n_1867)
);

OR2x6_ASAP7_75t_L g1868 ( 
.A(n_1724),
.B(n_1230),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1649),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1716),
.A2(n_1155),
.B1(n_1220),
.B2(n_1130),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1667),
.B(n_1122),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1656),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1667),
.B(n_1123),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1825),
.B(n_1178),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_SL g1875 ( 
.A(n_1735),
.B(n_1129),
.Y(n_1875)
);

AOI221x1_ASAP7_75t_L g1876 ( 
.A1(n_1790),
.A2(n_1185),
.B1(n_1190),
.B2(n_1182),
.C(n_1174),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1738),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1839),
.A2(n_1211),
.B(n_1197),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1843),
.A2(n_1232),
.B(n_1245),
.C(n_1226),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1821),
.A2(n_972),
.B(n_970),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_R g1881 ( 
.A(n_1743),
.B(n_1131),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1749),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1744),
.B(n_1188),
.Y(n_1883)
);

NOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1840),
.B(n_1263),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1769),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1866),
.A2(n_1139),
.B1(n_1143),
.B2(n_1137),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1767),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1777),
.B(n_1196),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1763),
.A2(n_975),
.B(n_973),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1826),
.A2(n_1301),
.B(n_1307),
.C(n_1284),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1737),
.Y(n_1891)
);

NOR2xp67_ASAP7_75t_L g1892 ( 
.A(n_1853),
.B(n_1533),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1772),
.B(n_1208),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1827),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1835),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1776),
.B(n_1531),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1775),
.B(n_1773),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1760),
.B(n_1526),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1831),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1848),
.B(n_1534),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1739),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1775),
.B(n_1146),
.Y(n_1902)
);

A2O1A1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1837),
.A2(n_1312),
.B(n_1315),
.C(n_1308),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1838),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1756),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1834),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1748),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1812),
.A2(n_977),
.B(n_976),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1842),
.B(n_1209),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1836),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1756),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1860),
.B(n_1224),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1828),
.B(n_1151),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1871),
.B(n_1229),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1873),
.A2(n_1352),
.B(n_1334),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1740),
.A2(n_1291),
.B1(n_1299),
.B2(n_1272),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1841),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1759),
.A2(n_1375),
.B1(n_1387),
.B2(n_1358),
.Y(n_1918)
);

O2A1O1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1734),
.A2(n_1241),
.B(n_1243),
.C(n_1239),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1846),
.B(n_1252),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1867),
.A2(n_1154),
.B1(n_1156),
.B2(n_1153),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1858),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1845),
.Y(n_1923)
);

NAND2x1p5_ASAP7_75t_L g1924 ( 
.A(n_1850),
.B(n_1545),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1755),
.B(n_1253),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1741),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1844),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1779),
.A2(n_984),
.B(n_982),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1820),
.B(n_1267),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1852),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1791),
.A2(n_1405),
.B(n_1395),
.C(n_1273),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1847),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1862),
.Y(n_1933)
);

OR2x6_ASAP7_75t_SL g1934 ( 
.A(n_1794),
.B(n_1167),
.Y(n_1934)
);

AOI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1747),
.A2(n_1399),
.B(n_1261),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1817),
.B(n_1302),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1754),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1859),
.B(n_1158),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1872),
.B(n_1310),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1757),
.B(n_1339),
.C(n_1248),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1803),
.B(n_1325),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1748),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1764),
.B(n_1332),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1805),
.A2(n_1351),
.B(n_1356),
.C(n_1338),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1765),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1746),
.B(n_1766),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1799),
.A2(n_1161),
.B1(n_1166),
.B2(n_1159),
.Y(n_1947)
);

INVx4_ASAP7_75t_L g1948 ( 
.A(n_1751),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1865),
.B(n_1172),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1829),
.B(n_1542),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1810),
.A2(n_1380),
.B(n_1386),
.C(n_1378),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1751),
.Y(n_1952)
);

A2O1A1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1750),
.A2(n_1390),
.B(n_1393),
.C(n_1389),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1869),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_SL g1955 ( 
.A(n_1758),
.B(n_1177),
.C(n_1176),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1854),
.B(n_1548),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1801),
.B(n_1397),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1753),
.B(n_1398),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1833),
.A2(n_1187),
.B1(n_1198),
.B2(n_1186),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1861),
.B(n_1543),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1766),
.B(n_1200),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1770),
.B(n_1560),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1736),
.B(n_1205),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1783),
.A2(n_986),
.B(n_985),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1854),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1752),
.A2(n_1414),
.B(n_1407),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1851),
.B(n_1213),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1830),
.B(n_1428),
.Y(n_1968)
);

OAI21xp33_ASAP7_75t_L g1969 ( 
.A1(n_1792),
.A2(n_1304),
.B(n_1290),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1813),
.A2(n_1856),
.B(n_1855),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1857),
.A2(n_1002),
.B(n_989),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1809),
.B(n_1429),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1868),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1807),
.A2(n_1216),
.B1(n_1217),
.B2(n_1215),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1866),
.B(n_1219),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1824),
.B(n_1228),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1761),
.A2(n_1369),
.B(n_1361),
.C(n_1026),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1782),
.A2(n_1240),
.B1(n_1246),
.B2(n_1237),
.C(n_1233),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1868),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1771),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1832),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1785),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1864),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1774),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1797),
.B(n_1251),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1819),
.B(n_1254),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1811),
.A2(n_1012),
.B(n_1009),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1866),
.B(n_1787),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1778),
.A2(n_1260),
.B1(n_1262),
.B2(n_1255),
.Y(n_1989)
);

NOR2xp67_ASAP7_75t_L g1990 ( 
.A(n_1796),
.B(n_1013),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1814),
.B(n_1266),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1796),
.B(n_1202),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1863),
.Y(n_1993)
);

AOI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1822),
.A2(n_1024),
.B(n_1017),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1795),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1786),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1793),
.A2(n_1033),
.B(n_1031),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1802),
.B(n_1268),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1800),
.A2(n_1041),
.B(n_1037),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1762),
.B(n_1275),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1804),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_L g2002 ( 
.A(n_1798),
.B(n_1238),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1806),
.B(n_1283),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1787),
.B(n_1293),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1780),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1816),
.Y(n_2006)
);

BUFx4f_ASAP7_75t_L g2007 ( 
.A(n_1781),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1745),
.A2(n_1296),
.B1(n_1297),
.B2(n_1295),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1818),
.A2(n_1319),
.B(n_1354),
.C(n_1322),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1823),
.A2(n_1069),
.B(n_1064),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1781),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1784),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1808),
.B(n_1309),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1784),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1787),
.A2(n_1074),
.B(n_1072),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1788),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1788),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1815),
.A2(n_1347),
.B1(n_1348),
.B2(n_1323),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1768),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1788),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1768),
.B(n_1349),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_SL g2022 ( 
.A1(n_1742),
.A2(n_1365),
.B1(n_1371),
.B2(n_1350),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1870),
.B(n_1379),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1789),
.Y(n_2024)
);

INVxp67_ASAP7_75t_L g2025 ( 
.A(n_1849),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1825),
.B(n_1383),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1825),
.B(n_1388),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1775),
.B(n_1396),
.Y(n_2028)
);

BUFx12f_ASAP7_75t_L g2029 ( 
.A(n_1743),
.Y(n_2029)
);

BUFx4f_ASAP7_75t_L g2030 ( 
.A(n_1756),
.Y(n_2030)
);

O2A1O1Ixp33_ASAP7_75t_L g2031 ( 
.A1(n_1825),
.A2(n_1046),
.B(n_1056),
.C(n_1023),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1825),
.A2(n_1409),
.B1(n_1419),
.B2(n_1408),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1825),
.B(n_1421),
.Y(n_2033)
);

AO221x2_ASAP7_75t_L g2034 ( 
.A1(n_1740),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.C(n_26),
.Y(n_2034)
);

O2A1O1Ixp33_ASAP7_75t_L g2035 ( 
.A1(n_1825),
.A2(n_1141),
.B(n_1234),
.C(n_1091),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1825),
.B(n_1078),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1775),
.B(n_1079),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1840),
.B(n_1316),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1821),
.A2(n_1083),
.B(n_1082),
.Y(n_2039)
);

OR2x6_ASAP7_75t_L g2040 ( 
.A(n_1858),
.B(n_1342),
.Y(n_2040)
);

O2A1O1Ixp33_ASAP7_75t_L g2041 ( 
.A1(n_1825),
.A2(n_1404),
.B(n_1416),
.C(n_1345),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1827),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1821),
.A2(n_1090),
.B(n_1089),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1737),
.Y(n_2044)
);

AOI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1839),
.A2(n_1425),
.B(n_1121),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1840),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1825),
.B(n_1096),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1821),
.A2(n_1113),
.B(n_1105),
.Y(n_2048)
);

OAI21xp33_ASAP7_75t_SL g2049 ( 
.A1(n_1777),
.A2(n_28),
.B(n_25),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1737),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1775),
.B(n_1118),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1840),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1894),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_2042),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_2045),
.A2(n_1121),
.B(n_1080),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_1923),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1885),
.B(n_23),
.Y(n_2057)
);

AOI22x1_ASAP7_75t_L g2058 ( 
.A1(n_1970),
.A2(n_1132),
.B1(n_1138),
.B2(n_1136),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1995),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1901),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1877),
.Y(n_2061)
);

BUFx3_ASAP7_75t_L g2062 ( 
.A(n_2030),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_2029),
.Y(n_2063)
);

AO21x2_ASAP7_75t_L g2064 ( 
.A1(n_1878),
.A2(n_1121),
.B(n_1080),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_2046),
.B(n_1116),
.Y(n_2065)
);

BUFx3_ASAP7_75t_L g2066 ( 
.A(n_2046),
.Y(n_2066)
);

BUFx12f_ASAP7_75t_L g2067 ( 
.A(n_1930),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_2027),
.B(n_2033),
.Y(n_2068)
);

AOI22x1_ASAP7_75t_L g2069 ( 
.A1(n_1908),
.A2(n_1140),
.B1(n_1148),
.B2(n_1142),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_2052),
.Y(n_2070)
);

BUFx8_ASAP7_75t_L g2071 ( 
.A(n_1993),
.Y(n_2071)
);

OR2x6_ASAP7_75t_L g2072 ( 
.A(n_1922),
.B(n_1905),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1965),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1891),
.Y(n_2074)
);

AO21x2_ASAP7_75t_L g2075 ( 
.A1(n_1935),
.A2(n_1121),
.B(n_1080),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_1911),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1907),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1966),
.A2(n_1121),
.B(n_1080),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_2036),
.A2(n_1171),
.B(n_1169),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1907),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1942),
.Y(n_2081)
);

NAND2x1p5_ASAP7_75t_L g2082 ( 
.A(n_2007),
.B(n_1116),
.Y(n_2082)
);

OAI21x1_ASAP7_75t_L g2083 ( 
.A1(n_1982),
.A2(n_1080),
.B(n_660),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_1948),
.B(n_1116),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1881),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1942),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1874),
.B(n_2026),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1882),
.Y(n_2088)
);

INVx8_ASAP7_75t_L g2089 ( 
.A(n_2040),
.Y(n_2089)
);

OA21x2_ASAP7_75t_L g2090 ( 
.A1(n_1876),
.A2(n_1183),
.B(n_1181),
.Y(n_2090)
);

AO21x2_ASAP7_75t_L g2091 ( 
.A1(n_1915),
.A2(n_1344),
.B(n_1288),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2001),
.A2(n_2006),
.B(n_1957),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1952),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_1981),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1895),
.Y(n_2095)
);

OAI21x1_ASAP7_75t_L g2096 ( 
.A1(n_2017),
.A2(n_661),
.B(n_657),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_2014),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1887),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1897),
.Y(n_2099)
);

AO21x2_ASAP7_75t_L g2100 ( 
.A1(n_1909),
.A2(n_1344),
.B(n_1288),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1904),
.Y(n_2101)
);

AOI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1912),
.A2(n_1344),
.B(n_1288),
.Y(n_2102)
);

BUFx8_ASAP7_75t_SL g2103 ( 
.A(n_2021),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_1899),
.A2(n_664),
.B(n_663),
.Y(n_2104)
);

CKINVDCx11_ASAP7_75t_R g2105 ( 
.A(n_1934),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1900),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_SL g2107 ( 
.A1(n_1988),
.A2(n_28),
.B(n_29),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_1906),
.A2(n_666),
.B(n_665),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1910),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1927),
.Y(n_2110)
);

NAND2x1p5_ASAP7_75t_L g2111 ( 
.A(n_1983),
.B(n_1381),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1917),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_2014),
.Y(n_2113)
);

CKINVDCx20_ASAP7_75t_R g2114 ( 
.A(n_2022),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1932),
.Y(n_2115)
);

INVx6_ASAP7_75t_L g2116 ( 
.A(n_1898),
.Y(n_2116)
);

OAI21x1_ASAP7_75t_L g2117 ( 
.A1(n_1920),
.A2(n_668),
.B(n_667),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1886),
.B(n_1377),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1926),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_2012),
.A2(n_670),
.B(n_669),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1933),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_1937),
.A2(n_672),
.B(n_671),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1925),
.B(n_30),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_1945),
.A2(n_674),
.B(n_673),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_2005),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_2040),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_2016),
.Y(n_2127)
);

CKINVDCx20_ASAP7_75t_R g2128 ( 
.A(n_1973),
.Y(n_2128)
);

AO21x2_ASAP7_75t_L g2129 ( 
.A1(n_1914),
.A2(n_1381),
.B(n_679),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_1946),
.A2(n_680),
.B(n_678),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_1996),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2011),
.A2(n_683),
.B(n_681),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_2016),
.Y(n_2133)
);

OAI21x1_ASAP7_75t_L g2134 ( 
.A1(n_1954),
.A2(n_688),
.B(n_686),
.Y(n_2134)
);

INVx1_ASAP7_75t_SL g2135 ( 
.A(n_1979),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2044),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_2038),
.B(n_30),
.Y(n_2137)
);

AO21x2_ASAP7_75t_L g2138 ( 
.A1(n_2047),
.A2(n_1381),
.B(n_691),
.Y(n_2138)
);

AOI22x1_ASAP7_75t_L g2139 ( 
.A1(n_1928),
.A2(n_1195),
.B1(n_1206),
.B2(n_1193),
.Y(n_2139)
);

OAI21x1_ASAP7_75t_L g2140 ( 
.A1(n_2050),
.A2(n_692),
.B(n_690),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2034),
.A2(n_1221),
.B1(n_1227),
.B2(n_1214),
.Y(n_2141)
);

OAI21x1_ASAP7_75t_L g2142 ( 
.A1(n_1994),
.A2(n_696),
.B(n_693),
.Y(n_2142)
);

INVxp67_ASAP7_75t_SL g2143 ( 
.A(n_1896),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_2031),
.A2(n_698),
.B(n_697),
.Y(n_2144)
);

CKINVDCx16_ASAP7_75t_R g2145 ( 
.A(n_1875),
.Y(n_2145)
);

BUFx2_ASAP7_75t_L g2146 ( 
.A(n_1960),
.Y(n_2146)
);

BUFx12f_ASAP7_75t_L g2147 ( 
.A(n_1962),
.Y(n_2147)
);

AO21x2_ASAP7_75t_L g2148 ( 
.A1(n_1883),
.A2(n_701),
.B(n_699),
.Y(n_2148)
);

INVx6_ASAP7_75t_L g2149 ( 
.A(n_1939),
.Y(n_2149)
);

INVx2_ASAP7_75t_SL g2150 ( 
.A(n_1950),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1980),
.Y(n_2151)
);

NAND2x1p5_ASAP7_75t_L g2152 ( 
.A(n_2020),
.B(n_702),
.Y(n_2152)
);

AO21x2_ASAP7_75t_L g2153 ( 
.A1(n_1888),
.A2(n_1893),
.B(n_1943),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_2019),
.Y(n_2154)
);

AO21x2_ASAP7_75t_L g2155 ( 
.A1(n_1964),
.A2(n_705),
.B(n_704),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1984),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2035),
.A2(n_709),
.B(n_707),
.Y(n_2157)
);

AO21x2_ASAP7_75t_L g2158 ( 
.A1(n_1929),
.A2(n_711),
.B(n_710),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1956),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1976),
.A2(n_1242),
.B1(n_1256),
.B2(n_1231),
.Y(n_2160)
);

AO21x2_ASAP7_75t_L g2161 ( 
.A1(n_1890),
.A2(n_714),
.B(n_712),
.Y(n_2161)
);

BUFx2_ASAP7_75t_SL g2162 ( 
.A(n_1892),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1958),
.B(n_1968),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1884),
.B(n_1902),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1936),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1924),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1941),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_1972),
.A2(n_1424),
.B(n_1422),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_2024),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_2020),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2028),
.B(n_1992),
.Y(n_2171)
);

AO21x2_ASAP7_75t_L g2172 ( 
.A1(n_1903),
.A2(n_716),
.B(n_715),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1953),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1949),
.B(n_1264),
.Y(n_2174)
);

INVx8_ASAP7_75t_L g2175 ( 
.A(n_2013),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1879),
.A2(n_1269),
.B(n_1265),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1986),
.B(n_32),
.Y(n_2177)
);

AO21x2_ASAP7_75t_L g2178 ( 
.A1(n_1880),
.A2(n_718),
.B(n_717),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1955),
.Y(n_2179)
);

OAI21xp33_ASAP7_75t_L g2180 ( 
.A1(n_2032),
.A2(n_1276),
.B(n_1271),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1977),
.Y(n_2181)
);

AO21x2_ASAP7_75t_L g2182 ( 
.A1(n_2039),
.A2(n_721),
.B(n_720),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1916),
.B(n_1978),
.Y(n_2183)
);

AO21x2_ASAP7_75t_L g2184 ( 
.A1(n_2043),
.A2(n_723),
.B(n_722),
.Y(n_2184)
);

OAI21x1_ASAP7_75t_L g2185 ( 
.A1(n_2041),
.A2(n_725),
.B(n_724),
.Y(n_2185)
);

OAI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_2048),
.A2(n_1279),
.B(n_1277),
.Y(n_2186)
);

AO21x2_ASAP7_75t_L g2187 ( 
.A1(n_1998),
.A2(n_727),
.B(n_726),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_1940),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1944),
.Y(n_2189)
);

BUFx8_ASAP7_75t_L g2190 ( 
.A(n_2025),
.Y(n_2190)
);

NAND2x1p5_ASAP7_75t_L g2191 ( 
.A(n_2037),
.B(n_730),
.Y(n_2191)
);

INVx3_ASAP7_75t_L g2192 ( 
.A(n_1975),
.Y(n_2192)
);

BUFx4_ASAP7_75t_SL g2193 ( 
.A(n_1985),
.Y(n_2193)
);

HB1xp67_ASAP7_75t_L g2194 ( 
.A(n_2056),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2061),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2062),
.Y(n_2196)
);

CKINVDCx20_ASAP7_75t_R g2197 ( 
.A(n_2085),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2059),
.Y(n_2198)
);

CKINVDCx14_ASAP7_75t_R g2199 ( 
.A(n_2105),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_2067),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_2066),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2088),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2068),
.A2(n_1918),
.B1(n_1967),
.B2(n_1963),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2167),
.B(n_1919),
.Y(n_2204)
);

CKINVDCx9p33_ASAP7_75t_R g2205 ( 
.A(n_2053),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_2073),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_2080),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2060),
.Y(n_2208)
);

NAND2x1p5_ASAP7_75t_L g2209 ( 
.A(n_2070),
.B(n_2051),
.Y(n_2209)
);

AOI21x1_ASAP7_75t_L g2210 ( 
.A1(n_2102),
.A2(n_2002),
.B(n_1961),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_2086),
.Y(n_2211)
);

OAI21x1_ASAP7_75t_L g2212 ( 
.A1(n_2055),
.A2(n_1889),
.B(n_1997),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_2081),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2165),
.B(n_1951),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_2081),
.Y(n_2215)
);

INVxp67_ASAP7_75t_SL g2216 ( 
.A(n_2143),
.Y(n_2216)
);

NAND2x1p5_ASAP7_75t_L g2217 ( 
.A(n_2054),
.B(n_1913),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2098),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2089),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2174),
.A2(n_1959),
.B1(n_1969),
.B2(n_1931),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2109),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2163),
.B(n_1990),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2146),
.B(n_2000),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2112),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2094),
.Y(n_2225)
);

AOI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2183),
.A2(n_1947),
.B1(n_2023),
.B2(n_2003),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_2116),
.Y(n_2227)
);

OAI21x1_ASAP7_75t_L g2228 ( 
.A1(n_2078),
.A2(n_2004),
.B(n_1987),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2125),
.B(n_1938),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2137),
.B(n_1921),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2177),
.A2(n_1989),
.B1(n_2018),
.B2(n_2008),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2087),
.B(n_1974),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2145),
.B(n_2009),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2131),
.B(n_1991),
.Y(n_2234)
);

NAND2x1p5_ASAP7_75t_L g2235 ( 
.A(n_2093),
.B(n_2015),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2074),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2114),
.A2(n_2049),
.B1(n_1282),
.B2(n_1285),
.Y(n_2237)
);

BUFx3_ASAP7_75t_L g2238 ( 
.A(n_2125),
.Y(n_2238)
);

BUFx10_ASAP7_75t_L g2239 ( 
.A(n_2171),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2095),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_2071),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2150),
.B(n_1971),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2101),
.Y(n_2243)
);

NAND2x1p5_ASAP7_75t_L g2244 ( 
.A(n_2127),
.B(n_1999),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2149),
.A2(n_2010),
.B1(n_1286),
.B2(n_1292),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_SL g2246 ( 
.A1(n_2089),
.A2(n_1337),
.B1(n_1384),
.B2(n_1303),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2057),
.B(n_32),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2079),
.A2(n_1294),
.B(n_1281),
.Y(n_2248)
);

INVx5_ASAP7_75t_L g2249 ( 
.A(n_2065),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2141),
.A2(n_1306),
.B1(n_1314),
.B2(n_1305),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_SL g2251 ( 
.A1(n_2189),
.A2(n_1385),
.B1(n_1336),
.B2(n_1330),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2119),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2147),
.A2(n_1331),
.B1(n_1353),
.B2(n_1329),
.Y(n_2253)
);

BUFx2_ASAP7_75t_L g2254 ( 
.A(n_2128),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2099),
.B(n_33),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2136),
.Y(n_2256)
);

OAI21x1_ASAP7_75t_L g2257 ( 
.A1(n_2083),
.A2(n_734),
.B(n_731),
.Y(n_2257)
);

INVx6_ASAP7_75t_L g2258 ( 
.A(n_2190),
.Y(n_2258)
);

CKINVDCx11_ASAP7_75t_R g2259 ( 
.A(n_2072),
.Y(n_2259)
);

AOI21x1_ASAP7_75t_L g2260 ( 
.A1(n_2181),
.A2(n_1363),
.B(n_1355),
.Y(n_2260)
);

BUFx12f_ASAP7_75t_L g2261 ( 
.A(n_2126),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2154),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2110),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2156),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2115),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_SL g2266 ( 
.A1(n_2188),
.A2(n_1394),
.B1(n_1372),
.B2(n_1374),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2121),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2151),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2169),
.A2(n_1382),
.B1(n_1391),
.B2(n_1368),
.Y(n_2269)
);

BUFx8_ASAP7_75t_L g2270 ( 
.A(n_2127),
.Y(n_2270)
);

INVxp33_ASAP7_75t_SL g2271 ( 
.A(n_2193),
.Y(n_2271)
);

NAND2x1p5_ASAP7_75t_L g2272 ( 
.A(n_2133),
.B(n_735),
.Y(n_2272)
);

BUFx12f_ASAP7_75t_L g2273 ( 
.A(n_2133),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2175),
.A2(n_1401),
.B1(n_1412),
.B2(n_1400),
.Y(n_2274)
);

INVx1_ASAP7_75t_SL g2275 ( 
.A(n_2135),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2092),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2123),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2173),
.Y(n_2278)
);

AOI21x1_ASAP7_75t_L g2279 ( 
.A1(n_2090),
.A2(n_1420),
.B(n_738),
.Y(n_2279)
);

OR2x6_ASAP7_75t_L g2280 ( 
.A(n_2175),
.B(n_33),
.Y(n_2280)
);

AOI22xp33_ASAP7_75t_L g2281 ( 
.A1(n_2153),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2170),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_SL g2283 ( 
.A(n_2170),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2192),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2075),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2134),
.A2(n_739),
.B(n_736),
.Y(n_2286)
);

NAND2x1p5_ASAP7_75t_L g2287 ( 
.A(n_2076),
.B(n_2077),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_2176),
.A2(n_2164),
.B1(n_2180),
.B2(n_2118),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2097),
.B(n_35),
.Y(n_2289)
);

OA21x2_ASAP7_75t_L g2290 ( 
.A1(n_2144),
.A2(n_741),
.B(n_740),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2162),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2103),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2179),
.B(n_36),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2113),
.Y(n_2294)
);

OAI21x1_ASAP7_75t_L g2295 ( 
.A1(n_2140),
.A2(n_2124),
.B(n_2122),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2187),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2160),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2063),
.B(n_38),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2106),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2166),
.Y(n_2300)
);

OA21x2_ASAP7_75t_L g2301 ( 
.A1(n_2157),
.A2(n_743),
.B(n_742),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2082),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2148),
.Y(n_2303)
);

BUFx2_ASAP7_75t_L g2304 ( 
.A(n_2159),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2158),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2058),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2084),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2107),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2186),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2111),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_2310)
);

AO21x2_ASAP7_75t_L g2311 ( 
.A1(n_2064),
.A2(n_745),
.B(n_744),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2152),
.Y(n_2312)
);

INVx3_ASAP7_75t_SL g2313 ( 
.A(n_2191),
.Y(n_2313)
);

INVx11_ASAP7_75t_L g2314 ( 
.A(n_2130),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_2168),
.Y(n_2315)
);

NAND2x1p5_ASAP7_75t_L g2316 ( 
.A(n_2096),
.B(n_749),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2117),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2129),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2139),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2132),
.Y(n_2320)
);

NAND3xp33_ASAP7_75t_L g2321 ( 
.A(n_2069),
.B(n_45),
.C(n_47),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2120),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2142),
.Y(n_2323)
);

OA21x2_ASAP7_75t_L g2324 ( 
.A1(n_2185),
.A2(n_752),
.B(n_751),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2161),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2172),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2104),
.Y(n_2327)
);

INVx2_ASAP7_75t_SL g2328 ( 
.A(n_2178),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2182),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2091),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2184),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2108),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2155),
.Y(n_2333)
);

INVx4_ASAP7_75t_SL g2334 ( 
.A(n_2138),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2100),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2059),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2055),
.A2(n_755),
.B(n_754),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2061),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2163),
.B(n_48),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2059),
.Y(n_2340)
);

INVxp33_ASAP7_75t_L g2341 ( 
.A(n_2053),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2068),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_2342)
);

NAND2x1p5_ASAP7_75t_L g2343 ( 
.A(n_2062),
.B(n_756),
.Y(n_2343)
);

INVx2_ASAP7_75t_SL g2344 ( 
.A(n_2062),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2062),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2195),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2202),
.Y(n_2347)
);

NAND2xp33_ASAP7_75t_R g2348 ( 
.A(n_2271),
.B(n_950),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_2241),
.Y(n_2349)
);

BUFx3_ASAP7_75t_L g2350 ( 
.A(n_2270),
.Y(n_2350)
);

NOR3xp33_ASAP7_75t_SL g2351 ( 
.A(n_2292),
.B(n_50),
.C(n_53),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2218),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2221),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2345),
.Y(n_2354)
);

OAI21xp33_ASAP7_75t_L g2355 ( 
.A1(n_2203),
.A2(n_54),
.B(n_56),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_SL g2356 ( 
.A1(n_2220),
.A2(n_2237),
.B1(n_2309),
.B2(n_2233),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2230),
.B(n_54),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_SL g2358 ( 
.A(n_2298),
.B(n_56),
.C(n_57),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2224),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_2249),
.B(n_57),
.Y(n_2360)
);

BUFx3_ASAP7_75t_L g2361 ( 
.A(n_2345),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2194),
.B(n_58),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_SL g2363 ( 
.A1(n_2342),
.A2(n_58),
.B(n_59),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_2197),
.Y(n_2364)
);

OAI221xp5_ASAP7_75t_L g2365 ( 
.A1(n_2293),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.C(n_63),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2223),
.B(n_60),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_R g2367 ( 
.A(n_2306),
.B(n_757),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2216),
.B(n_61),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2225),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2198),
.Y(n_2370)
);

OR2x6_ASAP7_75t_L g2371 ( 
.A(n_2219),
.B(n_758),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_2208),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2338),
.Y(n_2373)
);

BUFx2_ASAP7_75t_L g2374 ( 
.A(n_2205),
.Y(n_2374)
);

XNOR2xp5_ASAP7_75t_L g2375 ( 
.A(n_2254),
.B(n_63),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2252),
.Y(n_2376)
);

CKINVDCx20_ASAP7_75t_R g2377 ( 
.A(n_2199),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2339),
.B(n_64),
.Y(n_2378)
);

OA21x2_ASAP7_75t_L g2379 ( 
.A1(n_2295),
.A2(n_66),
.B(n_67),
.Y(n_2379)
);

INVx8_ASAP7_75t_L g2380 ( 
.A(n_2283),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2226),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2381)
);

NAND3xp33_ASAP7_75t_SL g2382 ( 
.A(n_2231),
.B(n_68),
.C(n_69),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2256),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2255),
.B(n_2247),
.Y(n_2384)
);

INVx2_ASAP7_75t_SL g2385 ( 
.A(n_2207),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2249),
.B(n_70),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2264),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_R g2388 ( 
.A(n_2206),
.B(n_953),
.Y(n_2388)
);

AO21x2_ASAP7_75t_L g2389 ( 
.A1(n_2325),
.A2(n_761),
.B(n_759),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2232),
.A2(n_71),
.B(n_72),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2280),
.B(n_72),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2336),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2280),
.B(n_73),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2268),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_2259),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2204),
.B(n_2275),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2340),
.Y(n_2397)
);

OR2x4_ASAP7_75t_L g2398 ( 
.A(n_2213),
.B(n_74),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2277),
.B(n_74),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2261),
.Y(n_2400)
);

CKINVDCx8_ASAP7_75t_R g2401 ( 
.A(n_2262),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_R g2402 ( 
.A(n_2273),
.B(n_762),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2341),
.B(n_2213),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2211),
.Y(n_2404)
);

OR2x6_ASAP7_75t_L g2405 ( 
.A(n_2258),
.B(n_2344),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2215),
.B(n_2201),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2214),
.B(n_75),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2236),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2240),
.Y(n_2409)
);

NAND2xp33_ASAP7_75t_SL g2410 ( 
.A(n_2313),
.B(n_75),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2243),
.Y(n_2411)
);

OAI21xp33_ASAP7_75t_L g2412 ( 
.A1(n_2297),
.A2(n_76),
.B(n_77),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2215),
.B(n_76),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2263),
.Y(n_2414)
);

AO31x2_ASAP7_75t_L g2415 ( 
.A1(n_2318),
.A2(n_764),
.A3(n_766),
.B(n_763),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2282),
.B(n_77),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2265),
.Y(n_2417)
);

OAI21xp33_ASAP7_75t_L g2418 ( 
.A1(n_2281),
.A2(n_78),
.B(n_79),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2234),
.B(n_78),
.Y(n_2419)
);

OR2x2_ASAP7_75t_L g2420 ( 
.A(n_2278),
.B(n_79),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2267),
.Y(n_2421)
);

OR2x6_ASAP7_75t_L g2422 ( 
.A(n_2196),
.B(n_767),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2284),
.Y(n_2423)
);

OAI22xp33_ASAP7_75t_SL g2424 ( 
.A1(n_2242),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_2238),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2294),
.Y(n_2426)
);

NAND2xp33_ASAP7_75t_R g2427 ( 
.A(n_2222),
.B(n_955),
.Y(n_2427)
);

BUFx6f_ASAP7_75t_L g2428 ( 
.A(n_2304),
.Y(n_2428)
);

OR2x6_ASAP7_75t_L g2429 ( 
.A(n_2343),
.B(n_768),
.Y(n_2429)
);

AO31x2_ASAP7_75t_L g2430 ( 
.A1(n_2305),
.A2(n_770),
.A3(n_772),
.B(n_769),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_R g2431 ( 
.A(n_2200),
.B(n_774),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2227),
.B(n_80),
.Y(n_2432)
);

CKINVDCx20_ASAP7_75t_R g2433 ( 
.A(n_2300),
.Y(n_2433)
);

CKINVDCx16_ASAP7_75t_R g2434 ( 
.A(n_2239),
.Y(n_2434)
);

INVx4_ASAP7_75t_SL g2435 ( 
.A(n_2229),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_2287),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_2312),
.B(n_81),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2235),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2299),
.B(n_2289),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_R g2440 ( 
.A(n_2291),
.B(n_775),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2276),
.Y(n_2441)
);

NAND2xp33_ASAP7_75t_SL g2442 ( 
.A(n_2288),
.B(n_82),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2209),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2308),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_2217),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2248),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2210),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2269),
.B(n_83),
.Y(n_2448)
);

NOR3xp33_ASAP7_75t_SL g2449 ( 
.A(n_2321),
.B(n_2319),
.C(n_2250),
.Y(n_2449)
);

AOI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2266),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_2450)
);

NOR3xp33_ASAP7_75t_SL g2451 ( 
.A(n_2317),
.B(n_86),
.C(n_87),
.Y(n_2451)
);

NAND2xp33_ASAP7_75t_SL g2452 ( 
.A(n_2310),
.B(n_2274),
.Y(n_2452)
);

INVxp67_ASAP7_75t_L g2453 ( 
.A(n_2302),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2307),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_R g2455 ( 
.A(n_2260),
.B(n_776),
.Y(n_2455)
);

INVx4_ASAP7_75t_L g2456 ( 
.A(n_2272),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2322),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2244),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2253),
.B(n_88),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2279),
.Y(n_2460)
);

NOR2x1_ASAP7_75t_L g2461 ( 
.A(n_2326),
.B(n_88),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2245),
.B(n_89),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2246),
.B(n_89),
.Y(n_2463)
);

INVxp33_ASAP7_75t_SL g2464 ( 
.A(n_2251),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2285),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2315),
.B(n_90),
.Y(n_2466)
);

BUFx3_ASAP7_75t_L g2467 ( 
.A(n_2228),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2334),
.B(n_90),
.Y(n_2468)
);

NAND2xp33_ASAP7_75t_SL g2469 ( 
.A(n_2323),
.B(n_91),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2314),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2330),
.B(n_91),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2334),
.B(n_92),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_2320),
.B(n_93),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2316),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2257),
.B(n_93),
.Y(n_2475)
);

INVx8_ASAP7_75t_L g2476 ( 
.A(n_2323),
.Y(n_2476)
);

OAI21x1_ASAP7_75t_L g2477 ( 
.A1(n_2333),
.A2(n_2303),
.B(n_2329),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2311),
.B(n_94),
.Y(n_2478)
);

OR2x6_ASAP7_75t_L g2479 ( 
.A(n_2286),
.B(n_778),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2327),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_2332),
.Y(n_2481)
);

NAND3xp33_ASAP7_75t_SL g2482 ( 
.A(n_2296),
.B(n_94),
.C(n_95),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2331),
.A2(n_2328),
.B1(n_2335),
.B2(n_2290),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_R g2484 ( 
.A(n_2212),
.B(n_780),
.Y(n_2484)
);

CKINVDCx20_ASAP7_75t_R g2485 ( 
.A(n_2301),
.Y(n_2485)
);

INVx1_ASAP7_75t_SL g2486 ( 
.A(n_2324),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2370),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2404),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2372),
.B(n_2435),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2396),
.B(n_95),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2346),
.Y(n_2491)
);

NOR2x1_ASAP7_75t_L g2492 ( 
.A(n_2368),
.B(n_2337),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2384),
.B(n_2357),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2392),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_2369),
.B(n_2347),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2364),
.B(n_96),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2352),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2366),
.B(n_96),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2397),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2353),
.Y(n_2500)
);

OR2x2_ASAP7_75t_L g2501 ( 
.A(n_2359),
.B(n_97),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2481),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2378),
.B(n_97),
.Y(n_2503)
);

HB1xp67_ASAP7_75t_L g2504 ( 
.A(n_2373),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2403),
.B(n_98),
.Y(n_2505)
);

AOI221xp5_ASAP7_75t_L g2506 ( 
.A1(n_2365),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.C(n_101),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2404),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2408),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2376),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2383),
.B(n_2387),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2394),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2457),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2423),
.B(n_99),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2419),
.B(n_2420),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2374),
.B(n_100),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2409),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2467),
.Y(n_2517)
);

OR2x2_ASAP7_75t_L g2518 ( 
.A(n_2426),
.B(n_102),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2413),
.B(n_102),
.Y(n_2519)
);

BUFx2_ASAP7_75t_SL g2520 ( 
.A(n_2433),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2480),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2444),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2473),
.B(n_2406),
.Y(n_2523)
);

NOR2x1_ASAP7_75t_SL g2524 ( 
.A(n_2429),
.B(n_103),
.Y(n_2524)
);

OR2x2_ASAP7_75t_L g2525 ( 
.A(n_2362),
.B(n_103),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2416),
.B(n_104),
.Y(n_2526)
);

BUFx2_ASAP7_75t_L g2527 ( 
.A(n_2485),
.Y(n_2527)
);

HB1xp67_ASAP7_75t_L g2528 ( 
.A(n_2438),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2428),
.B(n_104),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2411),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2407),
.B(n_105),
.Y(n_2531)
);

INVx3_ASAP7_75t_L g2532 ( 
.A(n_2401),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2414),
.Y(n_2533)
);

BUFx2_ASAP7_75t_L g2534 ( 
.A(n_2476),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2428),
.B(n_105),
.Y(n_2535)
);

CKINVDCx11_ASAP7_75t_R g2536 ( 
.A(n_2377),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2391),
.B(n_2393),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2466),
.B(n_2356),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2417),
.Y(n_2539)
);

HB1xp67_ASAP7_75t_L g2540 ( 
.A(n_2458),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2421),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2454),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2439),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2441),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2361),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2447),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2465),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2472),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2461),
.Y(n_2549)
);

HB1xp67_ASAP7_75t_L g2550 ( 
.A(n_2470),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2399),
.B(n_106),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2443),
.B(n_106),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2445),
.B(n_107),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2453),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2468),
.Y(n_2555)
);

OAI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2363),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2385),
.B(n_108),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2476),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2478),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2379),
.Y(n_2560)
);

INVx4_ASAP7_75t_L g2561 ( 
.A(n_2380),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2477),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2415),
.Y(n_2563)
);

INVx4_ASAP7_75t_R g2564 ( 
.A(n_2350),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_2474),
.Y(n_2565)
);

INVxp67_ASAP7_75t_SL g2566 ( 
.A(n_2460),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_2380),
.B(n_781),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2358),
.B(n_109),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2475),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2432),
.B(n_110),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2415),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2430),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2463),
.B(n_110),
.Y(n_2573)
);

HB1xp67_ASAP7_75t_L g2574 ( 
.A(n_2486),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2430),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2435),
.B(n_782),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2360),
.B(n_112),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2543),
.B(n_2355),
.Y(n_2578)
);

AND2x4_ASAP7_75t_SL g2579 ( 
.A(n_2532),
.B(n_2405),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2508),
.Y(n_2580)
);

INVx2_ASAP7_75t_SL g2581 ( 
.A(n_2488),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2527),
.B(n_2405),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2500),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2527),
.B(n_2354),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2504),
.Y(n_2585)
);

HB1xp67_ASAP7_75t_L g2586 ( 
.A(n_2502),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2523),
.B(n_2425),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2538),
.A2(n_2452),
.B1(n_2442),
.B2(n_2464),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2545),
.Y(n_2589)
);

BUFx2_ASAP7_75t_SL g2590 ( 
.A(n_2561),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2559),
.B(n_2451),
.Y(n_2591)
);

OR2x2_ASAP7_75t_L g2592 ( 
.A(n_2495),
.B(n_2434),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2493),
.B(n_2386),
.Y(n_2593)
);

OAI21xp5_ASAP7_75t_SL g2594 ( 
.A1(n_2556),
.A2(n_2382),
.B(n_2375),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2537),
.B(n_2422),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2520),
.B(n_2395),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2510),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2522),
.Y(n_2598)
);

NOR2x1p5_ASAP7_75t_L g2599 ( 
.A(n_2549),
.B(n_2400),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2491),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2502),
.B(n_2422),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2497),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2516),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2550),
.B(n_2371),
.Y(n_2604)
);

OA21x2_ASAP7_75t_L g2605 ( 
.A1(n_2560),
.A2(n_2563),
.B(n_2571),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2530),
.Y(n_2606)
);

NOR3xp33_ASAP7_75t_L g2607 ( 
.A(n_2506),
.B(n_2446),
.C(n_2412),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2505),
.B(n_2371),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2536),
.B(n_2398),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2542),
.B(n_2390),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_SL g2611 ( 
.A(n_2534),
.B(n_2431),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2509),
.B(n_2424),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2511),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2515),
.B(n_2529),
.Y(n_2614)
);

NOR2x1_ASAP7_75t_R g2615 ( 
.A(n_2489),
.B(n_2349),
.Y(n_2615)
);

OAI21xp5_ASAP7_75t_SL g2616 ( 
.A1(n_2568),
.A2(n_2450),
.B(n_2381),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2512),
.Y(n_2617)
);

OAI21xp5_ASAP7_75t_SL g2618 ( 
.A1(n_2496),
.A2(n_2462),
.B(n_2448),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2535),
.B(n_2514),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2548),
.B(n_2554),
.Y(n_2620)
);

INVx2_ASAP7_75t_SL g2621 ( 
.A(n_2507),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2569),
.B(n_2565),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2521),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2501),
.B(n_2351),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2519),
.B(n_2436),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2517),
.B(n_2456),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2574),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2539),
.Y(n_2628)
);

OAI221xp5_ASAP7_75t_L g2629 ( 
.A1(n_2531),
.A2(n_2410),
.B1(n_2459),
.B2(n_2418),
.C(n_2367),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2546),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2498),
.B(n_2440),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2517),
.B(n_2429),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2533),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2503),
.B(n_2471),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2541),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2544),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2526),
.B(n_2437),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2555),
.B(n_2479),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2540),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2534),
.B(n_2528),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2487),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2573),
.B(n_2479),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2558),
.B(n_2389),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2552),
.B(n_2402),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2553),
.B(n_2484),
.Y(n_2645)
);

OR2x2_ASAP7_75t_L g2646 ( 
.A(n_2513),
.B(n_2482),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2577),
.B(n_2570),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2494),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2499),
.Y(n_2649)
);

NAND3xp33_ASAP7_75t_L g2650 ( 
.A(n_2551),
.B(n_2449),
.C(n_2469),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2547),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2566),
.Y(n_2652)
);

NOR2x1_ASAP7_75t_L g2653 ( 
.A(n_2518),
.B(n_2388),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2490),
.B(n_112),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2525),
.B(n_2483),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2562),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2492),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2557),
.B(n_2455),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2567),
.B(n_2572),
.Y(n_2659)
);

HB1xp67_ASAP7_75t_L g2660 ( 
.A(n_2575),
.Y(n_2660)
);

HB1xp67_ASAP7_75t_L g2661 ( 
.A(n_2586),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2623),
.Y(n_2662)
);

INVxp67_ASAP7_75t_SL g2663 ( 
.A(n_2657),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2640),
.B(n_2524),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2640),
.B(n_2567),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2627),
.B(n_113),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_2607),
.A2(n_2576),
.B1(n_2427),
.B2(n_2348),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_R g2668 ( 
.A(n_2611),
.B(n_2564),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2582),
.B(n_113),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2583),
.B(n_114),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2580),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2584),
.B(n_2601),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2603),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2653),
.B(n_115),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2606),
.Y(n_2675)
);

INVx1_ASAP7_75t_SL g2676 ( 
.A(n_2579),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2585),
.B(n_2597),
.Y(n_2677)
);

AND2x2_ASAP7_75t_SL g2678 ( 
.A(n_2632),
.B(n_115),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2626),
.Y(n_2679)
);

HB1xp67_ASAP7_75t_L g2680 ( 
.A(n_2622),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2598),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2595),
.B(n_116),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2620),
.B(n_117),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2626),
.B(n_118),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2600),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2592),
.B(n_118),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2619),
.B(n_119),
.Y(n_2687)
);

AND2x4_ASAP7_75t_SL g2688 ( 
.A(n_2587),
.B(n_119),
.Y(n_2688)
);

NOR3xp33_ASAP7_75t_SL g2689 ( 
.A(n_2594),
.B(n_120),
.C(n_121),
.Y(n_2689)
);

INVxp67_ASAP7_75t_L g2690 ( 
.A(n_2639),
.Y(n_2690)
);

AND2x2_ASAP7_75t_SL g2691 ( 
.A(n_2645),
.B(n_120),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2602),
.B(n_121),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2613),
.B(n_122),
.Y(n_2693)
);

AND2x4_ASAP7_75t_SL g2694 ( 
.A(n_2625),
.B(n_123),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2614),
.B(n_123),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2590),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2617),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2628),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2630),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2636),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2642),
.B(n_124),
.Y(n_2701)
);

INVxp67_ASAP7_75t_L g2702 ( 
.A(n_2589),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2610),
.B(n_124),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2659),
.B(n_2638),
.Y(n_2704)
);

AND2x4_ASAP7_75t_L g2705 ( 
.A(n_2599),
.B(n_125),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2633),
.Y(n_2706)
);

INVxp67_ASAP7_75t_L g2707 ( 
.A(n_2621),
.Y(n_2707)
);

NAND2x1p5_ASAP7_75t_L g2708 ( 
.A(n_2581),
.B(n_127),
.Y(n_2708)
);

OR2x2_ASAP7_75t_SL g2709 ( 
.A(n_2591),
.B(n_127),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2635),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2593),
.B(n_128),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2608),
.B(n_128),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2604),
.B(n_129),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2631),
.B(n_129),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2647),
.B(n_130),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2578),
.B(n_130),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2634),
.B(n_131),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2652),
.B(n_131),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2641),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2649),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2612),
.B(n_132),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2655),
.B(n_132),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2646),
.B(n_133),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2648),
.Y(n_2724)
);

NOR2xp67_ASAP7_75t_L g2725 ( 
.A(n_2596),
.B(n_133),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2651),
.Y(n_2726)
);

NOR2x1_ASAP7_75t_L g2727 ( 
.A(n_2650),
.B(n_134),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2658),
.B(n_134),
.Y(n_2728)
);

AND2x2_ASAP7_75t_SL g2729 ( 
.A(n_2644),
.B(n_135),
.Y(n_2729)
);

NAND2xp33_ASAP7_75t_R g2730 ( 
.A(n_2609),
.B(n_136),
.Y(n_2730)
);

HB1xp67_ASAP7_75t_L g2731 ( 
.A(n_2643),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2654),
.B(n_2618),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2637),
.B(n_136),
.Y(n_2733)
);

AND2x4_ASAP7_75t_SL g2734 ( 
.A(n_2615),
.B(n_137),
.Y(n_2734)
);

OR2x6_ASAP7_75t_L g2735 ( 
.A(n_2624),
.B(n_138),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2656),
.B(n_138),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2605),
.B(n_139),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2605),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2616),
.B(n_139),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2588),
.B(n_140),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2660),
.B(n_140),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2629),
.B(n_143),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2586),
.B(n_143),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2586),
.B(n_144),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2623),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2580),
.Y(n_2746)
);

BUFx2_ASAP7_75t_L g2747 ( 
.A(n_2586),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2679),
.B(n_2672),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2738),
.Y(n_2749)
);

OAI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_2739),
.A2(n_2732),
.B1(n_2735),
.B2(n_2722),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_2676),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2680),
.B(n_144),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2737),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2663),
.B(n_145),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2747),
.B(n_145),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2662),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2747),
.B(n_2661),
.Y(n_2757)
);

INVxp67_ASAP7_75t_L g2758 ( 
.A(n_2730),
.Y(n_2758)
);

NAND5xp2_ASAP7_75t_L g2759 ( 
.A(n_2689),
.B(n_148),
.C(n_146),
.D(n_147),
.E(n_149),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2745),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2664),
.B(n_146),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2671),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2681),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2685),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2742),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2690),
.B(n_150),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2727),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_2767)
);

O2A1O1Ixp33_ASAP7_75t_L g2768 ( 
.A1(n_2721),
.A2(n_154),
.B(n_151),
.C(n_153),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2697),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2696),
.B(n_154),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2698),
.Y(n_2771)
);

OAI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2735),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2772)
);

AND2x2_ASAP7_75t_SL g2773 ( 
.A(n_2678),
.B(n_155),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_SL g2774 ( 
.A(n_2729),
.B(n_157),
.Y(n_2774)
);

INVx1_ASAP7_75t_SL g2775 ( 
.A(n_2734),
.Y(n_2775)
);

OR2x2_ASAP7_75t_L g2776 ( 
.A(n_2677),
.B(n_158),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2665),
.B(n_158),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2699),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2731),
.B(n_159),
.Y(n_2779)
);

OA222x2_ASAP7_75t_L g2780 ( 
.A1(n_2740),
.A2(n_161),
.B1(n_164),
.B2(n_159),
.C1(n_160),
.C2(n_162),
.Y(n_2780)
);

INVx3_ASAP7_75t_L g2781 ( 
.A(n_2704),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2684),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2700),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2702),
.B(n_160),
.Y(n_2784)
);

OAI21xp33_ASAP7_75t_L g2785 ( 
.A1(n_2723),
.A2(n_2703),
.B(n_2716),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2710),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2707),
.B(n_164),
.Y(n_2787)
);

NOR2x1p5_ASAP7_75t_SL g2788 ( 
.A(n_2692),
.B(n_165),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2688),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2743),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2668),
.B(n_165),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2705),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2719),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2720),
.Y(n_2794)
);

HB1xp67_ASAP7_75t_L g2795 ( 
.A(n_2744),
.Y(n_2795)
);

INVxp67_ASAP7_75t_SL g2796 ( 
.A(n_2741),
.Y(n_2796)
);

AOI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2667),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.Y(n_2797)
);

INVxp67_ASAP7_75t_L g2798 ( 
.A(n_2666),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2724),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2691),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2683),
.B(n_170),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2726),
.Y(n_2802)
);

O2A1O1Ixp33_ASAP7_75t_SL g2803 ( 
.A1(n_2728),
.A2(n_173),
.B(n_170),
.C(n_172),
.Y(n_2803)
);

OAI21xp33_ASAP7_75t_SL g2804 ( 
.A1(n_2715),
.A2(n_2717),
.B(n_2670),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2673),
.Y(n_2805)
);

NOR2x1p5_ASAP7_75t_SL g2806 ( 
.A(n_2718),
.B(n_172),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2675),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2693),
.B(n_173),
.Y(n_2808)
);

INVx1_ASAP7_75t_SL g2809 ( 
.A(n_2714),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2706),
.B(n_2746),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2736),
.Y(n_2811)
);

INVxp67_ASAP7_75t_L g2812 ( 
.A(n_2725),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2687),
.B(n_174),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2709),
.B(n_174),
.Y(n_2814)
);

NAND3xp33_ASAP7_75t_L g2815 ( 
.A(n_2686),
.B(n_175),
.C(n_176),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2713),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2733),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2712),
.Y(n_2818)
);

AND2x4_ASAP7_75t_L g2819 ( 
.A(n_2701),
.B(n_176),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2695),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2669),
.B(n_177),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2682),
.B(n_177),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2711),
.B(n_178),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2674),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2694),
.B(n_178),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2708),
.B(n_179),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2679),
.B(n_179),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2739),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2679),
.B(n_181),
.Y(n_2829)
);

INVx3_ASAP7_75t_SL g2830 ( 
.A(n_2696),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2676),
.Y(n_2831)
);

OA222x2_ASAP7_75t_L g2832 ( 
.A1(n_2735),
.A2(n_185),
.B1(n_187),
.B2(n_182),
.C1(n_184),
.C2(n_186),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2662),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2662),
.Y(n_2834)
);

INVx4_ASAP7_75t_L g2835 ( 
.A(n_2696),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2680),
.B(n_185),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2738),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2662),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2679),
.B(n_187),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2662),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2662),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2662),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2679),
.B(n_188),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2679),
.B(n_188),
.Y(n_2844)
);

AOI32xp33_ASAP7_75t_L g2845 ( 
.A1(n_2727),
.A2(n_191),
.A3(n_189),
.B1(n_190),
.B2(n_194),
.Y(n_2845)
);

HB1xp67_ASAP7_75t_L g2846 ( 
.A(n_2747),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2662),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2662),
.Y(n_2848)
);

AND2x4_ASAP7_75t_SL g2849 ( 
.A(n_2665),
.B(n_190),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2662),
.Y(n_2850)
);

INVx1_ASAP7_75t_SL g2851 ( 
.A(n_2676),
.Y(n_2851)
);

NAND4xp75_ASAP7_75t_L g2852 ( 
.A(n_2727),
.B(n_195),
.C(n_191),
.D(n_194),
.Y(n_2852)
);

AOI32xp33_ASAP7_75t_L g2853 ( 
.A1(n_2727),
.A2(n_198),
.A3(n_195),
.B1(n_196),
.B2(n_199),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2662),
.Y(n_2854)
);

AOI211xp5_ASAP7_75t_L g2855 ( 
.A1(n_2739),
.A2(n_207),
.B(n_215),
.C(n_196),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2680),
.B(n_198),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2662),
.Y(n_2857)
);

OAI21xp33_ASAP7_75t_L g2858 ( 
.A1(n_2845),
.A2(n_199),
.B(n_200),
.Y(n_2858)
);

A2O1A1Ixp33_ASAP7_75t_L g2859 ( 
.A1(n_2814),
.A2(n_211),
.B(n_220),
.C(n_200),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2751),
.B(n_2831),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2763),
.Y(n_2861)
);

AOI211xp5_ASAP7_75t_SL g2862 ( 
.A1(n_2772),
.A2(n_204),
.B(n_201),
.C(n_203),
.Y(n_2862)
);

AOI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2774),
.A2(n_208),
.B1(n_204),
.B2(n_205),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2796),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2764),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2753),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2769),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2749),
.Y(n_2868)
);

INVxp67_ASAP7_75t_L g2869 ( 
.A(n_2756),
.Y(n_2869)
);

AOI221xp5_ASAP7_75t_L g2870 ( 
.A1(n_2768),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.C(n_214),
.Y(n_2870)
);

OAI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2804),
.A2(n_212),
.B(n_214),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2771),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2760),
.B(n_2833),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2778),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2783),
.Y(n_2875)
);

AO21x1_ASAP7_75t_L g2876 ( 
.A1(n_2750),
.A2(n_216),
.B(n_217),
.Y(n_2876)
);

AOI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2773),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2877)
);

OAI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2767),
.A2(n_218),
.B(n_219),
.Y(n_2878)
);

INVx1_ASAP7_75t_SL g2879 ( 
.A(n_2830),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2800),
.A2(n_222),
.B1(n_219),
.B2(n_221),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2834),
.Y(n_2881)
);

OAI21xp33_ASAP7_75t_SL g2882 ( 
.A1(n_2757),
.A2(n_221),
.B(n_222),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2797),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2838),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2840),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2758),
.A2(n_227),
.B1(n_224),
.B2(n_226),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2828),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_2887)
);

OAI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_2809),
.A2(n_230),
.B1(n_231),
.B2(n_229),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2841),
.Y(n_2889)
);

OAI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2776),
.A2(n_231),
.B1(n_232),
.B2(n_230),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2842),
.Y(n_2891)
);

OAI22xp33_ASAP7_75t_L g2892 ( 
.A1(n_2765),
.A2(n_2752),
.B1(n_2818),
.B2(n_2812),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2837),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2847),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2846),
.Y(n_2895)
);

OAI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2815),
.A2(n_228),
.B(n_233),
.Y(n_2896)
);

INVx1_ASAP7_75t_SL g2897 ( 
.A(n_2851),
.Y(n_2897)
);

NAND3xp33_ASAP7_75t_L g2898 ( 
.A(n_2855),
.B(n_234),
.C(n_235),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2798),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2848),
.Y(n_2900)
);

XNOR2x1_ASAP7_75t_L g2901 ( 
.A(n_2819),
.B(n_236),
.Y(n_2901)
);

AOI221xp5_ASAP7_75t_L g2902 ( 
.A1(n_2803),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2790),
.B(n_237),
.Y(n_2903)
);

INVx1_ASAP7_75t_SL g2904 ( 
.A(n_2789),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2792),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2850),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2854),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2759),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_2908)
);

XOR2x2_ASAP7_75t_L g2909 ( 
.A(n_2791),
.B(n_242),
.Y(n_2909)
);

OAI21xp33_ASAP7_75t_L g2910 ( 
.A1(n_2853),
.A2(n_242),
.B(n_243),
.Y(n_2910)
);

INVxp67_ASAP7_75t_SL g2911 ( 
.A(n_2795),
.Y(n_2911)
);

OAI21xp33_ASAP7_75t_L g2912 ( 
.A1(n_2788),
.A2(n_244),
.B(n_245),
.Y(n_2912)
);

XOR2xp5_ASAP7_75t_L g2913 ( 
.A(n_2819),
.B(n_244),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2857),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2785),
.A2(n_249),
.B1(n_246),
.B2(n_247),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2786),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2748),
.Y(n_2917)
);

AOI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2852),
.A2(n_250),
.B1(n_246),
.B2(n_249),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2824),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2919)
);

NAND4xp75_ASAP7_75t_L g2920 ( 
.A(n_2806),
.B(n_255),
.C(n_251),
.D(n_254),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2793),
.Y(n_2921)
);

NOR3xp33_ASAP7_75t_L g2922 ( 
.A(n_2754),
.B(n_254),
.C(n_256),
.Y(n_2922)
);

INVxp67_ASAP7_75t_L g2923 ( 
.A(n_2755),
.Y(n_2923)
);

OAI22xp33_ASAP7_75t_SL g2924 ( 
.A1(n_2823),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2924)
);

OAI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2782),
.A2(n_261),
.B1(n_258),
.B2(n_259),
.Y(n_2925)
);

XNOR2x1_ASAP7_75t_L g2926 ( 
.A(n_2822),
.B(n_2775),
.Y(n_2926)
);

OAI221xp5_ASAP7_75t_L g2927 ( 
.A1(n_2801),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2927)
);

OAI21xp33_ASAP7_75t_L g2928 ( 
.A1(n_2766),
.A2(n_262),
.B(n_263),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2835),
.B(n_264),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2810),
.Y(n_2930)
);

NAND3xp33_ASAP7_75t_SL g2931 ( 
.A(n_2779),
.B(n_266),
.C(n_267),
.Y(n_2931)
);

A2O1A1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2780),
.A2(n_274),
.B(n_283),
.C(n_266),
.Y(n_2932)
);

AO21x1_ASAP7_75t_SL g2933 ( 
.A1(n_2836),
.A2(n_267),
.B(n_268),
.Y(n_2933)
);

NOR3xp33_ASAP7_75t_L g2934 ( 
.A(n_2856),
.B(n_269),
.C(n_270),
.Y(n_2934)
);

OAI221xp5_ASAP7_75t_L g2935 ( 
.A1(n_2808),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_272),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2794),
.Y(n_2936)
);

OAI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2826),
.A2(n_271),
.B(n_272),
.Y(n_2937)
);

OAI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2784),
.A2(n_273),
.B(n_274),
.Y(n_2938)
);

OAI22xp33_ASAP7_75t_L g2939 ( 
.A1(n_2817),
.A2(n_276),
.B1(n_278),
.B2(n_275),
.Y(n_2939)
);

AOI211xp5_ASAP7_75t_L g2940 ( 
.A1(n_2832),
.A2(n_278),
.B(n_273),
.C(n_276),
.Y(n_2940)
);

OAI211xp5_ASAP7_75t_L g2941 ( 
.A1(n_2770),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2941)
);

OAI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2784),
.A2(n_2825),
.B(n_2761),
.Y(n_2942)
);

XNOR2x1_ASAP7_75t_L g2943 ( 
.A(n_2816),
.B(n_279),
.Y(n_2943)
);

AOI211xp5_ASAP7_75t_SL g2944 ( 
.A1(n_2827),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_2944)
);

XNOR2x2_ASAP7_75t_L g2945 ( 
.A(n_2821),
.B(n_282),
.Y(n_2945)
);

AOI211xp5_ASAP7_75t_L g2946 ( 
.A1(n_2813),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2811),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2947)
);

OAI221xp5_ASAP7_75t_SL g2948 ( 
.A1(n_2820),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.C(n_290),
.Y(n_2948)
);

AOI221xp5_ASAP7_75t_SL g2949 ( 
.A1(n_2787),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.C(n_290),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2799),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_2950)
);

OAI31xp33_ASAP7_75t_L g2951 ( 
.A1(n_2849),
.A2(n_293),
.A3(n_294),
.B(n_292),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2781),
.A2(n_2839),
.B1(n_2843),
.B2(n_2829),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2802),
.A2(n_296),
.B1(n_291),
.B2(n_295),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2844),
.A2(n_2777),
.B(n_2807),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2762),
.B(n_295),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2805),
.B(n_296),
.Y(n_2956)
);

AOI22xp33_ASAP7_75t_L g2957 ( 
.A1(n_2759),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_2957)
);

AOI21xp33_ASAP7_75t_L g2958 ( 
.A1(n_2768),
.A2(n_300),
.B(n_301),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2790),
.B(n_302),
.Y(n_2959)
);

INVxp67_ASAP7_75t_SL g2960 ( 
.A(n_2846),
.Y(n_2960)
);

OAI21xp33_ASAP7_75t_L g2961 ( 
.A1(n_2845),
.A2(n_302),
.B(n_303),
.Y(n_2961)
);

OAI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2796),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2962)
);

OAI221xp5_ASAP7_75t_L g2963 ( 
.A1(n_2774),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.C(n_307),
.Y(n_2963)
);

XNOR2xp5_ASAP7_75t_L g2964 ( 
.A(n_2773),
.B(n_306),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2751),
.B(n_307),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2763),
.Y(n_2966)
);

OAI21xp5_ASAP7_75t_SL g2967 ( 
.A1(n_2845),
.A2(n_308),
.B(n_309),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2814),
.A2(n_308),
.B(n_309),
.Y(n_2968)
);

AOI221xp5_ASAP7_75t_L g2969 ( 
.A1(n_2768),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.C(n_313),
.Y(n_2969)
);

OAI22xp33_ASAP7_75t_SL g2970 ( 
.A1(n_2758),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2763),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2763),
.Y(n_2972)
);

AOI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2774),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2763),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2756),
.B(n_314),
.Y(n_2975)
);

OAI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2814),
.A2(n_315),
.B(n_317),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2911),
.B(n_317),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2932),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_2978)
);

NOR2x1_ASAP7_75t_L g2979 ( 
.A(n_2903),
.B(n_2871),
.Y(n_2979)
);

OAI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_2967),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_2980)
);

AOI221xp5_ASAP7_75t_L g2981 ( 
.A1(n_2958),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.C(n_324),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2897),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2879),
.B(n_325),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2869),
.B(n_326),
.Y(n_2984)
);

INVxp67_ASAP7_75t_L g2985 ( 
.A(n_2933),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2881),
.B(n_328),
.Y(n_2986)
);

OR2x2_ASAP7_75t_L g2987 ( 
.A(n_2873),
.B(n_328),
.Y(n_2987)
);

OAI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2944),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2988)
);

AOI322xp5_ASAP7_75t_L g2989 ( 
.A1(n_2949),
.A2(n_335),
.A3(n_334),
.B1(n_332),
.B2(n_329),
.C1(n_330),
.C2(n_333),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2861),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2905),
.B(n_332),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2865),
.Y(n_2992)
);

NOR2x1_ASAP7_75t_L g2993 ( 
.A(n_2860),
.B(n_333),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2867),
.Y(n_2994)
);

INVx1_ASAP7_75t_SL g2995 ( 
.A(n_2926),
.Y(n_2995)
);

OAI211xp5_ASAP7_75t_L g2996 ( 
.A1(n_2940),
.A2(n_2882),
.B(n_2957),
.C(n_2908),
.Y(n_2996)
);

A2O1A1Ixp33_ASAP7_75t_L g2997 ( 
.A1(n_2858),
.A2(n_337),
.B(n_334),
.C(n_336),
.Y(n_2997)
);

INVxp67_ASAP7_75t_SL g2998 ( 
.A(n_2876),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2884),
.B(n_2885),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2889),
.B(n_336),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2872),
.Y(n_3001)
);

INVxp33_ASAP7_75t_L g3002 ( 
.A(n_2929),
.Y(n_3002)
);

A2O1A1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2910),
.A2(n_2961),
.B(n_2912),
.C(n_2968),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2866),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2891),
.B(n_337),
.Y(n_3005)
);

OAI21xp5_ASAP7_75t_SL g3006 ( 
.A1(n_2862),
.A2(n_339),
.B(n_340),
.Y(n_3006)
);

INVx1_ASAP7_75t_SL g3007 ( 
.A(n_2901),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2894),
.B(n_339),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2874),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2875),
.Y(n_3010)
);

AOI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2965),
.A2(n_341),
.B(n_343),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2900),
.B(n_2906),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2892),
.A2(n_345),
.B1(n_341),
.B2(n_343),
.Y(n_3013)
);

OAI32xp33_ASAP7_75t_L g3014 ( 
.A1(n_2922),
.A2(n_348),
.A3(n_346),
.B1(n_347),
.B2(n_350),
.Y(n_3014)
);

AOI32xp33_ASAP7_75t_L g3015 ( 
.A1(n_2934),
.A2(n_2943),
.A3(n_2946),
.B1(n_2888),
.B2(n_2890),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2916),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2970),
.A2(n_2928),
.B(n_2976),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2921),
.Y(n_3018)
);

AOI22xp5_ASAP7_75t_L g3019 ( 
.A1(n_2898),
.A2(n_350),
.B1(n_346),
.B2(n_348),
.Y(n_3019)
);

OAI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2877),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_3020)
);

OAI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_2923),
.A2(n_354),
.B1(n_351),
.B2(n_352),
.Y(n_3021)
);

OAI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2905),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2936),
.Y(n_3023)
);

NOR2xp67_ASAP7_75t_SL g3024 ( 
.A(n_2920),
.B(n_355),
.Y(n_3024)
);

HB1xp67_ASAP7_75t_L g3025 ( 
.A(n_2895),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2907),
.B(n_356),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2904),
.B(n_357),
.Y(n_3027)
);

O2A1O1Ixp5_ASAP7_75t_L g3028 ( 
.A1(n_2960),
.A2(n_360),
.B(n_358),
.C(n_359),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2966),
.Y(n_3029)
);

A2O1A1Ixp33_ASAP7_75t_L g3030 ( 
.A1(n_2878),
.A2(n_360),
.B(n_358),
.C(n_359),
.Y(n_3030)
);

OAI22xp33_ASAP7_75t_SL g3031 ( 
.A1(n_2935),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2917),
.B(n_362),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2913),
.Y(n_3033)
);

OAI221xp5_ASAP7_75t_L g3034 ( 
.A1(n_2964),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.C(n_366),
.Y(n_3034)
);

AOI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2880),
.A2(n_369),
.B1(n_366),
.B2(n_368),
.Y(n_3035)
);

OAI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2859),
.A2(n_2896),
.B(n_2886),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2914),
.B(n_368),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2971),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2972),
.B(n_370),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2931),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2974),
.B(n_371),
.Y(n_3041)
);

AOI221xp5_ASAP7_75t_L g3042 ( 
.A1(n_2924),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.C(n_375),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2959),
.B(n_373),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2975),
.B(n_374),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2955),
.B(n_2956),
.Y(n_3045)
);

INVx1_ASAP7_75t_SL g3046 ( 
.A(n_2909),
.Y(n_3046)
);

AOI211xp5_ASAP7_75t_L g3047 ( 
.A1(n_2927),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2956),
.Y(n_3048)
);

OAI22x1_ASAP7_75t_L g3049 ( 
.A1(n_2863),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3049)
);

INVxp67_ASAP7_75t_L g3050 ( 
.A(n_2945),
.Y(n_3050)
);

INVxp67_ASAP7_75t_L g3051 ( 
.A(n_2942),
.Y(n_3051)
);

NAND2x1p5_ASAP7_75t_L g3052 ( 
.A(n_2973),
.B(n_378),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2941),
.B(n_379),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2868),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2893),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_2952),
.Y(n_3056)
);

O2A1O1Ixp33_ASAP7_75t_SL g3057 ( 
.A1(n_2938),
.A2(n_2962),
.B(n_2864),
.C(n_2937),
.Y(n_3057)
);

AOI221x1_ASAP7_75t_L g3058 ( 
.A1(n_2899),
.A2(n_2925),
.B1(n_2954),
.B2(n_2930),
.C(n_2948),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2947),
.B(n_379),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2953),
.Y(n_3060)
);

OAI21xp33_ASAP7_75t_SL g3061 ( 
.A1(n_2887),
.A2(n_380),
.B(n_381),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2870),
.A2(n_2969),
.B(n_2902),
.Y(n_3062)
);

NOR3xp33_ASAP7_75t_L g3063 ( 
.A(n_2963),
.B(n_380),
.C(n_381),
.Y(n_3063)
);

AOI21xp33_ASAP7_75t_L g3064 ( 
.A1(n_2939),
.A2(n_382),
.B(n_383),
.Y(n_3064)
);

OA21x2_ASAP7_75t_L g3065 ( 
.A1(n_2883),
.A2(n_383),
.B(n_384),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2919),
.Y(n_3066)
);

OAI221xp5_ASAP7_75t_SL g3067 ( 
.A1(n_2951),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.C(n_387),
.Y(n_3067)
);

XNOR2x2_ASAP7_75t_L g3068 ( 
.A(n_2918),
.B(n_385),
.Y(n_3068)
);

OAI321xp33_ASAP7_75t_L g3069 ( 
.A1(n_2915),
.A2(n_2950),
.A3(n_389),
.B1(n_391),
.B2(n_387),
.C(n_388),
.Y(n_3069)
);

NOR3xp33_ASAP7_75t_SL g3070 ( 
.A(n_2882),
.B(n_388),
.C(n_390),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2911),
.B(n_391),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2911),
.B(n_392),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2866),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2866),
.Y(n_3074)
);

AOI321xp33_ASAP7_75t_L g3075 ( 
.A1(n_2940),
.A2(n_395),
.A3(n_397),
.B1(n_393),
.B2(n_394),
.C(n_396),
.Y(n_3075)
);

OAI22xp33_ASAP7_75t_SL g3076 ( 
.A1(n_2871),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2873),
.Y(n_3077)
);

OAI322xp33_ASAP7_75t_L g3078 ( 
.A1(n_2945),
.A2(n_401),
.A3(n_400),
.B1(n_398),
.B2(n_396),
.C1(n_397),
.C2(n_399),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2873),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2866),
.Y(n_3080)
);

INVx1_ASAP7_75t_SL g3081 ( 
.A(n_2897),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2873),
.Y(n_3082)
);

INVxp67_ASAP7_75t_L g3083 ( 
.A(n_2933),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2873),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2932),
.A2(n_402),
.B1(n_398),
.B2(n_400),
.Y(n_3085)
);

AOI21xp33_ASAP7_75t_L g3086 ( 
.A1(n_2858),
.A2(n_402),
.B(n_403),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_SL g3087 ( 
.A(n_2879),
.B(n_404),
.Y(n_3087)
);

AOI222xp33_ASAP7_75t_L g3088 ( 
.A1(n_2967),
.A2(n_406),
.B1(n_408),
.B2(n_404),
.C1(n_405),
.C2(n_407),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2873),
.Y(n_3089)
);

BUFx2_ASAP7_75t_L g3090 ( 
.A(n_2911),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2879),
.B(n_405),
.Y(n_3091)
);

A2O1A1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2932),
.A2(n_410),
.B(n_406),
.C(n_409),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2911),
.B(n_409),
.Y(n_3093)
);

INVxp67_ASAP7_75t_L g3094 ( 
.A(n_2933),
.Y(n_3094)
);

AOI221xp5_ASAP7_75t_L g3095 ( 
.A1(n_2932),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.C(n_413),
.Y(n_3095)
);

OAI21xp33_ASAP7_75t_L g3096 ( 
.A1(n_2967),
.A2(n_412),
.B(n_413),
.Y(n_3096)
);

NAND3xp33_ASAP7_75t_L g3097 ( 
.A(n_2932),
.B(n_415),
.C(n_416),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2879),
.B(n_415),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2911),
.B(n_416),
.Y(n_3099)
);

INVx2_ASAP7_75t_SL g3100 ( 
.A(n_2897),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2897),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2905),
.B(n_417),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2911),
.B(n_417),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2873),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2932),
.A2(n_418),
.B(n_419),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2873),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2866),
.Y(n_3107)
);

AOI221x1_ASAP7_75t_SL g3108 ( 
.A1(n_2940),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.C(n_421),
.Y(n_3108)
);

OAI211xp5_ASAP7_75t_L g3109 ( 
.A1(n_2967),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_3109)
);

INVx1_ASAP7_75t_SL g3110 ( 
.A(n_2897),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2873),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2866),
.Y(n_3112)
);

A2O1A1Ixp33_ASAP7_75t_L g3113 ( 
.A1(n_2932),
.A2(n_426),
.B(n_422),
.C(n_425),
.Y(n_3113)
);

OAI221xp5_ASAP7_75t_L g3114 ( 
.A1(n_2932),
.A2(n_428),
.B1(n_425),
.B2(n_427),
.C(n_429),
.Y(n_3114)
);

AOI21xp33_ASAP7_75t_SL g3115 ( 
.A1(n_2860),
.A2(n_427),
.B(n_428),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2873),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2967),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_3117)
);

OAI22xp33_ASAP7_75t_SL g3118 ( 
.A1(n_2871),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_3118)
);

AOI221x1_ASAP7_75t_L g3119 ( 
.A1(n_2932),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.C(n_435),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2873),
.Y(n_3120)
);

OAI21xp33_ASAP7_75t_L g3121 ( 
.A1(n_2967),
.A2(n_433),
.B(n_434),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2879),
.B(n_435),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2873),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2873),
.Y(n_3124)
);

A2O1A1Ixp33_ASAP7_75t_L g3125 ( 
.A1(n_2932),
.A2(n_438),
.B(n_436),
.C(n_437),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_SL g3126 ( 
.A(n_2897),
.B(n_436),
.Y(n_3126)
);

AO21x1_ASAP7_75t_L g3127 ( 
.A1(n_2943),
.A2(n_437),
.B(n_438),
.Y(n_3127)
);

AOI21xp33_ASAP7_75t_L g3128 ( 
.A1(n_2858),
.A2(n_439),
.B(n_440),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2866),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2911),
.B(n_439),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_2911),
.B(n_440),
.Y(n_3131)
);

AOI222xp33_ASAP7_75t_L g3132 ( 
.A1(n_2967),
.A2(n_443),
.B1(n_446),
.B2(n_441),
.C1(n_442),
.C2(n_444),
.Y(n_3132)
);

AOI311xp33_ASAP7_75t_L g3133 ( 
.A1(n_2922),
.A2(n_443),
.A3(n_441),
.B(n_442),
.C(n_444),
.Y(n_3133)
);

OAI211xp5_ASAP7_75t_L g3134 ( 
.A1(n_2967),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_3134)
);

OAI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_2932),
.A2(n_450),
.B1(n_447),
.B2(n_448),
.Y(n_3135)
);

O2A1O1Ixp33_ASAP7_75t_L g3136 ( 
.A1(n_2932),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_3136)
);

INVxp67_ASAP7_75t_SL g3137 ( 
.A(n_2876),
.Y(n_3137)
);

OAI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2932),
.A2(n_452),
.B(n_454),
.Y(n_3138)
);

OAI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2967),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2911),
.B(n_456),
.Y(n_3140)
);

AOI221xp5_ASAP7_75t_L g3141 ( 
.A1(n_2932),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.C(n_461),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2911),
.B(n_460),
.Y(n_3142)
);

OAI33xp33_ASAP7_75t_L g3143 ( 
.A1(n_2970),
.A2(n_464),
.A3(n_466),
.B1(n_462),
.B2(n_463),
.B3(n_465),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2911),
.B(n_462),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2873),
.Y(n_3145)
);

OAI32xp33_ASAP7_75t_L g3146 ( 
.A1(n_2882),
.A2(n_465),
.A3(n_463),
.B1(n_464),
.B2(n_466),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2873),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2911),
.B(n_467),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2905),
.B(n_468),
.Y(n_3149)
);

AOI221xp5_ASAP7_75t_L g3150 ( 
.A1(n_2998),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.C(n_472),
.Y(n_3150)
);

AOI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_3137),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_3050),
.A2(n_472),
.B(n_474),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2999),
.Y(n_3153)
);

AOI221xp5_ASAP7_75t_L g3154 ( 
.A1(n_3108),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.C(n_478),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_3081),
.B(n_476),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3012),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2990),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_SL g3158 ( 
.A(n_2995),
.B(n_478),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_L g3159 ( 
.A(n_2985),
.B(n_479),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_3083),
.B(n_479),
.Y(n_3160)
);

AOI21xp33_ASAP7_75t_SL g3161 ( 
.A1(n_3094),
.A2(n_480),
.B(n_481),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2992),
.Y(n_3162)
);

NAND2xp33_ASAP7_75t_SL g3163 ( 
.A(n_3100),
.B(n_481),
.Y(n_3163)
);

NAND3xp33_ASAP7_75t_L g3164 ( 
.A(n_3058),
.B(n_482),
.C(n_483),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_3101),
.B(n_484),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_3110),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_3090),
.Y(n_3167)
);

NOR2x1_ASAP7_75t_SL g3168 ( 
.A(n_3131),
.B(n_484),
.Y(n_3168)
);

NOR2x1_ASAP7_75t_L g3169 ( 
.A(n_2993),
.B(n_485),
.Y(n_3169)
);

NOR3xp33_ASAP7_75t_L g3170 ( 
.A(n_3109),
.B(n_485),
.C(n_486),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_3056),
.B(n_486),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_3002),
.B(n_487),
.Y(n_3172)
);

NAND3xp33_ASAP7_75t_SL g3173 ( 
.A(n_3127),
.B(n_488),
.C(n_489),
.Y(n_3173)
);

NOR3x1_ASAP7_75t_L g3174 ( 
.A(n_3006),
.B(n_488),
.C(n_489),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_2987),
.B(n_490),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_3046),
.B(n_490),
.Y(n_3176)
);

NOR3xp33_ASAP7_75t_L g3177 ( 
.A(n_3134),
.B(n_491),
.C(n_492),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_2979),
.B(n_493),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_3144),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3025),
.B(n_493),
.Y(n_3180)
);

HB1xp67_ASAP7_75t_L g3181 ( 
.A(n_3051),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_3087),
.B(n_494),
.Y(n_3182)
);

OAI21xp33_ASAP7_75t_L g3183 ( 
.A1(n_3096),
.A2(n_495),
.B(n_497),
.Y(n_3183)
);

AOI211xp5_ASAP7_75t_SL g3184 ( 
.A1(n_2980),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_3184)
);

OAI211xp5_ASAP7_75t_L g3185 ( 
.A1(n_3133),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3185)
);

INVx8_ASAP7_75t_L g3186 ( 
.A(n_2991),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3077),
.B(n_500),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_3079),
.B(n_501),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3082),
.B(n_502),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2994),
.Y(n_3190)
);

OAI211xp5_ASAP7_75t_L g3191 ( 
.A1(n_3121),
.A2(n_504),
.B(n_502),
.C(n_503),
.Y(n_3191)
);

NOR2x1_ASAP7_75t_SL g3192 ( 
.A(n_3039),
.B(n_503),
.Y(n_3192)
);

AOI221xp5_ASAP7_75t_L g3193 ( 
.A1(n_3143),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.C(n_508),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_3033),
.Y(n_3194)
);

AOI221xp5_ASAP7_75t_L g3195 ( 
.A1(n_3003),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.C(n_509),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_3084),
.B(n_509),
.Y(n_3196)
);

HB1xp67_ASAP7_75t_L g3197 ( 
.A(n_3001),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_2986),
.B(n_510),
.Y(n_3198)
);

AOI221xp5_ASAP7_75t_L g3199 ( 
.A1(n_3062),
.A2(n_513),
.B1(n_510),
.B2(n_511),
.C(n_514),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3009),
.Y(n_3200)
);

NAND2x1_ASAP7_75t_L g3201 ( 
.A(n_3010),
.B(n_515),
.Y(n_3201)
);

XOR2x2_ASAP7_75t_L g3202 ( 
.A(n_3068),
.B(n_515),
.Y(n_3202)
);

NOR3xp33_ASAP7_75t_SL g3203 ( 
.A(n_2996),
.B(n_516),
.C(n_517),
.Y(n_3203)
);

O2A1O1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_3139),
.A2(n_521),
.B(n_519),
.C(n_520),
.Y(n_3204)
);

AOI221xp5_ASAP7_75t_L g3205 ( 
.A1(n_3078),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.C(n_523),
.Y(n_3205)
);

NOR2xp67_ASAP7_75t_L g3206 ( 
.A(n_3013),
.B(n_523),
.Y(n_3206)
);

OAI221xp5_ASAP7_75t_L g3207 ( 
.A1(n_3036),
.A2(n_527),
.B1(n_524),
.B2(n_526),
.C(n_528),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_3089),
.B(n_524),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3016),
.Y(n_3209)
);

AOI221xp5_ASAP7_75t_L g3210 ( 
.A1(n_3031),
.A2(n_3017),
.B1(n_3057),
.B2(n_3138),
.C(n_3136),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3104),
.B(n_527),
.Y(n_3211)
);

AOI21xp33_ASAP7_75t_L g3212 ( 
.A1(n_3088),
.A2(n_3132),
.B(n_3118),
.Y(n_3212)
);

XNOR2xp5_ASAP7_75t_L g3213 ( 
.A(n_3007),
.B(n_528),
.Y(n_3213)
);

NOR3x1_ASAP7_75t_L g3214 ( 
.A(n_3097),
.B(n_529),
.C(n_530),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3106),
.B(n_529),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3018),
.Y(n_3216)
);

AOI221x1_ASAP7_75t_L g3217 ( 
.A1(n_3105),
.A2(n_3063),
.B1(n_3135),
.B2(n_3085),
.C(n_2978),
.Y(n_3217)
);

OAI221xp5_ASAP7_75t_L g3218 ( 
.A1(n_3015),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.C(n_534),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_SL g3219 ( 
.A(n_3111),
.B(n_531),
.Y(n_3219)
);

OR2x2_ASAP7_75t_L g3220 ( 
.A(n_3116),
.B(n_532),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3032),
.B(n_533),
.Y(n_3221)
);

NAND4xp25_ASAP7_75t_L g3222 ( 
.A(n_3117),
.B(n_536),
.C(n_534),
.D(n_535),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3120),
.B(n_535),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3023),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_3123),
.B(n_3124),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3029),
.Y(n_3226)
);

NOR3xp33_ASAP7_75t_SL g3227 ( 
.A(n_2988),
.B(n_536),
.C(n_537),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_3038),
.Y(n_3228)
);

NOR2xp33_ASAP7_75t_L g3229 ( 
.A(n_3000),
.B(n_538),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_3102),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_3005),
.B(n_539),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_3008),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_3026),
.B(n_539),
.Y(n_3233)
);

AOI211xp5_ASAP7_75t_L g3234 ( 
.A1(n_3014),
.A2(n_542),
.B(n_540),
.C(n_541),
.Y(n_3234)
);

NOR3x1_ASAP7_75t_L g3235 ( 
.A(n_3027),
.B(n_541),
.C(n_542),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3145),
.Y(n_3236)
);

NOR2xp67_ASAP7_75t_L g3237 ( 
.A(n_2977),
.B(n_543),
.Y(n_3237)
);

AOI211xp5_ASAP7_75t_L g3238 ( 
.A1(n_3076),
.A2(n_547),
.B(n_544),
.C(n_546),
.Y(n_3238)
);

AOI221xp5_ASAP7_75t_L g3239 ( 
.A1(n_3086),
.A2(n_548),
.B1(n_544),
.B2(n_547),
.C(n_549),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3048),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3147),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3054),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_3037),
.B(n_548),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3055),
.Y(n_3244)
);

NAND2xp33_ASAP7_75t_L g3245 ( 
.A(n_3070),
.B(n_550),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3060),
.B(n_551),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3071),
.B(n_3072),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2984),
.Y(n_3248)
);

OAI21xp33_ASAP7_75t_L g3249 ( 
.A1(n_2989),
.A2(n_551),
.B(n_552),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3041),
.Y(n_3250)
);

NAND3xp33_ASAP7_75t_L g3251 ( 
.A(n_3075),
.B(n_553),
.C(n_554),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3126),
.A2(n_553),
.B(n_554),
.Y(n_3252)
);

O2A1O1Ixp33_ASAP7_75t_L g3253 ( 
.A1(n_2997),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_L g3254 ( 
.A(n_3044),
.B(n_556),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3092),
.A2(n_3125),
.B(n_3113),
.Y(n_3255)
);

AOI221xp5_ASAP7_75t_L g3256 ( 
.A1(n_3128),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.C(n_561),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_3043),
.B(n_558),
.Y(n_3257)
);

OR2x2_ASAP7_75t_L g3258 ( 
.A(n_3093),
.B(n_3099),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3103),
.B(n_559),
.Y(n_3259)
);

NOR3xp33_ASAP7_75t_SL g3260 ( 
.A(n_2983),
.B(n_560),
.C(n_562),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3028),
.A2(n_562),
.B(n_563),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3130),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3140),
.B(n_563),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3142),
.B(n_564),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_3149),
.B(n_564),
.Y(n_3265)
);

INVxp33_ASAP7_75t_SL g3266 ( 
.A(n_3091),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3148),
.B(n_3066),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3065),
.B(n_3059),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_SL g3269 ( 
.A(n_3067),
.B(n_565),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3065),
.B(n_566),
.Y(n_3270)
);

NOR4xp25_ASAP7_75t_L g3271 ( 
.A(n_3034),
.B(n_569),
.C(n_566),
.D(n_568),
.Y(n_3271)
);

OAI221xp5_ASAP7_75t_L g3272 ( 
.A1(n_3061),
.A2(n_571),
.B1(n_568),
.B2(n_570),
.C(n_572),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3053),
.B(n_570),
.Y(n_3273)
);

AOI221xp5_ASAP7_75t_L g3274 ( 
.A1(n_3114),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.C(n_574),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3045),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3115),
.B(n_573),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3021),
.B(n_574),
.Y(n_3277)
);

NAND4xp25_ASAP7_75t_L g3278 ( 
.A(n_3164),
.B(n_3098),
.C(n_3122),
.D(n_3047),
.Y(n_3278)
);

OAI21xp33_ASAP7_75t_SL g3279 ( 
.A1(n_3181),
.A2(n_3040),
.B(n_3019),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3194),
.B(n_3042),
.Y(n_3280)
);

NOR2x1_ASAP7_75t_L g3281 ( 
.A(n_3173),
.B(n_2982),
.Y(n_3281)
);

OAI211xp5_ASAP7_75t_SL g3282 ( 
.A1(n_3210),
.A2(n_3141),
.B(n_3095),
.C(n_3011),
.Y(n_3282)
);

NOR3xp33_ASAP7_75t_L g3283 ( 
.A(n_3185),
.B(n_3069),
.C(n_3020),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3179),
.B(n_3119),
.Y(n_3284)
);

NOR3x1_ASAP7_75t_L g3285 ( 
.A(n_3230),
.B(n_3022),
.C(n_3024),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3249),
.A2(n_3052),
.B1(n_3049),
.B2(n_3035),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3192),
.Y(n_3287)
);

AOI211xp5_ASAP7_75t_L g3288 ( 
.A1(n_3212),
.A2(n_3146),
.B(n_3064),
.C(n_3030),
.Y(n_3288)
);

NOR3xp33_ASAP7_75t_L g3289 ( 
.A(n_3251),
.B(n_2981),
.C(n_3004),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3197),
.Y(n_3290)
);

NOR2x1p5_ASAP7_75t_L g3291 ( 
.A(n_3166),
.B(n_3073),
.Y(n_3291)
);

CKINVDCx6p67_ASAP7_75t_R g3292 ( 
.A(n_3259),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3228),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3179),
.B(n_3167),
.Y(n_3294)
);

OA22x2_ASAP7_75t_L g3295 ( 
.A1(n_3217),
.A2(n_3080),
.B1(n_3107),
.B2(n_3074),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3178),
.A2(n_3129),
.B(n_3112),
.Y(n_3296)
);

OAI222xp33_ASAP7_75t_L g3297 ( 
.A1(n_3268),
.A2(n_577),
.B1(n_579),
.B2(n_575),
.C1(n_576),
.C2(n_578),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3266),
.B(n_575),
.Y(n_3298)
);

OAI21xp33_ASAP7_75t_SL g3299 ( 
.A1(n_3225),
.A2(n_576),
.B(n_577),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3157),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3152),
.A2(n_578),
.B(n_579),
.Y(n_3301)
);

AO22x2_ASAP7_75t_L g3302 ( 
.A1(n_3262),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_3186),
.Y(n_3303)
);

AOI31xp33_ASAP7_75t_L g3304 ( 
.A1(n_3154),
.A2(n_582),
.A3(n_580),
.B(n_581),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3162),
.Y(n_3305)
);

NOR2x1_ASAP7_75t_L g3306 ( 
.A(n_3155),
.B(n_583),
.Y(n_3306)
);

OAI21xp5_ASAP7_75t_SL g3307 ( 
.A1(n_3184),
.A2(n_583),
.B(n_584),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3255),
.A2(n_584),
.B(n_585),
.Y(n_3308)
);

NOR3x1_ASAP7_75t_L g3309 ( 
.A(n_3218),
.B(n_3275),
.C(n_3261),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_3203),
.A2(n_586),
.B(n_587),
.Y(n_3310)
);

OAI22xp33_ASAP7_75t_SL g3311 ( 
.A1(n_3158),
.A2(n_590),
.B1(n_586),
.B2(n_588),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3163),
.A2(n_588),
.B(n_590),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3232),
.B(n_591),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3271),
.B(n_591),
.Y(n_3314)
);

OAI222xp33_ASAP7_75t_L g3315 ( 
.A1(n_3151),
.A2(n_595),
.B1(n_598),
.B2(n_592),
.C1(n_594),
.C2(n_597),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3172),
.B(n_592),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3190),
.Y(n_3317)
);

OAI21xp33_ASAP7_75t_SL g3318 ( 
.A1(n_3153),
.A2(n_594),
.B(n_597),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3250),
.B(n_598),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_3202),
.A2(n_599),
.B(n_600),
.Y(n_3320)
);

AOI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3193),
.A2(n_603),
.B1(n_599),
.B2(n_600),
.Y(n_3321)
);

NOR2x1_ASAP7_75t_L g3322 ( 
.A(n_3169),
.B(n_603),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3248),
.B(n_604),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3245),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3171),
.A2(n_605),
.B(n_606),
.Y(n_3325)
);

NOR2x1_ASAP7_75t_L g3326 ( 
.A(n_3201),
.B(n_607),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3220),
.B(n_607),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3200),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3209),
.Y(n_3329)
);

INVxp67_ASAP7_75t_L g3330 ( 
.A(n_3168),
.Y(n_3330)
);

BUFx2_ASAP7_75t_L g3331 ( 
.A(n_3186),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_3165),
.A2(n_608),
.B(n_609),
.Y(n_3332)
);

AOI22x1_ASAP7_75t_L g3333 ( 
.A1(n_3156),
.A2(n_612),
.B1(n_608),
.B2(n_611),
.Y(n_3333)
);

OAI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3258),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3334)
);

NOR3xp33_ASAP7_75t_L g3335 ( 
.A(n_3191),
.B(n_614),
.C(n_615),
.Y(n_3335)
);

AND4x1_ASAP7_75t_L g3336 ( 
.A(n_3174),
.B(n_616),
.C(n_614),
.D(n_615),
.Y(n_3336)
);

AOI21xp33_ASAP7_75t_SL g3337 ( 
.A1(n_3186),
.A2(n_616),
.B(n_617),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_3273),
.A2(n_617),
.B(n_618),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3216),
.Y(n_3339)
);

AOI21xp33_ASAP7_75t_L g3340 ( 
.A1(n_3236),
.A2(n_618),
.B(n_619),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3247),
.B(n_619),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3302),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_SL g3343 ( 
.A(n_3330),
.B(n_3176),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3331),
.B(n_3159),
.Y(n_3344)
);

AOI221xp5_ASAP7_75t_L g3345 ( 
.A1(n_3304),
.A2(n_3205),
.B1(n_3195),
.B2(n_3177),
.C(n_3170),
.Y(n_3345)
);

AOI221xp5_ASAP7_75t_L g3346 ( 
.A1(n_3283),
.A2(n_3284),
.B1(n_3279),
.B2(n_3282),
.C(n_3318),
.Y(n_3346)
);

OAI322xp33_ASAP7_75t_L g3347 ( 
.A1(n_3295),
.A2(n_3269),
.A3(n_3277),
.B1(n_3276),
.B2(n_3219),
.C1(n_3196),
.C2(n_3188),
.Y(n_3347)
);

OAI22x1_ASAP7_75t_L g3348 ( 
.A1(n_3336),
.A2(n_3240),
.B1(n_3213),
.B2(n_3265),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_R g3349 ( 
.A(n_3303),
.B(n_3160),
.Y(n_3349)
);

AOI211xp5_ASAP7_75t_SL g3350 ( 
.A1(n_3303),
.A2(n_3183),
.B(n_3234),
.C(n_3150),
.Y(n_3350)
);

NOR4xp25_ASAP7_75t_L g3351 ( 
.A(n_3314),
.B(n_3222),
.C(n_3204),
.D(n_3253),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3281),
.A2(n_3206),
.B1(n_3237),
.B2(n_3238),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3320),
.A2(n_3270),
.B(n_3267),
.Y(n_3353)
);

OAI211xp5_ASAP7_75t_L g3354 ( 
.A1(n_3307),
.A2(n_3161),
.B(n_3227),
.C(n_3199),
.Y(n_3354)
);

OAI211xp5_ASAP7_75t_L g3355 ( 
.A1(n_3299),
.A2(n_3252),
.B(n_3207),
.C(n_3274),
.Y(n_3355)
);

AOI221xp5_ASAP7_75t_L g3356 ( 
.A1(n_3308),
.A2(n_3272),
.B1(n_3189),
.B2(n_3215),
.C(n_3211),
.Y(n_3356)
);

AOI21xp33_ASAP7_75t_L g3357 ( 
.A1(n_3288),
.A2(n_3241),
.B(n_3242),
.Y(n_3357)
);

AOI221xp5_ASAP7_75t_SL g3358 ( 
.A1(n_3337),
.A2(n_3208),
.B1(n_3180),
.B2(n_3182),
.C(n_3224),
.Y(n_3358)
);

NOR2x1_ASAP7_75t_L g3359 ( 
.A(n_3326),
.B(n_3187),
.Y(n_3359)
);

OAI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3312),
.A2(n_3260),
.B(n_3175),
.Y(n_3360)
);

O2A1O1Ixp5_ASAP7_75t_L g3361 ( 
.A1(n_3294),
.A2(n_3226),
.B(n_3229),
.C(n_3198),
.Y(n_3361)
);

AOI221xp5_ASAP7_75t_L g3362 ( 
.A1(n_3289),
.A2(n_3223),
.B1(n_3243),
.B2(n_3233),
.C(n_3231),
.Y(n_3362)
);

OAI21xp33_ASAP7_75t_SL g3363 ( 
.A1(n_3290),
.A2(n_3264),
.B(n_3263),
.Y(n_3363)
);

AOI221xp5_ASAP7_75t_SL g3364 ( 
.A1(n_3278),
.A2(n_3239),
.B1(n_3256),
.B2(n_3257),
.C(n_3246),
.Y(n_3364)
);

AOI221xp5_ASAP7_75t_L g3365 ( 
.A1(n_3297),
.A2(n_3254),
.B1(n_3244),
.B2(n_3221),
.C(n_3214),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3287),
.Y(n_3366)
);

NAND3xp33_ASAP7_75t_L g3367 ( 
.A(n_3335),
.B(n_3310),
.C(n_3321),
.Y(n_3367)
);

AOI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_3322),
.A2(n_3235),
.B(n_620),
.Y(n_3368)
);

AOI221xp5_ASAP7_75t_L g3369 ( 
.A1(n_3301),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.C(n_623),
.Y(n_3369)
);

OAI211xp5_ASAP7_75t_SL g3370 ( 
.A1(n_3293),
.A2(n_626),
.B(n_622),
.C(n_624),
.Y(n_3370)
);

AOI221xp5_ASAP7_75t_L g3371 ( 
.A1(n_3280),
.A2(n_627),
.B1(n_624),
.B2(n_626),
.C(n_628),
.Y(n_3371)
);

NAND4xp75_ASAP7_75t_L g3372 ( 
.A(n_3285),
.B(n_629),
.C(n_627),
.D(n_628),
.Y(n_3372)
);

AOI21xp33_ASAP7_75t_SL g3373 ( 
.A1(n_3298),
.A2(n_629),
.B(n_631),
.Y(n_3373)
);

OAI21xp33_ASAP7_75t_L g3374 ( 
.A1(n_3286),
.A2(n_631),
.B(n_632),
.Y(n_3374)
);

AOI221xp5_ASAP7_75t_L g3375 ( 
.A1(n_3338),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.C(n_635),
.Y(n_3375)
);

AOI221xp5_ASAP7_75t_SL g3376 ( 
.A1(n_3332),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.C(n_636),
.Y(n_3376)
);

NOR4xp25_ASAP7_75t_L g3377 ( 
.A(n_3300),
.B(n_639),
.C(n_637),
.D(n_638),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3344),
.B(n_3292),
.Y(n_3378)
);

NOR2x1_ASAP7_75t_L g3379 ( 
.A(n_3372),
.B(n_3323),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3342),
.Y(n_3380)
);

AO22x2_ASAP7_75t_L g3381 ( 
.A1(n_3353),
.A2(n_3317),
.B1(n_3328),
.B2(n_3305),
.Y(n_3381)
);

NOR4xp25_ASAP7_75t_L g3382 ( 
.A(n_3346),
.B(n_3315),
.C(n_3339),
.D(n_3329),
.Y(n_3382)
);

AOI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3343),
.A2(n_3306),
.B1(n_3291),
.B2(n_3324),
.Y(n_3383)
);

AND2x2_ASAP7_75t_SL g3384 ( 
.A(n_3351),
.B(n_3309),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3366),
.Y(n_3385)
);

NOR2x1_ASAP7_75t_L g3386 ( 
.A(n_3354),
.B(n_3319),
.Y(n_3386)
);

NOR2x1_ASAP7_75t_L g3387 ( 
.A(n_3347),
.B(n_3313),
.Y(n_3387)
);

INVxp33_ASAP7_75t_L g3388 ( 
.A(n_3349),
.Y(n_3388)
);

AOI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3352),
.A2(n_3302),
.B1(n_3341),
.B2(n_3311),
.Y(n_3389)
);

NAND3xp33_ASAP7_75t_L g3390 ( 
.A(n_3367),
.B(n_3333),
.C(n_3340),
.Y(n_3390)
);

NOR2x1_ASAP7_75t_L g3391 ( 
.A(n_3370),
.B(n_3316),
.Y(n_3391)
);

AOI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3348),
.A2(n_3345),
.B1(n_3355),
.B2(n_3356),
.Y(n_3392)
);

AOI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_3365),
.A2(n_3296),
.B1(n_3334),
.B2(n_3325),
.Y(n_3393)
);

NOR2x1_ASAP7_75t_L g3394 ( 
.A(n_3359),
.B(n_3327),
.Y(n_3394)
);

AOI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_3364),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_3395)
);

NOR2x1_ASAP7_75t_L g3396 ( 
.A(n_3368),
.B(n_640),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3374),
.Y(n_3397)
);

NOR2x1_ASAP7_75t_L g3398 ( 
.A(n_3378),
.B(n_3360),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3384),
.Y(n_3399)
);

AOI211xp5_ASAP7_75t_SL g3400 ( 
.A1(n_3392),
.A2(n_3357),
.B(n_3375),
.C(n_3369),
.Y(n_3400)
);

AND3x2_ASAP7_75t_L g3401 ( 
.A(n_3382),
.B(n_3377),
.C(n_3371),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3380),
.Y(n_3402)
);

AND3x2_ASAP7_75t_L g3403 ( 
.A(n_3385),
.B(n_3362),
.C(n_3376),
.Y(n_3403)
);

AOI211xp5_ASAP7_75t_L g3404 ( 
.A1(n_3390),
.A2(n_3363),
.B(n_3358),
.C(n_3373),
.Y(n_3404)
);

NOR3xp33_ASAP7_75t_SL g3405 ( 
.A(n_3397),
.B(n_3388),
.C(n_3381),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3394),
.B(n_3350),
.Y(n_3406)
);

NAND2xp33_ASAP7_75t_SL g3407 ( 
.A(n_3381),
.B(n_3361),
.Y(n_3407)
);

NOR3xp33_ASAP7_75t_SL g3408 ( 
.A(n_3386),
.B(n_641),
.C(n_643),
.Y(n_3408)
);

BUFx2_ASAP7_75t_L g3409 ( 
.A(n_3407),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3398),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3399),
.B(n_3391),
.Y(n_3411)
);

AOI22x1_ASAP7_75t_L g3412 ( 
.A1(n_3402),
.A2(n_3400),
.B1(n_3405),
.B2(n_3401),
.Y(n_3412)
);

CKINVDCx5p33_ASAP7_75t_R g3413 ( 
.A(n_3408),
.Y(n_3413)
);

BUFx6f_ASAP7_75t_L g3414 ( 
.A(n_3406),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3403),
.Y(n_3415)
);

BUFx6f_ASAP7_75t_L g3416 ( 
.A(n_3404),
.Y(n_3416)
);

CKINVDCx14_ASAP7_75t_R g3417 ( 
.A(n_3399),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3398),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3410),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3418),
.Y(n_3420)
);

AND2x4_ASAP7_75t_L g3421 ( 
.A(n_3414),
.B(n_3396),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3412),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3417),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3415),
.Y(n_3424)
);

AO22x2_ASAP7_75t_L g3425 ( 
.A1(n_3423),
.A2(n_3411),
.B1(n_3409),
.B2(n_3413),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3420),
.Y(n_3426)
);

OAI22x1_ASAP7_75t_L g3427 ( 
.A1(n_3421),
.A2(n_3395),
.B1(n_3387),
.B2(n_3389),
.Y(n_3427)
);

OAI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3426),
.A2(n_3414),
.B1(n_3424),
.B2(n_3422),
.Y(n_3428)
);

OAI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_3425),
.A2(n_3419),
.B(n_3393),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_SL g3430 ( 
.A1(n_3427),
.A2(n_3416),
.B1(n_3383),
.B2(n_3379),
.Y(n_3430)
);

XNOR2x1_ASAP7_75t_L g3431 ( 
.A(n_3427),
.B(n_3416),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3431),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3430),
.A2(n_644),
.B1(n_641),
.B2(n_643),
.Y(n_3433)
);

OAI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3433),
.A2(n_3429),
.B(n_3428),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3434),
.A2(n_3432),
.B1(n_646),
.B2(n_644),
.Y(n_3435)
);

OR2x6_ASAP7_75t_L g3436 ( 
.A(n_3435),
.B(n_645),
.Y(n_3436)
);

AOI31xp33_ASAP7_75t_L g3437 ( 
.A1(n_3436),
.A2(n_648),
.A3(n_645),
.B(n_647),
.Y(n_3437)
);


endmodule