module real_aes_8471_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_1), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_1), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_2), .A2(n_148), .B(n_153), .C(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_3), .A2(n_143), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g505 ( .A(n_4), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_5), .B(n_181), .Y(n_247) );
AOI21xp33_ASAP7_75t_L g512 ( .A1(n_6), .A2(n_143), .B(n_513), .Y(n_512) );
AND2x6_ASAP7_75t_L g148 ( .A(n_7), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_8), .A2(n_278), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g160 ( .A(n_9), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_10), .B(n_43), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_11), .A2(n_33), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_11), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_12), .B(n_158), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_13), .B(n_205), .Y(n_484) );
INVx1_ASAP7_75t_L g517 ( .A(n_14), .Y(n_517) );
INVx1_ASAP7_75t_L g141 ( .A(n_15), .Y(n_141) );
INVx1_ASAP7_75t_L g496 ( .A(n_16), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_17), .A2(n_161), .B(n_175), .C(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_18), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_19), .B(n_475), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_20), .B(n_143), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_21), .B(n_287), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_22), .A2(n_205), .B(n_206), .C(n_208), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_23), .B(n_181), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_24), .B(n_158), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_25), .A2(n_177), .B(n_179), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_26), .B(n_158), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_27), .Y(n_229) );
INVx1_ASAP7_75t_L g217 ( .A(n_28), .Y(n_217) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_29), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_30), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_31), .B(n_158), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_32), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g460 ( .A(n_33), .Y(n_460) );
INVx1_ASAP7_75t_L g283 ( .A(n_34), .Y(n_283) );
INVx1_ASAP7_75t_L g525 ( .A(n_35), .Y(n_525) );
INVx2_ASAP7_75t_L g146 ( .A(n_36), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_37), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_38), .A2(n_205), .B(n_243), .C(n_245), .Y(n_242) );
INVxp67_ASAP7_75t_L g284 ( .A(n_39), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_40), .A2(n_153), .B(n_216), .C(n_222), .Y(n_215) );
CKINVDCx14_ASAP7_75t_R g241 ( .A(n_41), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_42), .A2(n_148), .B(n_153), .C(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g524 ( .A(n_44), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_45), .A2(n_157), .B(n_159), .C(n_162), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_46), .B(n_158), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_47), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_48), .Y(n_280) );
INVx1_ASAP7_75t_L g203 ( .A(n_49), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_50), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_51), .B(n_143), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_52), .A2(n_153), .B1(n_208), .B2(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_53), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_54), .Y(n_502) );
CKINVDCx14_ASAP7_75t_R g151 ( .A(n_55), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_56), .A2(n_157), .B(n_245), .C(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_57), .Y(n_562) );
INVx1_ASAP7_75t_L g514 ( .A(n_58), .Y(n_514) );
INVx1_ASAP7_75t_L g149 ( .A(n_59), .Y(n_149) );
INVx1_ASAP7_75t_L g140 ( .A(n_60), .Y(n_140) );
INVx1_ASAP7_75t_SL g244 ( .A(n_61), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_62), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_63), .B(n_181), .Y(n_210) );
INVx1_ASAP7_75t_L g232 ( .A(n_64), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_SL g533 ( .A1(n_65), .A2(n_245), .B(n_475), .C(n_534), .Y(n_533) );
INVxp67_ASAP7_75t_L g535 ( .A(n_66), .Y(n_535) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_68), .A2(n_143), .B(n_150), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_69), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_70), .A2(n_143), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_71), .Y(n_528) );
INVx1_ASAP7_75t_L g556 ( .A(n_72), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_73), .A2(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g173 ( .A(n_74), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_75), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_76), .A2(n_77), .B1(n_444), .B2(n_445), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_76), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_77), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_78), .A2(n_148), .B(n_153), .C(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_SL g451 ( .A1(n_79), .A2(n_122), .B1(n_452), .B2(n_745), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_143), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g176 ( .A(n_81), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_82), .B(n_218), .Y(n_473) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx1_ASAP7_75t_L g192 ( .A(n_84), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_85), .B(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_86), .A2(n_148), .B(n_153), .C(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g108 ( .A(n_87), .Y(n_108) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_88), .A2(n_153), .B(n_231), .C(n_234), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_89), .A2(n_91), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_89), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_90), .B(n_137), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_91), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_92), .A2(n_148), .B(n_153), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_93), .Y(n_488) );
INVx1_ASAP7_75t_L g532 ( .A(n_94), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_95), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_96), .B(n_218), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_97), .A2(n_105), .B1(n_114), .B2(n_750), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_98), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_99), .B(n_166), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g207 ( .A(n_101), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_102), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_102), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_103), .A2(n_143), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_106), .Y(n_751) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
INVx1_ASAP7_75t_L g743 ( .A(n_108), .Y(n_743) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_108), .B(n_122), .Y(n_747) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g123 ( .A(n_113), .B(n_124), .Y(n_123) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_450), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g749 ( .A(n_117), .Y(n_749) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_125), .B(n_447), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_121), .Y(n_449) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_130), .B2(n_446), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_126), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_127), .B(n_186), .Y(n_508) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
XOR2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_443), .Y(n_130) );
INVx2_ASAP7_75t_L g744 ( .A(n_131), .Y(n_744) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_373), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_288), .C(n_320), .D(n_337), .E(n_360), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_211), .B1(n_248), .B2(n_252), .C(n_256), .Y(n_133) );
INVx1_ASAP7_75t_L g400 ( .A(n_134), .Y(n_400) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_183), .Y(n_134) );
AND3x2_ASAP7_75t_L g375 ( .A(n_135), .B(n_185), .C(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_136), .B(n_254), .Y(n_253) );
BUFx3_ASAP7_75t_L g263 ( .A(n_136), .Y(n_263) );
AND2x2_ASAP7_75t_L g267 ( .A(n_136), .B(n_199), .Y(n_267) );
INVx2_ASAP7_75t_L g297 ( .A(n_136), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_136), .B(n_200), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_136), .B(n_184), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_136), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g387 ( .A(n_136), .B(n_200), .Y(n_387) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_142), .B(n_165), .Y(n_136) );
INVx1_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_137), .A2(n_189), .B(n_214), .C(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g237 ( .A(n_137), .Y(n_237) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_137), .A2(n_491), .B(n_497), .Y(n_490) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_L g167 ( .A(n_138), .B(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx2_ASAP7_75t_L g278 ( .A(n_143), .Y(n_278) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_144), .B(n_148), .Y(n_189) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx3_ASAP7_75t_L g161 ( .A(n_147), .Y(n_161) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g475 ( .A(n_147), .Y(n_475) );
INVx4_ASAP7_75t_SL g164 ( .A(n_148), .Y(n_164) );
BUFx3_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_164), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_152), .A2(n_164), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_152), .A2(n_164), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_152), .A2(n_164), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_152), .A2(n_164), .B(n_280), .C(n_281), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_152), .A2(n_164), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_152), .A2(n_164), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_152), .A2(n_164), .B(n_532), .C(n_533), .Y(n_531) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx5_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_161), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_161), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
INVx1_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_164), .A2(n_189), .B1(n_522), .B2(n_526), .Y(n_521) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_166), .Y(n_170) );
INVx4_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_166), .A2(n_530), .B(n_536), .Y(n_529) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g275 ( .A(n_167), .Y(n_275) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_168), .Y(n_266) );
AND2x2_ASAP7_75t_L g328 ( .A(n_168), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_168), .B(n_184), .Y(n_347) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g255 ( .A(n_169), .B(n_184), .Y(n_255) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_169), .Y(n_262) );
AND2x2_ASAP7_75t_L g314 ( .A(n_169), .B(n_200), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_169), .B(n_183), .C(n_297), .Y(n_339) );
AND2x2_ASAP7_75t_L g404 ( .A(n_169), .B(n_185), .Y(n_404) );
AND2x2_ASAP7_75t_L g438 ( .A(n_169), .B(n_184), .Y(n_438) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_180), .Y(n_169) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_170), .A2(n_201), .B(n_210), .Y(n_200) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_170), .A2(n_239), .B(n_247), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_177), .B(n_207), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_177), .A2(n_218), .B1(n_283), .B2(n_284), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_177), .B(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g523 ( .A1(n_178), .A2(n_194), .B1(n_524), .B2(n_525), .Y(n_523) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_181), .A2(n_512), .B(n_518), .Y(n_511) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_182), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_182), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_182), .A2(n_228), .B(n_235), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g476 ( .A(n_182), .B(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_184), .B(n_297), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_184), .B(n_328), .Y(n_336) );
AND2x2_ASAP7_75t_L g386 ( .A(n_184), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g414 ( .A(n_184), .Y(n_414) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g321 ( .A(n_185), .B(n_314), .Y(n_321) );
BUFx3_ASAP7_75t_L g353 ( .A(n_185), .Y(n_353) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_186), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_186), .B(n_562), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_189), .A2(n_229), .B(n_230), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_189), .A2(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_189), .A2(n_556), .B(n_557), .Y(n_555) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_193), .A2(n_196), .B(n_232), .C(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_196), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_196), .A2(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g329 ( .A(n_199), .Y(n_329) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_205), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g507 ( .A(n_208), .Y(n_507) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_211), .A2(n_389), .B1(n_391), .B2(n_392), .Y(n_388) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
AND2x2_ASAP7_75t_L g248 ( .A(n_212), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_SL g259 ( .A(n_212), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_212), .B(n_292), .Y(n_324) );
OR2x2_ASAP7_75t_L g343 ( .A(n_212), .B(n_226), .Y(n_343) );
AND2x2_ASAP7_75t_L g348 ( .A(n_212), .B(n_300), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_212), .B(n_293), .Y(n_351) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_238), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_212), .B(n_227), .Y(n_379) );
AND2x4_ASAP7_75t_L g382 ( .A(n_212), .B(n_250), .Y(n_382) );
OR2x2_ASAP7_75t_L g399 ( .A(n_212), .B(n_335), .Y(n_399) );
OR2x2_ASAP7_75t_L g430 ( .A(n_212), .B(n_272), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_212), .B(n_358), .Y(n_432) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .C(n_220), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_218), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_221), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g306 ( .A(n_225), .B(n_270), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_225), .B(n_293), .Y(n_425) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_238), .Y(n_225) );
AND2x2_ASAP7_75t_L g258 ( .A(n_226), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g292 ( .A(n_226), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_226), .B(n_272), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_226), .B(n_250), .Y(n_318) );
OR2x2_ASAP7_75t_L g335 ( .A(n_226), .B(n_293), .Y(n_335) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
BUFx2_ASAP7_75t_L g251 ( .A(n_227), .Y(n_251) );
AND2x2_ASAP7_75t_L g358 ( .A(n_227), .B(n_238), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_237), .A2(n_480), .B(n_487), .Y(n_479) );
INVx2_ASAP7_75t_L g250 ( .A(n_238), .Y(n_250) );
INVx1_ASAP7_75t_L g370 ( .A(n_238), .Y(n_370) );
AND2x2_ASAP7_75t_L g420 ( .A(n_238), .B(n_259), .Y(n_420) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_246), .Y(n_485) );
AND2x2_ASAP7_75t_L g269 ( .A(n_249), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g304 ( .A(n_249), .B(n_259), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_249), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g291 ( .A(n_250), .B(n_259), .Y(n_291) );
OR2x2_ASAP7_75t_L g407 ( .A(n_251), .B(n_381), .Y(n_407) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_254), .B(n_387), .Y(n_393) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OAI32xp33_ASAP7_75t_L g349 ( .A1(n_255), .A2(n_350), .A3(n_352), .B1(n_354), .B2(n_355), .Y(n_349) );
OR2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_308), .Y(n_366) );
OAI21xp33_ASAP7_75t_SL g391 ( .A1(n_255), .A2(n_265), .B(n_296), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B1(n_265), .B2(n_268), .Y(n_256) );
INVxp33_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_258), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_259), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g317 ( .A(n_259), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g417 ( .A(n_259), .B(n_358), .Y(n_417) );
OR2x2_ASAP7_75t_L g441 ( .A(n_259), .B(n_335), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_260), .A2(n_323), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_262), .B(n_267), .Y(n_319) );
AND2x2_ASAP7_75t_L g341 ( .A(n_263), .B(n_314), .Y(n_341) );
INVx1_ASAP7_75t_L g354 ( .A(n_263), .Y(n_354) );
OR2x2_ASAP7_75t_L g359 ( .A(n_263), .B(n_293), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_266), .B(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_267), .A2(n_290), .B1(n_295), .B2(n_299), .Y(n_289) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_270), .A2(n_332), .B1(n_339), .B2(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g416 ( .A(n_270), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_272), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g435 ( .A(n_272), .B(n_318), .Y(n_435) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_285), .Y(n_272) );
INVx1_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_273), .A2(n_555), .B(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI21xp5_ASAP7_75t_SL g469 ( .A1(n_274), .A2(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_275), .A2(n_501), .B(n_508), .Y(n_500) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_275), .A2(n_521), .B(n_527), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_275), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_277), .A2(n_286), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_301), .B1(n_302), .B2(n_307), .C(n_309), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_291), .B(n_293), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_291), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_292), .A2(n_398), .B(n_399), .C(n_400), .Y(n_397) );
AND2x2_ASAP7_75t_L g402 ( .A(n_292), .B(n_382), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_SL g440 ( .A1(n_292), .A2(n_381), .B(n_441), .C(n_442), .Y(n_440) );
BUFx3_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_296), .B(n_353), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_296), .A2(n_416), .B(n_418), .C(n_424), .Y(n_415) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVxp67_ASAP7_75t_L g376 ( .A(n_298), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_300), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
AOI211xp5_ASAP7_75t_L g320 ( .A1(n_304), .A2(n_321), .B(n_322), .C(n_330), .Y(n_320) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g405 ( .A(n_308), .Y(n_405) );
OR2x2_ASAP7_75t_L g422 ( .A(n_308), .B(n_352), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_316), .B2(n_319), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_311), .A2(n_323), .B1(n_324), .B2(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
OR2x2_ASAP7_75t_L g409 ( .A(n_313), .B(n_353), .Y(n_409) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g364 ( .A(n_314), .B(n_354), .Y(n_364) );
INVx1_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_318), .B(n_332), .Y(n_380) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_328), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g437 ( .A(n_329), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_332), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_332), .B(n_363), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_332), .B(n_358), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_332), .B(n_379), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g394 ( .A1(n_332), .A2(n_342), .B(n_382), .C(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_342), .B1(n_344), .B2(n_348), .C(n_349), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_346), .B(n_354), .Y(n_428) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_348), .A2(n_363), .B(n_365), .C(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_351), .B(n_358), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_352), .B(n_405), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
INVxp33_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_357), .A2(n_369), .B(n_371), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_357), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_358), .B(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B1(n_365), .B2(n_367), .C(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_364), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
NAND5xp2_ASAP7_75t_L g373 ( .A(n_374), .B(n_401), .C(n_415), .D(n_426), .E(n_439), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_384), .C(n_397), .Y(n_374) );
INVx2_ASAP7_75t_SL g421 ( .A(n_375), .Y(n_421) );
NAND4xp25_ASAP7_75t_SL g377 ( .A(n_378), .B(n_380), .C(n_381), .D(n_383), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_383), .A2(n_385), .B(n_388), .C(n_394), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_386), .A2(n_427), .B1(n_429), .B2(n_431), .C(n_433), .Y(n_426) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_409), .A2(n_432), .B1(n_434), .B2(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_447), .B(n_451), .C(n_748), .Y(n_450) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
XOR2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_711), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_604), .C(n_677), .Y(n_464) );
OAI211xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_498), .B(n_537), .C(n_588), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g553 ( .A(n_468), .B(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g571 ( .A(n_468), .Y(n_571) );
INVx2_ASAP7_75t_L g586 ( .A(n_468), .Y(n_586) );
INVx1_ASAP7_75t_L g616 ( .A(n_468), .Y(n_616) );
AND2x2_ASAP7_75t_L g666 ( .A(n_468), .B(n_587), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g693 ( .A1(n_468), .A2(n_621), .A3(n_694), .B1(n_696), .B2(n_697), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_468), .B(n_543), .Y(n_699) );
AND2x2_ASAP7_75t_L g726 ( .A(n_468), .B(n_569), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_468), .B(n_735), .Y(n_734) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_476), .Y(n_468) );
AND2x2_ASAP7_75t_L g615 ( .A(n_478), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g637 ( .A(n_478), .Y(n_637) );
AND2x2_ASAP7_75t_L g722 ( .A(n_478), .B(n_553), .Y(n_722) );
AND2x2_ASAP7_75t_L g725 ( .A(n_478), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
INVx2_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_479), .B(n_569), .Y(n_575) );
AND2x2_ASAP7_75t_L g585 ( .A(n_479), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g621 ( .A(n_479), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_486), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_485), .Y(n_482) );
AND2x2_ASAP7_75t_L g563 ( .A(n_489), .B(n_545), .Y(n_563) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g546 ( .A(n_490), .Y(n_546) );
AND2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_569), .Y(n_587) );
AND2x2_ASAP7_75t_L g656 ( .A(n_490), .B(n_554), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
OR2x2_ASAP7_75t_L g551 ( .A(n_499), .B(n_520), .Y(n_551) );
INVx1_ASAP7_75t_L g629 ( .A(n_499), .Y(n_629) );
AND2x2_ASAP7_75t_L g643 ( .A(n_499), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_499), .B(n_519), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_499), .B(n_641), .Y(n_695) );
AND2x2_ASAP7_75t_L g703 ( .A(n_499), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g541 ( .A(n_500), .Y(n_541) );
AND2x2_ASAP7_75t_L g610 ( .A(n_500), .B(n_520), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_509), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g737 ( .A(n_509), .Y(n_737) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_510), .B(n_581), .Y(n_603) );
OR2x2_ASAP7_75t_L g632 ( .A(n_510), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g664 ( .A(n_510), .B(n_644), .Y(n_664) );
INVx1_ASAP7_75t_SL g684 ( .A(n_510), .Y(n_684) );
AND2x2_ASAP7_75t_L g688 ( .A(n_510), .B(n_550), .Y(n_688) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_511), .B(n_519), .Y(n_542) );
AND2x2_ASAP7_75t_L g549 ( .A(n_511), .B(n_529), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g591 ( .A(n_511), .B(n_573), .Y(n_591) );
INVx1_ASAP7_75t_SL g598 ( .A(n_511), .Y(n_598) );
BUFx2_ASAP7_75t_L g609 ( .A(n_511), .Y(n_609) );
AND2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_541), .Y(n_625) );
AND2x2_ASAP7_75t_L g640 ( .A(n_511), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g704 ( .A(n_511), .B(n_520), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_519), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g628 ( .A(n_519), .B(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_519), .A2(n_646), .B1(n_649), .B2(n_652), .C(n_657), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_519), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
INVx3_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
BUFx2_ASAP7_75t_L g583 ( .A(n_529), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_529), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g614 ( .A(n_529), .Y(n_614) );
OR2x2_ASAP7_75t_L g633 ( .A(n_529), .B(n_573), .Y(n_633) );
INVx3_ASAP7_75t_L g641 ( .A(n_529), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_529), .B(n_573), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_543), .B1(n_547), .B2(n_552), .C(n_564), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_540), .B(n_613), .Y(n_738) );
OR2x2_ASAP7_75t_L g741 ( .A(n_540), .B(n_572), .Y(n_741) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_541), .A2(n_565), .B1(n_572), .B2(n_574), .C(n_577), .Y(n_564) );
AND2x2_ASAP7_75t_L g581 ( .A(n_541), .B(n_573), .Y(n_581) );
AND2x2_ASAP7_75t_L g589 ( .A(n_541), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_541), .B(n_597), .Y(n_596) );
NAND2x1_ASAP7_75t_L g639 ( .A(n_541), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g691 ( .A(n_541), .B(n_633), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_543), .A2(n_651), .B1(n_680), .B2(n_682), .Y(n_679) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI322xp5_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_553), .A3(n_589), .B1(n_592), .B2(n_595), .C1(n_599), .C2(n_602), .Y(n_588) );
OR2x2_ASAP7_75t_L g600 ( .A(n_544), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_545), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g579 ( .A(n_545), .B(n_554), .Y(n_579) );
INVx1_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
AND2x2_ASAP7_75t_L g660 ( .A(n_545), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g570 ( .A(n_546), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g661 ( .A(n_546), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_546), .B(n_569), .Y(n_735) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_550), .B(n_684), .Y(n_683) );
INVx3_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g635 ( .A(n_551), .B(n_582), .Y(n_635) );
OR2x2_ASAP7_75t_L g732 ( .A(n_551), .B(n_583), .Y(n_732) );
INVx1_ASAP7_75t_L g713 ( .A(n_552), .Y(n_713) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_563), .Y(n_552) );
INVx4_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_553), .B(n_620), .Y(n_626) );
INVx2_ASAP7_75t_L g569 ( .A(n_554), .Y(n_569) );
INVx1_ASAP7_75t_L g651 ( .A(n_563), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_563), .B(n_623), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g638 ( .A1(n_565), .A2(n_639), .B(n_642), .Y(n_638) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g623 ( .A(n_569), .Y(n_623) );
INVx1_ASAP7_75t_L g650 ( .A(n_569), .Y(n_650) );
INVx1_ASAP7_75t_L g576 ( .A(n_570), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_570), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g674 ( .A(n_571), .B(n_660), .Y(n_674) );
AND2x2_ASAP7_75t_L g696 ( .A(n_571), .B(n_656), .Y(n_696) );
BUFx2_ASAP7_75t_L g648 ( .A(n_573), .Y(n_648) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AOI32xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .A3(n_581), .B1(n_582), .B2(n_584), .Y(n_577) );
INVx1_ASAP7_75t_L g658 ( .A(n_578), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_578), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_581), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_581), .B(n_640), .Y(n_681) );
AND2x2_ASAP7_75t_L g728 ( .A(n_581), .B(n_613), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_582), .B(n_629), .Y(n_676) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g729 ( .A(n_584), .Y(n_729) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g654 ( .A(n_585), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_587), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g701 ( .A(n_587), .B(n_621), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_587), .B(n_616), .Y(n_708) );
INVx1_ASAP7_75t_SL g690 ( .A(n_589), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_590), .B(n_641), .Y(n_668) );
NOR4xp25_ASAP7_75t_L g714 ( .A(n_590), .B(n_613), .C(n_715), .D(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_591), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_L g671 ( .A(n_594), .Y(n_671) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_597), .A2(n_688), .B(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g613 ( .A(n_598), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g662 ( .A(n_601), .Y(n_662) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND4xp25_ASAP7_75t_SL g604 ( .A(n_605), .B(n_630), .C(n_645), .D(n_665), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_611), .B(n_615), .C(n_617), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g697 ( .A(n_610), .B(n_640), .Y(n_697) );
AND2x2_ASAP7_75t_L g706 ( .A(n_610), .B(n_684), .Y(n_706) );
INVx3_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_613), .B(n_648), .Y(n_710) );
AND2x2_ASAP7_75t_L g622 ( .A(n_616), .B(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_624), .B1(n_626), .B2(n_627), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g720 ( .A(n_620), .B(n_666), .Y(n_720) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_622), .B(n_671), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_623), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_636), .C(n_638), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_631), .A2(n_666), .B1(n_667), .B2(n_669), .C(n_672), .Y(n_665) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_639), .A2(n_724), .B1(n_727), .B2(n_729), .C(n_730), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_640), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_648), .B(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g678 ( .A(n_650), .Y(n_678) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_653), .A2(n_673), .B1(n_675), .B2(n_676), .Y(n_672) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_662), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_673), .A2(n_699), .B1(n_737), .B2(n_738), .C(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g718 ( .A(n_675), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_685), .C(n_705), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_689), .C(n_698), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B(n_692), .C(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g717 ( .A(n_695), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_696), .A2(n_722), .B(n_740), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g731 ( .A1(n_708), .A2(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_723), .C(n_736), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_719), .C(n_721), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
CKINVDCx14_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule