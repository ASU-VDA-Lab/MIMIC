module fake_jpeg_6662_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx11_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_18),
.B(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_9),
.B1(n_8),
.B2(n_12),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_24),
.B(n_25),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_6),
.B(n_10),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_9),
.C(n_12),
.Y(n_25)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_10),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_33),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_9),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_25),
.B(n_6),
.Y(n_37)
);

NOR4xp25_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.C(n_11),
.D(n_36),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_7),
.B1(n_11),
.B2(n_34),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_11),
.B(n_31),
.Y(n_40)
);


endmodule