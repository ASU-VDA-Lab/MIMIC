module fake_jpeg_3721_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_13;
wire n_21;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_27),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_17),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_39),
.B1(n_23),
.B2(n_18),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_59),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_14),
.B(n_24),
.C(n_33),
.D(n_15),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_16),
.A3(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_61),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_18),
.Y(n_59)
);

OR2x4_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_24),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_79),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_47),
.A3(n_25),
.B1(n_26),
.B2(n_43),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_23),
.B(n_36),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_28),
.B1(n_31),
.B2(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_39),
.B1(n_61),
.B2(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_50),
.B1(n_57),
.B2(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_101),
.B1(n_102),
.B2(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_95),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_64),
.B1(n_62),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_104),
.B1(n_41),
.B2(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_23),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_26),
.B(n_25),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_44),
.B1(n_54),
.B2(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_65),
.B1(n_63),
.B2(n_43),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_119),
.B1(n_81),
.B2(n_30),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_80),
.B1(n_67),
.B2(n_63),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_124),
.B1(n_103),
.B2(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_80),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_114),
.C(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_46),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_48),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_101),
.C(n_48),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_98),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_81),
.B1(n_83),
.B2(n_36),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_95),
.B(n_115),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_131),
.B(n_139),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_134),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_146),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_20),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_103),
.B1(n_86),
.B2(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_96),
.B1(n_89),
.B2(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_94),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_99),
.B(n_94),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_138),
.B(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_118),
.C(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_110),
.B1(n_41),
.B2(n_72),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_154),
.C(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_157),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_128),
.B1(n_146),
.B2(n_129),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_123),
.C(n_72),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_72),
.C(n_30),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_160),
.B1(n_165),
.B2(n_130),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_166),
.Y(n_179)
);

AO21x2_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_24),
.B(n_16),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_24),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_164),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_24),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_16),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_24),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_22),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_0),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_147),
.B1(n_143),
.B2(n_145),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_173),
.B1(n_170),
.B2(n_160),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_184),
.B(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_141),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_135),
.B1(n_136),
.B2(n_140),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_145),
.B1(n_131),
.B2(n_127),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_141),
.C(n_16),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_164),
.C(n_161),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_16),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_165),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_163),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_166),
.C(n_159),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_201),
.B(n_22),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_200),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_158),
.B(n_154),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_199),
.B(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_182),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_160),
.B1(n_169),
.B2(n_152),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_162),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_180),
.C(n_179),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_161),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.C(n_191),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_184),
.C(n_179),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_215),
.B(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_184),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_225),
.B1(n_13),
.B2(n_201),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_26),
.C(n_25),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_26),
.C(n_25),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_21),
.B(n_19),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_13),
.B(n_21),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_230),
.C(n_236),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_203),
.C(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_11),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_1),
.B(n_2),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_226),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_1),
.B(n_2),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_214),
.B(n_3),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_212),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_224),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_252),
.B(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_251),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_234),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_3),
.C(n_4),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_4),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_4),
.C(n_5),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_4),
.B(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_259),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_263),
.B(n_6),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_228),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_232),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_7),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_5),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_7),
.Y(n_270)
);

AOI221xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_243),
.B1(n_260),
.B2(n_255),
.C(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_5),
.B(n_6),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_269),
.B(n_271),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_7),
.C(n_8),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_266),
.B(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_7),
.C(n_8),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_9),
.B1(n_10),
.B2(n_277),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_280),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_9),
.B(n_10),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_278),
.Y(n_284)
);


endmodule