module real_jpeg_15723_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_6),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_2),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_3),
.A2(n_108),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_3),
.A2(n_108),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_4),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_183),
.B1(n_187),
.B2(n_192),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_7),
.Y(n_169)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_7),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_7),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_8),
.A2(n_171),
.B1(n_175),
.B2(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_178),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_9),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_9),
.Y(n_309)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_9),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_10),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_107),
.B1(n_141),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_10),
.A2(n_141),
.B1(n_184),
.B2(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_194),
.A3(n_197),
.B1(n_201),
.B2(n_208),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_12),
.B(n_27),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_12),
.A2(n_284),
.A3(n_288),
.B1(n_289),
.B2(n_292),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_12),
.A2(n_56),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_12),
.B(n_67),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_12),
.B(n_395),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_12),
.B(n_148),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_13),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_13),
.A2(n_60),
.B1(n_235),
.B2(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_13),
.A2(n_60),
.B1(n_357),
.B2(n_363),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_13),
.A2(n_60),
.B1(n_397),
.B2(n_401),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_15),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_15),
.A2(n_150),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_16),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

BUFx4f_ASAP7_75t_L g174 ( 
.A(n_16),
.Y(n_174)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_16),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_278),
.B1(n_428),
.B2(n_429),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_21),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_277),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_243),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_23),
.B(n_243),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_158),
.C(n_214),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_24),
.B(n_424),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_64),
.Y(n_24)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_25),
.B(n_65),
.C(n_116),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_48),
.B1(n_57),
.B2(n_63),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_26),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_27),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_27)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_28),
.Y(n_321)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_29),
.Y(n_240)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_50),
.Y(n_252)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_55),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_56),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_56),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_56),
.B(n_129),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_56),
.A2(n_344),
.B(n_354),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_56),
.A2(n_162),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_57),
.Y(n_247)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_62),
.A2(n_100),
.B1(n_104),
.B2(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_116),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_95),
.B1(n_105),
.B2(n_115),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_66),
.Y(n_241)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_66),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_66),
.A2(n_115),
.B1(n_234),
.B2(n_315),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_80),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_73),
.Y(n_291)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_75),
.Y(n_270)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_76),
.Y(n_274)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_95),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_100),
.A2(n_104),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_100),
.A2(n_104),
.B1(n_187),
.B2(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_103),
.Y(n_259)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_112),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_115),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_115),
.B(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_147),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_117),
.A2(n_130),
.B1(n_303),
.B2(n_310),
.Y(n_302)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_118),
.B(n_149),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_118),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_118),
.A2(n_148),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_118),
.A2(n_148),
.B1(n_304),
.B2(n_356),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_130),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_123),
.B1(n_125),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_121),
.Y(n_339)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_122),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_122),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_124),
.Y(n_343)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_129),
.Y(n_313)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_130),
.B(n_138),
.Y(n_327)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_133),
.Y(n_350)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_145),
.Y(n_288)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_148),
.B(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_158),
.A2(n_159),
.B1(n_214),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_193),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_160),
.B(n_193),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_170),
.B1(n_179),
.B2(n_182),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_161),
.A2(n_182),
.B(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_161),
.A2(n_264),
.B(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_161),
.A2(n_383),
.B1(n_387),
.B2(n_388),
.Y(n_382)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_162),
.A2(n_367),
.B(n_373),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_162),
.A2(n_384),
.B1(n_396),
.B2(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_167),
.B(n_222),
.Y(n_264)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_168),
.Y(n_411)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_216),
.B(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_173),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_174),
.Y(n_370)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_174),
.Y(n_400)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_185),
.Y(n_372)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_185),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_189),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_214),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_231),
.C(n_233),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_215),
.A2(n_231),
.B1(n_232),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g376 ( 
.A(n_219),
.Y(n_376)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_219),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_233),
.B(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_261),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_260),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_278),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_422),
.B(n_427),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_333),
.B(n_421),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_322),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_281),
.B(n_322),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_302),
.C(n_314),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_282),
.B(n_419),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_298),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_298),
.Y(n_324)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_300),
.B(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_302),
.B(n_314),
.Y(n_419)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_328),
.B1(n_329),
.B2(n_332),
.Y(n_322)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_324),
.B(n_325),
.C(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_416),
.B(n_420),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_380),
.B(n_415),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_365),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_336),
.B(n_365),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_351),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_337),
.A2(n_351),
.B1(n_352),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_340),
.A3(n_341),
.B1(n_344),
.B2(n_345),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_377),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_378),
.C(n_379),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

OAI21x1_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_391),
.B(n_414),
.Y(n_380)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_389),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_389),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_407),
.B(n_413),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_402),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_412),
.Y(n_413)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_417),
.B(n_418),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_426),
.Y(n_427)
);


endmodule