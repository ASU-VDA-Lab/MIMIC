module fake_netlist_5_15_n_1743 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1743);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1743;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_83),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_54),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_40),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_46),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_26),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_33),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_21),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_16),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_53),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_105),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_22),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_102),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_118),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_35),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_43),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_35),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_146),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_106),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_28),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_61),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_81),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_37),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_73),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_30),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_34),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_4),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_20),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_94),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_8),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_38),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_53),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_87),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_101),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_67),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_92),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_153),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_141),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_57),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_58),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_21),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_32),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_129),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_52),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_12),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_16),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_124),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_29),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_38),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_89),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_10),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_45),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_26),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_98),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_69),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_96),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_14),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_17),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_127),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_10),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_60),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_41),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_80),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_46),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_48),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_64),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_70),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_44),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_123),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_32),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_72),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_22),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_29),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_132),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_45),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_82),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_56),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_66),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_156),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_171),
.B(n_0),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_196),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_157),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_158),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_167),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_175),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_179),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_205),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_208),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_165),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_180),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_302),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_219),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_186),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_188),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_267),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_242),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_192),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_198),
.B(n_0),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_202),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_211),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_276),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_204),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_214),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_215),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_287),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_216),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_290),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_173),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_191),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_222),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_191),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_240),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_178),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_174),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_288),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_198),
.B(n_1),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_240),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_220),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_241),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_221),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_159),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_163),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_163),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_166),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_231),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_192),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_166),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_234),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_189),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_189),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_194),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_224),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_224),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_244),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_334),
.A2(n_164),
.B1(n_252),
.B2(n_274),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_348),
.B(n_244),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_353),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_312),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_358),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_348),
.B(n_243),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_245),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_246),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_348),
.B(n_247),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_321),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_323),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_383),
.B(n_160),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_383),
.B(n_160),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_168),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_323),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_329),
.Y(n_442)
);

AND3x2_ASAP7_75t_L g443 ( 
.A(n_371),
.B(n_218),
.C(n_233),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_329),
.A2(n_203),
.B(n_194),
.Y(n_445)
);

AND2x4_ASAP7_75t_SL g446 ( 
.A(n_377),
.B(n_239),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_325),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_338),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_338),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_350),
.B(n_345),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_168),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_339),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_170),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_366),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_394),
.B(n_331),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_412),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_319),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_310),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_336),
.B1(n_316),
.B2(n_343),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_445),
.A2(n_313),
.B1(n_303),
.B2(n_251),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_394),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_417),
.B(n_320),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_203),
.B1(n_206),
.B2(n_209),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_430),
.B(n_324),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_327),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_170),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_176),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_445),
.A2(n_438),
.B1(n_439),
.B2(n_435),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

AND3x2_ASAP7_75t_L g490 ( 
.A(n_421),
.B(n_177),
.C(n_176),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_419),
.B(n_328),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_430),
.B(n_330),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_394),
.B(n_335),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_435),
.B(n_438),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_411),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_395),
.B(n_372),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_419),
.B(n_337),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_395),
.B(n_341),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_408),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_427),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_436),
.B(n_344),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_400),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_404),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_446),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_411),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_406),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_395),
.B(n_351),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_427),
.B(n_355),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_400),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_436),
.B(n_356),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_447),
.A2(n_353),
.B1(n_370),
.B2(n_184),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_436),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_416),
.B(n_375),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_396),
.B(n_230),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_390),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_440),
.B(n_206),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

AND3x2_ASAP7_75t_L g547 ( 
.A(n_421),
.B(n_182),
.C(n_177),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_376),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_446),
.B(n_182),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_440),
.A2(n_362),
.B1(n_360),
.B2(n_357),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_390),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_425),
.B(n_373),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_408),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_390),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_402),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_396),
.B(n_230),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_447),
.B(n_385),
.C(n_382),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_425),
.B(n_386),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_390),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_425),
.B(n_193),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_438),
.A2(n_270),
.B1(n_209),
.B2(n_303),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_446),
.B(n_370),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_408),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_402),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_390),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_443),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_439),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_446),
.B(n_248),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_413),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_443),
.B(n_210),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_406),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_461),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_456),
.B(n_293),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_415),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_402),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_439),
.B(n_184),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_461),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_439),
.B(n_250),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_461),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_455),
.B(n_253),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_433),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_415),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_433),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_418),
.B(n_376),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_433),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_456),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_401),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_441),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_441),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_254),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_455),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_449),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_455),
.B(n_255),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_415),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_262),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_415),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_458),
.B(n_212),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_405),
.A2(n_259),
.B1(n_197),
.B2(n_195),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_474),
.B(n_468),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_482),
.A2(n_227),
.B1(n_298),
.B2(n_270),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_475),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_509),
.B(n_458),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_474),
.B(n_317),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_488),
.B(n_458),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_466),
.B(n_301),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_510),
.B(n_318),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_576),
.B(n_162),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_476),
.B(n_458),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_415),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_572),
.B(n_183),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_579),
.B(n_401),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_535),
.B(n_549),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_538),
.B(n_332),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_504),
.B(n_420),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_491),
.B(n_415),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_506),
.B(n_415),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_563),
.A2(n_405),
.B(n_449),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_549),
.B(n_340),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_531),
.B(n_415),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_486),
.A2(n_449),
.B(n_429),
.Y(n_635)
);

BUFx8_ASAP7_75t_L g636 ( 
.A(n_538),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_493),
.B(n_185),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_529),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_471),
.B(n_199),
.C(n_187),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_507),
.B(n_201),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_477),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_550),
.B(n_346),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_481),
.B(n_429),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_467),
.B(n_354),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_529),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

INVx8_ASAP7_75t_L g648 ( 
.A(n_501),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_481),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_484),
.B(n_429),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_420),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_473),
.B(n_359),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_484),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_559),
.B(n_361),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_486),
.B(n_429),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_525),
.B(n_207),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_552),
.B(n_265),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_479),
.B(n_213),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_560),
.B(n_429),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_492),
.B(n_228),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_565),
.B(n_212),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_482),
.B(n_190),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_423),
.Y(n_664)
);

BUFx5_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_555),
.B(n_190),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_472),
.B(n_429),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_523),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_472),
.B(n_429),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_536),
.B(n_271),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_539),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_472),
.B(n_278),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_541),
.B(n_429),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_391),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_551),
.B(n_391),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_534),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_551),
.B(n_392),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_543),
.B(n_229),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_543),
.B(n_232),
.Y(n_681)
);

INVx8_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_543),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_554),
.B(n_392),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_548),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_554),
.B(n_295),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_487),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_467),
.Y(n_688)
);

AND2x4_ASAP7_75t_SL g689 ( 
.A(n_516),
.B(n_239),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_562),
.B(n_397),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_610),
.B(n_256),
.C(n_299),
.Y(n_692)
);

O2A1O1Ixp5_ASAP7_75t_L g693 ( 
.A1(n_483),
.A2(n_414),
.B(n_397),
.C(n_403),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_562),
.B(n_297),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_485),
.Y(n_695)
);

AO21x1_ASAP7_75t_L g696 ( 
.A1(n_470),
.A2(n_200),
.B(n_256),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_564),
.B(n_478),
.C(n_608),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_485),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_516),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_608),
.B(n_237),
.C(n_249),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_592),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_555),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_569),
.B(n_403),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_558),
.B(n_407),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_558),
.B(n_407),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_586),
.A2(n_305),
.B1(n_304),
.B2(n_226),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_485),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_483),
.B(n_409),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_483),
.B(n_495),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_604),
.A2(n_223),
.B1(n_200),
.B2(n_294),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_528),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_561),
.B(n_423),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_596),
.B(n_236),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_561),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_566),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_495),
.B(n_409),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_566),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_570),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_577),
.B(n_424),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_495),
.B(n_410),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_SL g722 ( 
.A(n_574),
.B(n_172),
.C(n_238),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_502),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_502),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_503),
.B(n_424),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_501),
.B(n_230),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_502),
.B(n_410),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_512),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_512),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_587),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_512),
.B(n_414),
.Y(n_731)
);

INVx4_ASAP7_75t_SL g732 ( 
.A(n_501),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_570),
.B(n_223),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_573),
.A2(n_226),
.B1(n_299),
.B2(n_272),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_584),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_573),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_490),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_501),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_470),
.B(n_217),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_465),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_601),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_516),
.B(n_426),
.Y(n_742)
);

INVx8_ASAP7_75t_L g743 ( 
.A(n_503),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_487),
.B(n_230),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_470),
.B(n_459),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_588),
.B(n_426),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_465),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_600),
.B(n_257),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_601),
.A2(n_285),
.B1(n_275),
.B2(n_272),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_601),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_606),
.B(n_459),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_522),
.B(n_428),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_522),
.B(n_428),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_601),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_464),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_584),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_497),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_497),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_513),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_513),
.B(n_258),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_568),
.B(n_459),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_568),
.B(n_459),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_515),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_568),
.B(n_459),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_553),
.A2(n_463),
.B(n_462),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_527),
.B(n_260),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_459),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_487),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_527),
.A2(n_275),
.B1(n_294),
.B2(n_285),
.Y(n_769)
);

OAI221xp5_ASAP7_75t_L g770 ( 
.A1(n_540),
.A2(n_217),
.B1(n_225),
.B2(n_227),
.C(n_251),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_532),
.B(n_261),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_532),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_614),
.A2(n_567),
.B(n_553),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_SL g774 ( 
.A(n_688),
.B(n_578),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_748),
.B(n_533),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_625),
.A2(n_557),
.B(n_540),
.C(n_537),
.Y(n_777)
);

AOI21x1_ASAP7_75t_L g778 ( 
.A1(n_635),
.A2(n_542),
.B(n_537),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_621),
.A2(n_616),
.B(n_745),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_641),
.B(n_544),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_649),
.B(n_544),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_653),
.B(n_545),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_668),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_627),
.B(n_546),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_757),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_627),
.B(n_546),
.Y(n_787)
);

BUFx8_ASAP7_75t_SL g788 ( 
.A(n_699),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_658),
.B(n_578),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_743),
.Y(n_791)
);

AOI21xp33_ASAP7_75t_L g792 ( 
.A1(n_659),
.A2(n_557),
.B(n_264),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_622),
.A2(n_567),
.B(n_553),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_715),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_665),
.B(n_464),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_758),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_720),
.B(n_547),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_671),
.B(n_590),
.Y(n_798)
);

AOI33xp33_ASAP7_75t_L g799 ( 
.A1(n_664),
.A2(n_389),
.A3(n_225),
.B1(n_284),
.B2(n_282),
.B3(n_298),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_676),
.B(n_590),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_SL g801 ( 
.A(n_644),
.B(n_280),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_685),
.B(n_607),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_607),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_628),
.A2(n_567),
.B(n_517),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_759),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_612),
.A2(n_284),
.B(n_282),
.C(n_286),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_701),
.B(n_607),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_743),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_629),
.A2(n_505),
.B(n_605),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_434),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_634),
.A2(n_505),
.B(n_605),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_660),
.A2(n_505),
.B(n_605),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_617),
.B(n_571),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_763),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_635),
.A2(n_609),
.B(n_575),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_652),
.A2(n_487),
.B1(n_583),
.B2(n_602),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_665),
.B(n_487),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_617),
.B(n_571),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_655),
.A2(n_520),
.B(n_580),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_730),
.B(n_434),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_658),
.B(n_239),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_665),
.B(n_738),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_679),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_751),
.A2(n_580),
.B(n_520),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_647),
.B(n_575),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_665),
.B(n_464),
.Y(n_827)
);

AO21x2_ASAP7_75t_L g828 ( 
.A1(n_696),
.A2(n_609),
.B(n_582),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_753),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_582),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_611),
.B(n_589),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_693),
.A2(n_595),
.B(n_602),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_692),
.A2(n_595),
.B(n_599),
.C(n_598),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_709),
.A2(n_517),
.B(n_520),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_693),
.A2(n_593),
.B(n_599),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_665),
.B(n_464),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_687),
.A2(n_580),
.B(n_517),
.Y(n_837)
);

NOR2x1_ASAP7_75t_L g838 ( 
.A(n_725),
.B(n_589),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_760),
.B(n_593),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_665),
.B(n_464),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_673),
.A2(n_496),
.B(n_499),
.Y(n_841)
);

AO21x1_ASAP7_75t_L g842 ( 
.A1(n_663),
.A2(n_598),
.B(n_277),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_612),
.A2(n_286),
.B(n_277),
.C(n_454),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_626),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_651),
.B(n_437),
.Y(n_845)
);

CKINVDCx10_ASAP7_75t_R g846 ( 
.A(n_699),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_760),
.B(n_766),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_667),
.A2(n_500),
.B(n_499),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_738),
.B(n_496),
.Y(n_849)
);

INVx11_ASAP7_75t_L g850 ( 
.A(n_636),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_437),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_669),
.A2(n_556),
.B(n_500),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_714),
.B(n_444),
.Y(n_853)
);

INVx11_ASAP7_75t_L g854 ( 
.A(n_636),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_692),
.A2(n_697),
.B(n_661),
.C(n_659),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_585),
.Y(n_856)
);

AO21x2_ASAP7_75t_L g857 ( 
.A1(n_630),
.A2(n_726),
.B(n_702),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_744),
.B(n_389),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_715),
.B(n_496),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_755),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_661),
.A2(n_444),
.B(n_451),
.C(n_454),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_732),
.B(n_496),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_771),
.B(n_603),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_746),
.A2(n_556),
.B(n_500),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_732),
.B(n_496),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_620),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_742),
.B(n_451),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_771),
.B(n_603),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_698),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_643),
.A2(n_581),
.B(n_499),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_624),
.B(n_585),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_615),
.B(n_591),
.Y(n_872)
);

NAND2x1_ASAP7_75t_L g873 ( 
.A(n_755),
.B(n_499),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_650),
.A2(n_556),
.B(n_500),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_712),
.B(n_597),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_716),
.B(n_597),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_722),
.B(n_591),
.Y(n_877)
);

NOR2x1p5_ASAP7_75t_SL g878 ( 
.A(n_707),
.B(n_469),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_715),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_630),
.A2(n_498),
.B(n_469),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_755),
.A2(n_500),
.B(n_581),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_718),
.B(n_487),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_739),
.A2(n_663),
.B1(n_682),
.B2(n_648),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_719),
.B(n_487),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_768),
.B(n_499),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_772),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_736),
.B(n_583),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_741),
.A2(n_583),
.B1(n_581),
.B2(n_556),
.Y(n_889)
);

NOR2x1_ASAP7_75t_R g890 ( 
.A(n_642),
.B(n_266),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_623),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_770),
.A2(n_489),
.B(n_519),
.C(n_514),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_755),
.A2(n_581),
.B(n_556),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_769),
.A2(n_489),
.B(n_519),
.C(n_514),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_723),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_674),
.A2(n_581),
.B(n_521),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_724),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_675),
.A2(n_521),
.B(n_518),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_743),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_623),
.B(n_583),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_651),
.B(n_583),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_708),
.A2(n_494),
.B(n_511),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_728),
.Y(n_903)
);

BUFx2_ASAP7_75t_SL g904 ( 
.A(n_711),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_678),
.A2(n_521),
.B(n_518),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_713),
.B(n_583),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_637),
.A2(n_268),
.B(n_269),
.C(n_273),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_729),
.Y(n_908)
);

NOR2x1p5_ASAP7_75t_L g909 ( 
.A(n_722),
.B(n_279),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_749),
.A2(n_494),
.B(n_511),
.C(n_498),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_684),
.A2(n_521),
.B(n_518),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_691),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_703),
.A2(n_521),
.B(n_518),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_761),
.A2(n_518),
.B(n_508),
.Y(n_914)
);

AOI21xp33_ASAP7_75t_L g915 ( 
.A1(n_637),
.A2(n_281),
.B(n_289),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_733),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_762),
.A2(n_764),
.B(n_682),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_739),
.A2(n_583),
.B(n_526),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_670),
.A2(n_463),
.B(n_462),
.C(n_457),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_648),
.A2(n_526),
.B(n_508),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_735),
.B(n_291),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_640),
.B(n_452),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_739),
.A2(n_300),
.B1(n_292),
.B2(n_307),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_SL g924 ( 
.A1(n_640),
.A2(n_452),
.B(n_453),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_648),
.A2(n_526),
.B(n_508),
.Y(n_925)
);

NOR2x1p5_ASAP7_75t_L g926 ( 
.A(n_639),
.B(n_296),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_682),
.A2(n_526),
.B(n_508),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_767),
.A2(n_526),
.B(n_508),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_677),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_656),
.B(n_452),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_750),
.A2(n_754),
.B(n_672),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_679),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_756),
.B(n_311),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_656),
.B(n_452),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_230),
.B1(n_453),
.B2(n_463),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_657),
.B(n_453),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_680),
.B(n_453),
.C(n_463),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_704),
.A2(n_705),
.B(n_717),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_710),
.B(n_462),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_721),
.B(n_462),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_727),
.A2(n_526),
.B(n_508),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_731),
.A2(n_457),
.B(n_459),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_686),
.A2(n_457),
.B(n_459),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_457),
.B(n_230),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_732),
.B(n_230),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_694),
.A2(n_460),
.B(n_230),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_619),
.B(n_1),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_756),
.B(n_680),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_L g949 ( 
.A(n_733),
.B(n_230),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_737),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_618),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_683),
.B(n_700),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_460),
.B(n_65),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_631),
.A2(n_460),
.B(n_68),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_638),
.B(n_645),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_646),
.A2(n_460),
.B(n_155),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_784),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_779),
.A2(n_818),
.B(n_837),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_845),
.B(n_683),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_847),
.A2(n_733),
.B1(n_632),
.B2(n_666),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_855),
.A2(n_681),
.B(n_706),
.C(n_752),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_845),
.B(n_662),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_778),
.A2(n_917),
.B(n_880),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_855),
.A2(n_681),
.B(n_734),
.C(n_654),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_884),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_891),
.B(n_662),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_793),
.A2(n_747),
.B(n_740),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_810),
.B(n_662),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_853),
.B(n_666),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_810),
.B(n_689),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_788),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_773),
.A2(n_460),
.B(n_666),
.Y(n_972)
);

AOI221xp5_ASAP7_75t_L g973 ( 
.A1(n_947),
.A2(n_460),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_776),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_829),
.B(n_666),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_884),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_809),
.A2(n_460),
.B(n_666),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_907),
.A2(n_4),
.B(n_9),
.C(n_13),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_789),
.B(n_844),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_947),
.A2(n_460),
.B(n_13),
.C(n_15),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_867),
.B(n_9),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_811),
.A2(n_75),
.B(n_144),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_915),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_899),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_L g985 ( 
.A(n_783),
.B(n_79),
.Y(n_985)
);

AO32x2_ASAP7_75t_L g986 ( 
.A1(n_883),
.A2(n_19),
.A3(n_23),
.B1(n_27),
.B2(n_30),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_789),
.B(n_27),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_821),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_L g989 ( 
.A1(n_792),
.A2(n_86),
.B(n_138),
.C(n_135),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_923),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.C(n_43),
.Y(n_990)
);

CKINVDCx8_ASAP7_75t_R g991 ( 
.A(n_846),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_948),
.B(n_36),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_861),
.A2(n_877),
.B(n_952),
.C(n_814),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_783),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_786),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_SL g997 ( 
.A1(n_952),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_871),
.B(n_49),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_804),
.A2(n_108),
.B(n_134),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_843),
.A2(n_103),
.B(n_133),
.C(n_131),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_884),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_871),
.B(n_50),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_SL g1003 ( 
.A1(n_858),
.A2(n_51),
.B(n_55),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_861),
.A2(n_877),
.B(n_819),
.C(n_872),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_796),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_783),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_825),
.A2(n_99),
.B(n_126),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_950),
.Y(n_1008)
);

AOI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_801),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.C(n_74),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_922),
.A2(n_111),
.B(n_112),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_912),
.B(n_117),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_815),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_813),
.A2(n_145),
.B(n_823),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_805),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_815),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_921),
.B(n_774),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_791),
.B(n_808),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_843),
.A2(n_806),
.B(n_945),
.C(n_900),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_823),
.A2(n_820),
.B(n_930),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_783),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_775),
.B(n_887),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_824),
.B(n_932),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_785),
.B(n_787),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_884),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_950),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_932),
.B(n_890),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_951),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_812),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_866),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_797),
.B(n_933),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_934),
.A2(n_827),
.B(n_840),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_812),
.B(n_901),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_812),
.B(n_858),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_795),
.A2(n_836),
.B(n_840),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_839),
.A2(n_812),
.B1(n_863),
.B2(n_856),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_822),
.B(n_831),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_794),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_795),
.A2(n_827),
.B(n_836),
.Y(n_1038)
);

AOI22x1_ASAP7_75t_L g1039 ( 
.A1(n_931),
.A2(n_864),
.B1(n_926),
.B2(n_848),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_909),
.B(n_799),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_798),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_SL g1042 ( 
.A1(n_944),
.A2(n_945),
.B(n_832),
.C(n_835),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_794),
.B(n_879),
.Y(n_1043)
);

OAI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_817),
.A2(n_868),
.B1(n_916),
.B2(n_906),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_879),
.B(n_838),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_850),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_916),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_903),
.A2(n_800),
.B1(n_807),
.B2(n_803),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_799),
.B(n_929),
.Y(n_1049)
);

OA21x2_ASAP7_75t_L g1050 ( 
.A1(n_816),
.A2(n_941),
.B(n_902),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_852),
.A2(n_841),
.B(n_870),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_860),
.B(n_780),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_SL g1053 ( 
.A(n_777),
.B(n_842),
.C(n_935),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_781),
.B(n_782),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_802),
.B(n_790),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_834),
.A2(n_849),
.B(n_896),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_849),
.A2(n_874),
.B(n_826),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_938),
.A2(n_830),
.B(n_881),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_869),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_953),
.B(n_888),
.C(n_885),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_857),
.A2(n_893),
.B(n_918),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_833),
.A2(n_919),
.B(n_949),
.C(n_946),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_889),
.A2(n_886),
.B1(n_859),
.B2(n_939),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_895),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_875),
.A2(n_876),
.B(n_924),
.C(n_936),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_857),
.A2(n_940),
.B(n_865),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_897),
.B(n_908),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_SL g1068 ( 
.A(n_882),
.B(n_956),
.C(n_954),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_886),
.B(n_859),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_955),
.B(n_937),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_862),
.B(n_865),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_862),
.B(n_911),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_873),
.A2(n_892),
.B1(n_894),
.B2(n_910),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_878),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_942),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_928),
.A2(n_914),
.B(n_913),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_828),
.B(n_898),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_828),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_854),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_905),
.A2(n_920),
.B(n_925),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_943),
.A2(n_855),
.B(n_847),
.C(n_947),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_927),
.A2(n_847),
.B1(n_855),
.B2(n_947),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_847),
.A2(n_612),
.B1(n_855),
.B2(n_488),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_784),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_845),
.B(n_810),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_797),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_884),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_855),
.B(n_801),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_776),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_847),
.A2(n_855),
.B1(n_891),
.B2(n_616),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_779),
.A2(n_818),
.B(n_614),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_851),
.B(n_853),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_851),
.B(n_853),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_784),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_884),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_SL g1096 ( 
.A(n_789),
.B(n_584),
.C(n_722),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_899),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_851),
.B(n_853),
.Y(n_1098)
);

INVx8_ASAP7_75t_L g1099 ( 
.A(n_783),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_776),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_855),
.A2(n_847),
.B(n_907),
.C(n_915),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1056),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_958),
.A2(n_1091),
.B(n_1019),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1054),
.A2(n_1035),
.B(n_1061),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_991),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1081),
.A2(n_1004),
.B(n_1021),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1051),
.A2(n_1057),
.B(n_967),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_1101),
.A2(n_987),
.B1(n_1083),
.B2(n_973),
.C(n_1090),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_963),
.A2(n_972),
.B(n_1058),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1084),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_957),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1099),
.B(n_1020),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1077),
.A2(n_1078),
.A3(n_1073),
.B(n_1066),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_SL g1116 ( 
.A1(n_1075),
.A2(n_1072),
.B(n_998),
.C(n_1002),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1039),
.A2(n_977),
.B(n_1013),
.Y(n_1117)
);

AO32x2_ASAP7_75t_L g1118 ( 
.A1(n_1048),
.A2(n_1083),
.A3(n_1073),
.B1(n_1063),
.B2(n_986),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1088),
.A2(n_1030),
.B1(n_1098),
.B2(n_1036),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_988),
.B(n_992),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_1094),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1089),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_971),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_984),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1050),
.A2(n_1065),
.B(n_1031),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1034),
.A2(n_1038),
.B(n_1042),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_988),
.B(n_968),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1082),
.A2(n_993),
.B(n_964),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_1088),
.B(n_1086),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1040),
.A2(n_968),
.B1(n_962),
.B2(n_979),
.Y(n_1130)
);

AOI221x1_ASAP7_75t_L g1131 ( 
.A1(n_961),
.A2(n_980),
.B1(n_1048),
.B2(n_1053),
.C(n_1060),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1082),
.A2(n_978),
.B(n_1044),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1009),
.B(n_990),
.C(n_1096),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_1046),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1070),
.A2(n_1074),
.B(n_989),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1063),
.A2(n_999),
.A3(n_1007),
.B(n_982),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_969),
.A2(n_1011),
.A3(n_1014),
.B(n_1041),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_960),
.A2(n_1052),
.B1(n_1023),
.B2(n_966),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1032),
.A2(n_1068),
.B(n_1010),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1047),
.A2(n_1100),
.B1(n_1033),
.B2(n_975),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1055),
.A2(n_1045),
.B(n_1071),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_983),
.B(n_981),
.C(n_1003),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1049),
.B(n_1064),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_996),
.A2(n_1015),
.A3(n_1012),
.B(n_1005),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_986),
.A2(n_997),
.A3(n_1003),
.B1(n_1006),
.B2(n_994),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1067),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1016),
.A2(n_1026),
.B(n_1086),
.C(n_1062),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_1099),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1085),
.B(n_959),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1027),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1059),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1017),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_1028),
.B(n_1087),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1022),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1018),
.A2(n_985),
.B(n_1024),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1043),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_959),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1037),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1069),
.A2(n_1000),
.B(n_1024),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1020),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_965),
.Y(n_1162)
);

CKINVDCx6p67_ASAP7_75t_R g1163 ( 
.A(n_1025),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_994),
.A2(n_1006),
.A3(n_986),
.B(n_1069),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1024),
.B(n_1047),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1079),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_970),
.B(n_995),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1099),
.A2(n_976),
.B(n_1001),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_970),
.B(n_1037),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1037),
.B(n_1028),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1097),
.B(n_976),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_976),
.A2(n_1001),
.B(n_1087),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1001),
.A2(n_1087),
.B(n_1095),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1095),
.B(n_1029),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1008),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1095),
.B(n_891),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1101),
.A2(n_855),
.B(n_847),
.C(n_961),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1092),
.A2(n_1093),
.B1(n_1098),
.B2(n_847),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1085),
.B(n_962),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1101),
.A2(n_855),
.B(n_847),
.C(n_961),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1046),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_958),
.A2(n_1091),
.B(n_779),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_964),
.A2(n_855),
.B(n_961),
.C(n_847),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_958),
.A2(n_1091),
.B(n_779),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_958),
.A2(n_1091),
.B(n_779),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_964),
.A2(n_855),
.B(n_468),
.C(n_847),
.Y(n_1186)
);

OAI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1088),
.A2(n_471),
.B1(n_468),
.B2(n_661),
.C(n_659),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_974),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_1088),
.B(n_801),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1017),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_974),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1058),
.A2(n_1066),
.B(n_1061),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1088),
.A2(n_947),
.B1(n_847),
.B2(n_1083),
.Y(n_1193)
);

AO21x1_ASAP7_75t_L g1194 ( 
.A1(n_1101),
.A2(n_1088),
.B(n_847),
.Y(n_1194)
);

AOI31xp67_ASAP7_75t_L g1195 ( 
.A1(n_1082),
.A2(n_1078),
.A3(n_1077),
.B(n_1072),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_SL g1196 ( 
.A(n_1088),
.B(n_468),
.C(n_801),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_988),
.B(n_668),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1099),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1061),
.A2(n_1077),
.A3(n_1078),
.B(n_1081),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_964),
.A2(n_855),
.B(n_961),
.C(n_847),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1061),
.A2(n_1077),
.A3(n_1078),
.B(n_1081),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1092),
.B(n_801),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1017),
.Y(n_1205)
);

BUFx4f_ASAP7_75t_L g1206 ( 
.A(n_1046),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_987),
.A2(n_947),
.B1(n_909),
.B2(n_966),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1088),
.A2(n_947),
.B1(n_847),
.B2(n_1083),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_958),
.A2(n_1091),
.B(n_779),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1101),
.A2(n_855),
.B(n_1042),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1101),
.A2(n_855),
.B(n_1042),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1088),
.A2(n_947),
.B1(n_847),
.B2(n_1083),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1017),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1099),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_987),
.A2(n_947),
.B1(n_909),
.B2(n_966),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1080),
.A2(n_778),
.B(n_1076),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1061),
.A2(n_1077),
.A3(n_1078),
.B(n_1081),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_957),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_957),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1061),
.A2(n_1077),
.A3(n_1078),
.B(n_1081),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_963),
.A2(n_1077),
.B(n_1061),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1101),
.A2(n_471),
.B1(n_450),
.B2(n_596),
.C(n_947),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1101),
.A2(n_855),
.B(n_1042),
.Y(n_1224)
);

NOR3xp33_ASAP7_75t_L g1225 ( 
.A(n_1030),
.B(n_722),
.C(n_468),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1088),
.A2(n_947),
.B1(n_847),
.B2(n_1083),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1061),
.A2(n_1077),
.A3(n_1078),
.B(n_1081),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_L g1228 ( 
.A1(n_1081),
.A2(n_847),
.B(n_855),
.C(n_998),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1092),
.B(n_801),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1101),
.A2(n_855),
.B(n_1042),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_987),
.A2(n_947),
.B1(n_909),
.B2(n_966),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_SL g1232 ( 
.A(n_991),
.B(n_688),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1085),
.B(n_962),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1092),
.A2(n_1093),
.B1(n_1098),
.B2(n_847),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_991),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_988),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1084),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_958),
.A2(n_1091),
.B(n_779),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1080),
.A2(n_778),
.B(n_1076),
.Y(n_1239)
);

INVx6_ASAP7_75t_L g1240 ( 
.A(n_1148),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1198),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1187),
.A2(n_1208),
.B1(n_1226),
.B2(n_1212),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1107),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1189),
.A2(n_1129),
.B1(n_1208),
.B2(n_1212),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1189),
.A2(n_1129),
.B1(n_1128),
.B2(n_1133),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1122),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1165),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_1105),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1235),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1223),
.A2(n_1196),
.B1(n_1110),
.B2(n_1225),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1188),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1191),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1148),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1182),
.A2(n_1185),
.B(n_1184),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1133),
.A2(n_1193),
.B1(n_1226),
.B2(n_1128),
.Y(n_1255)
);

INVx6_ASAP7_75t_L g1256 ( 
.A(n_1148),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1166),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1193),
.A2(n_1119),
.B1(n_1130),
.B2(n_1147),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1134),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1164),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1218),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1194),
.A2(n_1215),
.B1(n_1207),
.B2(n_1231),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1124),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1121),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1143),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1167),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1153),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1167),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1144),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1204),
.A2(n_1229),
.B1(n_1132),
.B2(n_1142),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1142),
.A2(n_1234),
.B1(n_1178),
.B2(n_1224),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1112),
.Y(n_1273)
);

BUFx8_ASAP7_75t_L g1274 ( 
.A(n_1181),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1123),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1123),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1158),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1236),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1109),
.A2(n_1197),
.B1(n_1219),
.B2(n_1201),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1190),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1177),
.A2(n_1180),
.B1(n_1186),
.B2(n_1120),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1210),
.A2(n_1230),
.B1(n_1224),
.B2(n_1211),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1210),
.A2(n_1230),
.B1(n_1211),
.B2(n_1106),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1171),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1214),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1163),
.Y(n_1286)
);

BUFx8_ASAP7_75t_L g1287 ( 
.A(n_1149),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1138),
.A2(n_1146),
.B1(n_1155),
.B2(n_1127),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1176),
.A2(n_1113),
.B1(n_1161),
.B2(n_1152),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1237),
.B(n_1179),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1104),
.A2(n_1151),
.B1(n_1140),
.B2(n_1156),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1205),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1179),
.A2(n_1233),
.B1(n_1183),
.B2(n_1202),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1233),
.A2(n_1161),
.B1(n_1135),
.B2(n_1157),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1214),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1213),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1114),
.B(n_1169),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1131),
.A2(n_1114),
.B1(n_1175),
.B2(n_1174),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1206),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1137),
.B(n_1159),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1162),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1228),
.A2(n_1116),
.B(n_1141),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1170),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1173),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1135),
.A2(n_1125),
.B1(n_1114),
.B2(n_1222),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_1206),
.B1(n_1172),
.B2(n_1238),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1150),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1150),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1137),
.B(n_1217),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1222),
.A2(n_1232),
.B1(n_1126),
.B2(n_1117),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1137),
.B(n_1203),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1150),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1103),
.A2(n_1209),
.B1(n_1139),
.B2(n_1118),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1118),
.A2(n_1160),
.B1(n_1199),
.B2(n_1154),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1154),
.A2(n_1168),
.B1(n_1108),
.B2(n_1216),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1154),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1118),
.A2(n_1111),
.B1(n_1239),
.B2(n_1102),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1145),
.A2(n_1203),
.B1(n_1221),
.B2(n_1217),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1145),
.A2(n_1203),
.B1(n_1221),
.B2(n_1217),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_1200),
.B1(n_1221),
.B2(n_1227),
.Y(n_1321)
);

CKINVDCx8_ASAP7_75t_R g1322 ( 
.A(n_1227),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1115),
.A2(n_1187),
.B1(n_1223),
.B2(n_1088),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1192),
.A2(n_1136),
.B1(n_1187),
.B2(n_1093),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1136),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1136),
.A2(n_1187),
.B1(n_1093),
.B2(n_1098),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1189),
.A2(n_1088),
.B1(n_1187),
.B2(n_801),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1107),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1187),
.A2(n_1189),
.B1(n_1088),
.B2(n_1129),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1187),
.A2(n_1223),
.B1(n_1088),
.B2(n_1196),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1189),
.A2(n_1088),
.B1(n_1187),
.B2(n_801),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1189),
.A2(n_1088),
.B1(n_1187),
.B2(n_801),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1121),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1124),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1165),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1189),
.A2(n_1187),
.B1(n_1088),
.B2(n_1196),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1187),
.A2(n_1223),
.B1(n_1088),
.B2(n_1196),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1107),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1235),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1198),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1189),
.A2(n_1187),
.B1(n_1088),
.B2(n_1129),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1235),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1124),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1235),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_1105),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1189),
.A2(n_1088),
.B1(n_1187),
.B2(n_801),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1134),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1187),
.A2(n_1189),
.B1(n_1196),
.B2(n_1088),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1189),
.A2(n_1088),
.B1(n_1187),
.B2(n_801),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1120),
.B(n_1149),
.Y(n_1351)
);

BUFx8_ASAP7_75t_L g1352 ( 
.A(n_1134),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1124),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1322),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1240),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1269),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1254),
.A2(n_1302),
.B(n_1305),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1325),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1305),
.A2(n_1310),
.B(n_1318),
.Y(n_1359)
);

AOI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1324),
.A2(n_1317),
.B(n_1326),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1325),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1300),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1260),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1283),
.B(n_1255),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1278),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1304),
.B(n_1315),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1316),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1327),
.A2(n_1350),
.B1(n_1331),
.B2(n_1332),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1309),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1242),
.A2(n_1329),
.B1(n_1258),
.B2(n_1281),
.Y(n_1370)
);

NOR2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1336),
.B(n_1247),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1316),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1283),
.B(n_1255),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1284),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1311),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1243),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1246),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1284),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1342),
.A2(n_1250),
.B(n_1244),
.C(n_1330),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1251),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1310),
.A2(n_1318),
.B(n_1313),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1313),
.A2(n_1282),
.B(n_1321),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1273),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1252),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1291),
.A2(n_1306),
.B(n_1319),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1297),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1249),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1328),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1282),
.B(n_1272),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1250),
.A2(n_1338),
.B(n_1330),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1240),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1241),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1343),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1291),
.A2(n_1319),
.B(n_1320),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1342),
.A2(n_1323),
.B(n_1350),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1323),
.B(n_1245),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1339),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1245),
.B(n_1262),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1297),
.B(n_1293),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1338),
.B(n_1320),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1253),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1253),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1321),
.B(n_1244),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1271),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1253),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1303),
.B(n_1337),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1270),
.B(n_1349),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1327),
.B(n_1331),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1332),
.B(n_1347),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1341),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1351),
.B(n_1296),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1261),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1347),
.B(n_1265),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1248),
.B(n_1346),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1294),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1275),
.B(n_1298),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1294),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1301),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1314),
.B(n_1288),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1256),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1279),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1285),
.B(n_1295),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1298),
.A2(n_1308),
.B1(n_1312),
.B2(n_1289),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1266),
.A2(n_1268),
.B(n_1290),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1287),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1247),
.B(n_1335),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1277),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1333),
.Y(n_1430)
);

NAND2x1_ASAP7_75t_L g1431 ( 
.A(n_1285),
.B(n_1295),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1423),
.B(n_1264),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1391),
.A2(n_1299),
.B(n_1280),
.C(n_1263),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_SL g1434 ( 
.A(n_1380),
.B(n_1267),
.C(n_1276),
.D(n_1286),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1361),
.B(n_1353),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1377),
.B(n_1307),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1356),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1386),
.B(n_1295),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1362),
.B(n_1344),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1365),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1357),
.A2(n_1285),
.B(n_1257),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1380),
.A2(n_1334),
.B(n_1287),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1366),
.Y(n_1443)
);

A2O1A1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1391),
.A2(n_1340),
.B(n_1259),
.C(n_1280),
.Y(n_1444)
);

INVx5_ASAP7_75t_L g1445 ( 
.A(n_1354),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1446)
);

INVxp33_ASAP7_75t_SL g1447 ( 
.A(n_1416),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1370),
.A2(n_1292),
.B(n_1274),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1375),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1362),
.B(n_1274),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1378),
.B(n_1345),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1368),
.B(n_1348),
.C(n_1352),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1396),
.A2(n_1418),
.B(n_1409),
.C(n_1411),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1396),
.A2(n_1425),
.B1(n_1411),
.B2(n_1409),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1384),
.Y(n_1458)
);

NAND4xp25_ASAP7_75t_L g1459 ( 
.A(n_1423),
.B(n_1407),
.C(n_1415),
.D(n_1418),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1405),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1425),
.A2(n_1399),
.B(n_1390),
.C(n_1408),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1413),
.B(n_1393),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_L g1463 ( 
.A(n_1397),
.B(n_1371),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1357),
.A2(n_1382),
.B(n_1359),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1397),
.A2(n_1399),
.B(n_1373),
.C(n_1364),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_SL g1466 ( 
.A(n_1369),
.B(n_1376),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1363),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1360),
.A2(n_1359),
.B(n_1382),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1390),
.A2(n_1408),
.B1(n_1364),
.B2(n_1373),
.C(n_1421),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1415),
.A2(n_1407),
.B1(n_1400),
.B2(n_1421),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1398),
.B(n_1389),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1426),
.A2(n_1386),
.B(n_1431),
.Y(n_1473)
);

AO32x2_ASAP7_75t_L g1474 ( 
.A1(n_1355),
.A2(n_1392),
.A3(n_1403),
.B1(n_1406),
.B2(n_1383),
.Y(n_1474)
);

AOI211xp5_ASAP7_75t_L g1475 ( 
.A1(n_1426),
.A2(n_1414),
.B(n_1428),
.C(n_1419),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1354),
.A2(n_1404),
.B(n_1395),
.C(n_1371),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_R g1477 ( 
.A(n_1388),
.B(n_1394),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_SL g1478 ( 
.A(n_1374),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1424),
.A2(n_1431),
.B(n_1354),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1420),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1405),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1361),
.B(n_1387),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1472),
.B(n_1369),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1437),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1474),
.B(n_1383),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1474),
.B(n_1366),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1474),
.B(n_1383),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1474),
.B(n_1383),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1467),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1455),
.B(n_1419),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1454),
.A2(n_1452),
.B1(n_1448),
.B2(n_1457),
.C(n_1461),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1366),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1468),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1482),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1466),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1443),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1395),
.Y(n_1500)
);

OR2x2_ASAP7_75t_SL g1501 ( 
.A(n_1441),
.B(n_1404),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1455),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1473),
.B(n_1354),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1438),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1438),
.B(n_1361),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1480),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1491),
.B(n_1449),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1484),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1494),
.A2(n_1434),
.B1(n_1469),
.B2(n_1459),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1506),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1501),
.B(n_1460),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1501),
.B(n_1458),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1501),
.B(n_1480),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1499),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_SL g1518 ( 
.A(n_1494),
.B(n_1433),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1504),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1503),
.A2(n_1444),
.B1(n_1465),
.B2(n_1442),
.C(n_1475),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1499),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1484),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1506),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1486),
.A2(n_1470),
.B1(n_1440),
.B2(n_1463),
.C(n_1471),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1503),
.A2(n_1447),
.B1(n_1358),
.B2(n_1478),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1492),
.B(n_1456),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1493),
.B(n_1483),
.Y(n_1528)
);

AOI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1496),
.A2(n_1479),
.B(n_1358),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

AOI211xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1498),
.A2(n_1463),
.B(n_1476),
.C(n_1450),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1504),
.A2(n_1445),
.B1(n_1450),
.B2(n_1432),
.Y(n_1532)
);

OAI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1503),
.A2(n_1462),
.B(n_1481),
.C(n_1439),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1487),
.B(n_1466),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1486),
.A2(n_1401),
.B1(n_1447),
.B2(n_1451),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1485),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1510),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1477),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1534),
.B(n_1487),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1513),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1534),
.B(n_1487),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1502),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1522),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1528),
.B(n_1493),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1522),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1519),
.B(n_1505),
.Y(n_1553)
);

NAND2x1_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1505),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1497),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1511),
.B(n_1374),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1451),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1513),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1509),
.B(n_1490),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1523),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1536),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1509),
.B(n_1490),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1536),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

NOR4xp25_ASAP7_75t_SL g1565 ( 
.A(n_1520),
.B(n_1498),
.C(n_1430),
.D(n_1429),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1549),
.B(n_1533),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1544),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1543),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1559),
.B(n_1515),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1549),
.A2(n_1511),
.B(n_1524),
.C(n_1531),
.Y(n_1573)
);

NOR2x1p5_ASAP7_75t_SL g1574 ( 
.A(n_1537),
.B(n_1529),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1557),
.B(n_1533),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1551),
.B(n_1535),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1544),
.B(n_1525),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1551),
.B(n_1535),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1507),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1559),
.B(n_1515),
.Y(n_1580)
);

NAND4xp75_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1524),
.C(n_1556),
.D(n_1505),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1508),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1562),
.B(n_1514),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1514),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1538),
.B(n_1545),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1374),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1537),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1545),
.B(n_1514),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1546),
.B(n_1531),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1553),
.A2(n_1516),
.B(n_1489),
.Y(n_1595)
);

AND2x2_ASAP7_75t_SL g1596 ( 
.A(n_1565),
.B(n_1453),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1547),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1547),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1564),
.B(n_1527),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1548),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1548),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1564),
.B(n_1527),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1553),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1564),
.B(n_1508),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1553),
.A2(n_1516),
.B(n_1489),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1587),
.B(n_1541),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1567),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1600),
.B(n_1541),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1597),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1597),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1553),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.B(n_1564),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1550),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1599),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1605),
.B(n_1558),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1599),
.Y(n_1620)
);

OAI321xp33_ASAP7_75t_L g1621 ( 
.A1(n_1573),
.A2(n_1525),
.A3(n_1532),
.B1(n_1529),
.B2(n_1565),
.C(n_1500),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_1560),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1596),
.B(n_1532),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1607),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1594),
.B(n_1560),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1607),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1577),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1576),
.B(n_1578),
.C(n_1589),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1552),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1379),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1606),
.B(n_1550),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1568),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1588),
.Y(n_1635)
);

CKINVDCx16_ASAP7_75t_R g1636 ( 
.A(n_1584),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1512),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1596),
.B(n_1512),
.Y(n_1638)
);

NAND2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1570),
.B(n_1554),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1571),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1595),
.B(n_1512),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1512),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1604),
.B(n_1550),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1617),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1630),
.A2(n_1519),
.B1(n_1530),
.B2(n_1504),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1621),
.A2(n_1604),
.B(n_1582),
.C(n_1580),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1617),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1623),
.A2(n_1604),
.B(n_1586),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1569),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1627),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1637),
.A2(n_1529),
.B(n_1570),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1639),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1622),
.A2(n_1580),
.B(n_1591),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1593),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1620),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1620),
.Y(n_1658)
);

OAI322xp33_ASAP7_75t_L g1659 ( 
.A1(n_1618),
.A2(n_1591),
.A3(n_1593),
.B1(n_1598),
.B2(n_1571),
.C1(n_1590),
.C2(n_1603),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1614),
.B(n_1569),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1625),
.A2(n_1603),
.B1(n_1598),
.B2(n_1590),
.C(n_1500),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1638),
.A2(n_1530),
.B1(n_1379),
.B2(n_1521),
.C(n_1517),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1636),
.A2(n_1615),
.B1(n_1644),
.B2(n_1631),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1634),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1639),
.B(n_1430),
.C(n_1453),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1612),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1609),
.A2(n_1530),
.B(n_1500),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1645),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1651),
.A2(n_1609),
.B1(n_1643),
.B2(n_1642),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1660),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1611),
.B1(n_1619),
.B2(n_1635),
.C(n_1626),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1651),
.B(n_1644),
.C(n_1640),
.D(n_1611),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1662),
.B(n_1631),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1662),
.B(n_1640),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1649),
.A2(n_1619),
.B(n_1613),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1655),
.B(n_1624),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1656),
.B(n_1624),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1648),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1654),
.B(n_1626),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1657),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1633),
.C(n_1632),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1661),
.B(n_1572),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1658),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1669),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_SL g1688 ( 
.A(n_1647),
.B(n_1629),
.C(n_1592),
.D(n_1585),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1629),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1663),
.A2(n_1641),
.B1(n_1530),
.B2(n_1436),
.C(n_1585),
.Y(n_1690)
);

OAI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1646),
.A2(n_1574),
.B(n_1641),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

INVxp33_ASAP7_75t_L g1693 ( 
.A(n_1675),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1673),
.B(n_1660),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1689),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1650),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1682),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1680),
.B(n_1653),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1684),
.B(n_1653),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1677),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1685),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1674),
.A2(n_1664),
.B1(n_1652),
.B2(n_1667),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1701),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1698),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1697),
.B(n_1687),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1693),
.B(n_1678),
.C(n_1694),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1695),
.B(n_1679),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1702),
.A2(n_1688),
.B(n_1678),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1696),
.B(n_1667),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1700),
.B(n_1671),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_SL g1711 ( 
.A1(n_1700),
.A2(n_1379),
.B1(n_1683),
.B2(n_1681),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1708),
.A2(n_1699),
.B(n_1672),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1706),
.A2(n_1691),
.B(n_1668),
.C(n_1690),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1705),
.A2(n_1672),
.B1(n_1659),
.B2(n_1692),
.C(n_1686),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1707),
.A2(n_1670),
.B(n_1668),
.C(n_1439),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1703),
.B(n_1572),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1713),
.A2(n_1709),
.B1(n_1704),
.B2(n_1710),
.C(n_1711),
.Y(n_1717)
);

O2A1O1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1712),
.A2(n_1427),
.B(n_1372),
.C(n_1367),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1716),
.B(n_1427),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1592),
.Y(n_1720)
);

NAND4xp25_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1427),
.C(n_1372),
.D(n_1367),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1716),
.Y(n_1722)
);

NOR2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1720),
.B(n_1367),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1722),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1719),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1718),
.B(n_1574),
.Y(n_1726)
);

NAND4xp75_ASAP7_75t_L g1727 ( 
.A(n_1717),
.B(n_1583),
.C(n_1579),
.D(n_1436),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1725),
.B(n_1372),
.Y(n_1728)
);

NAND4xp75_ASAP7_75t_L g1729 ( 
.A(n_1724),
.B(n_1721),
.C(n_1583),
.D(n_1579),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1727),
.A2(n_1723),
.B1(n_1726),
.B2(n_1435),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1729),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1731),
.Y(n_1732)
);

O2A1O1Ixp33_ASAP7_75t_SL g1733 ( 
.A1(n_1732),
.A2(n_1730),
.B(n_1728),
.C(n_1424),
.Y(n_1733)
);

XNOR2xp5_ASAP7_75t_L g1734 ( 
.A(n_1732),
.B(n_1435),
.Y(n_1734)
);

OAI22x1_ASAP7_75t_L g1735 ( 
.A1(n_1734),
.A2(n_1435),
.B1(n_1429),
.B2(n_1521),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1733),
.B(n_1523),
.C(n_1552),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1736),
.A2(n_1517),
.B1(n_1521),
.B2(n_1563),
.Y(n_1737)
);

AO21x2_ASAP7_75t_L g1738 ( 
.A1(n_1735),
.A2(n_1561),
.B(n_1563),
.Y(n_1738)
);

XNOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1737),
.B(n_1402),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1738),
.B(n_1428),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1740),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1392),
.B1(n_1355),
.B2(n_1402),
.C(n_1410),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1422),
.B(n_1410),
.C(n_1402),
.Y(n_1743)
);


endmodule