module fake_jpeg_24093_n_268 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_35),
.B1(n_17),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_52),
.B1(n_66),
.B2(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_20),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_17),
.B1(n_29),
.B2(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_59),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_16),
.B1(n_25),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_22),
.B1(n_32),
.B2(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_33),
.A2(n_30),
.B1(n_31),
.B2(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_81),
.B1(n_49),
.B2(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_88),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_20),
.B1(n_28),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_47),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_20),
.C(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_62),
.C(n_64),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_21),
.B1(n_26),
.B2(n_6),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_24),
.B1(n_23),
.B2(n_27),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_96),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_59),
.C(n_55),
.Y(n_129)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_63),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_109),
.C(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_58),
.B1(n_53),
.B2(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_86),
.B1(n_72),
.B2(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_76),
.Y(n_114)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_85),
.B1(n_88),
.B2(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_49),
.B1(n_70),
.B2(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_48),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_116),
.Y(n_138)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_123),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_97),
.B1(n_108),
.B2(n_51),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_129),
.C(n_97),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_125),
.B1(n_108),
.B2(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_92),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_82),
.B(n_50),
.C(n_23),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_96),
.Y(n_135)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_104),
.B1(n_75),
.B2(n_88),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_154),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_148),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_122),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_8),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_101),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_156),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_147),
.B1(n_160),
.B2(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_110),
.B(n_99),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_153),
.B(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_98),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_161),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_102),
.B1(n_100),
.B2(n_48),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_159),
.B1(n_154),
.B2(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_83),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_51),
.B1(n_50),
.B2(n_68),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_79),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_50),
.B(n_1),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_166),
.B1(n_171),
.B2(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_118),
.B1(n_125),
.B2(n_116),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_135),
.B1(n_126),
.B2(n_116),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_155),
.B1(n_152),
.B2(n_3),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_129),
.B1(n_126),
.B2(n_130),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_130),
.B(n_135),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_175),
.B(n_177),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_123),
.B1(n_115),
.B2(n_23),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_142),
.B1(n_149),
.B2(n_156),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_79),
.B(n_68),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_68),
.B(n_1),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_145),
.B(n_148),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_152),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_184),
.B(n_150),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

XOR2x2_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_141),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_193),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_9),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_200),
.B(n_202),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_201),
.B1(n_204),
.B2(n_168),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_158),
.C(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_183),
.C(n_171),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_181),
.B1(n_184),
.B2(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_145),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_185),
.B1(n_168),
.B2(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_208),
.C(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_180),
.C(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_191),
.B1(n_205),
.B2(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_170),
.B1(n_178),
.B2(n_3),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_216),
.B1(n_220),
.B2(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_178),
.C(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_193),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_203),
.B1(n_186),
.B2(n_191),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_0),
.C(n_2),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.C(n_200),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_230),
.C(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_201),
.C(n_202),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_233),
.C(n_234),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_232),
.B1(n_217),
.B2(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_188),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_218),
.B1(n_212),
.B2(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_237),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_219),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_212),
.C(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_188),
.C(n_10),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_234),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_231),
.B(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_12),
.C(n_14),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_232),
.B(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_251),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_225),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_10),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_15),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_14),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_251),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_12),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_256),
.A2(n_257),
.B1(n_15),
.B2(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_14),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_262),
.B(n_5),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_245),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_262),
.C(n_260),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_5),
.Y(n_268)
);


endmodule