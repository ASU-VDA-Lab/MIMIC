module fake_jpeg_6335_n_336 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_3),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_37),
.B(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_12),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_51),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_11),
.Y(n_103)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_59),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_62),
.Y(n_116)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_27),
.B(n_32),
.C(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_79),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_75),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_72),
.B(n_78),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_86),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_34),
.B1(n_33),
.B2(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_16),
.B1(n_31),
.B2(n_17),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_37),
.B(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_16),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_23),
.B1(n_14),
.B2(n_34),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_33),
.B1(n_22),
.B2(n_10),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_56),
.B1(n_52),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_23),
.Y(n_99)
);

CKINVDCx9p33_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_105),
.B(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_43),
.B(n_10),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_33),
.B1(n_22),
.B2(n_10),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_109),
.A2(n_118),
.B1(n_128),
.B2(n_130),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_102),
.B1(n_61),
.B2(n_104),
.Y(n_157)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_114),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_59),
.B1(n_74),
.B2(n_96),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_131),
.B1(n_133),
.B2(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_58),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_84),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_62),
.A2(n_0),
.B1(n_7),
.B2(n_8),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_7),
.B1(n_8),
.B2(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_143),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_73),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_151),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_78),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_65),
.B1(n_83),
.B2(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_112),
.B1(n_108),
.B2(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_71),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_60),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_160),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_72),
.B(n_61),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_163),
.B(n_168),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_162),
.B1(n_164),
.B2(n_143),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_159),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_80),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_80),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_81),
.C(n_77),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_108),
.C(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_110),
.A2(n_101),
.B(n_100),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_82),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_77),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_136),
.Y(n_180)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_175),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_112),
.A2(n_91),
.B1(n_97),
.B2(n_92),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_124),
.B1(n_138),
.B2(n_119),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_8),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_131),
.B(n_128),
.C(n_112),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_204),
.B(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_182),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_132),
.B1(n_114),
.B2(n_111),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_186),
.B1(n_196),
.B2(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_208),
.B1(n_178),
.B2(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_122),
.B1(n_129),
.B2(n_139),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_212),
.B1(n_187),
.B2(n_196),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_67),
.C(n_122),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_207),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_139),
.B1(n_79),
.B2(n_124),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_201),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_67),
.B(n_124),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_206),
.B(n_152),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_124),
.B1(n_138),
.B2(n_67),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_141),
.B(n_8),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_155),
.A2(n_86),
.B(n_121),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_86),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_142),
.A2(n_86),
.B1(n_121),
.B2(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_150),
.B(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_142),
.A2(n_145),
.B1(n_159),
.B2(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_144),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_231),
.B1(n_234),
.B2(n_241),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_221),
.A2(n_181),
.B1(n_194),
.B2(n_182),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_151),
.B(n_148),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_151),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_229),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_163),
.B(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_161),
.B(n_175),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_164),
.B(n_167),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_140),
.B(n_153),
.Y(n_241)
);

AOI32xp33_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_153),
.A3(n_173),
.B1(n_158),
.B2(n_156),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_243),
.B(n_200),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_SL g243 ( 
.A(n_180),
.B(n_153),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_195),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_254),
.Y(n_275)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_204),
.B(n_179),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_207),
.B(n_208),
.C(n_186),
.D(n_205),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_191),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_263),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_190),
.C(n_185),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_219),
.C(n_241),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_184),
.B1(n_209),
.B2(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_232),
.B1(n_240),
.B2(n_221),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_218),
.B(n_177),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_188),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_179),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_266),
.B1(n_267),
.B2(n_251),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_225),
.B(n_229),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_257),
.C(n_252),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_216),
.B1(n_228),
.B2(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_216),
.B1(n_235),
.B2(n_226),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_219),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_280),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_226),
.B1(n_218),
.B2(n_236),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_265),
.B1(n_253),
.B2(n_254),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_237),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_247),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_245),
.B(n_177),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_233),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.C(n_260),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_202),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_258),
.B(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_250),
.B(n_246),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_279),
.B(n_275),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_250),
.B(n_267),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_289),
.A2(n_291),
.B(n_274),
.C(n_272),
.Y(n_311)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_294),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_273),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_298),
.B(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_270),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_257),
.C(n_280),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_278),
.A2(n_265),
.B(n_244),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_302),
.B(n_308),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_268),
.B1(n_285),
.B2(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_284),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_217),
.B1(n_255),
.B2(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_255),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_259),
.B(n_244),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_291),
.B1(n_293),
.B2(n_289),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_259),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_317),
.B(n_263),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_304),
.B1(n_296),
.B2(n_302),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_245),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_282),
.C(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_262),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_288),
.B(n_292),
.C(n_311),
.D(n_289),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_318),
.B1(n_315),
.B2(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_319),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.A3(n_329),
.B1(n_323),
.B2(n_314),
.C1(n_330),
.C2(n_262),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_314),
.C(n_330),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_262),
.B(n_183),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_211),
.Y(n_336)
);


endmodule