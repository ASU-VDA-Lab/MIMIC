module real_jpeg_2148_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_2),
.B(n_19),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_2),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_6),
.B(n_93),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_8),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_40),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_75),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_52),
.B(n_74),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_31),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.C(n_29),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_17),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_17),
.A2(n_18),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_20),
.Y(n_17)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_28),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_41),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_42),
.C(n_46),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_34),
.B(n_37),
.C(n_38),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_48),
.B(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_65),
.B(n_73),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_64),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_100),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_103),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_90),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);


endmodule