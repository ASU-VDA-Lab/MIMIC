module real_jpeg_20968_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_53),
.B1(n_59),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_0),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_97),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_0),
.A2(n_29),
.B1(n_31),
.B2(n_97),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_97),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_55),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_16),
.B(n_29),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_108),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_27),
.B1(n_33),
.B2(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_1),
.B(n_75),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_1),
.A2(n_57),
.B(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_3),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_60),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_60),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_68),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_53),
.B1(n_59),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_63),
.Y(n_194)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_7),
.A2(n_53),
.B1(n_59),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_119),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_119),
.Y(n_177)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_8),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_46),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_12),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_14),
.A2(n_40),
.A3(n_57),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_15),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_29),
.B1(n_31),
.B2(n_41),
.Y(n_42)
);

BUFx3_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_98),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_21),
.B(n_98),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_76),
.B2(n_77),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_47),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_27),
.A2(n_34),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_27),
.A2(n_33),
.B1(n_88),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_27),
.A2(n_80),
.B1(n_111),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_27),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_27),
.A2(n_33),
.B1(n_162),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_27),
.A2(n_33),
.B1(n_164),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_27),
.A2(n_28),
.B1(n_151),
.B2(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_31),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_37),
.A2(n_42),
.B1(n_45),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_37),
.A2(n_42),
.B1(n_43),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_37),
.A2(n_42),
.B1(n_90),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_37),
.A2(n_42),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_37),
.A2(n_42),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_37),
.A2(n_42),
.B1(n_192),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_37),
.A2(n_42),
.B1(n_130),
.B2(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_39),
.B(n_71),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_40),
.A2(n_41),
.B(n_108),
.C(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_42),
.B(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_58),
.B1(n_61),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_50),
.A2(n_61),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_51),
.A2(n_55),
.B1(n_107),
.B2(n_118),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_53),
.B(n_108),
.CON(n_107),
.SN(n_107)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_56),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_56),
.B(n_108),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_69),
.A2(n_75),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_73),
.B1(n_93),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_73),
.B1(n_114),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_70),
.A2(n_73),
.B1(n_146),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_80),
.B(n_108),
.Y(n_180)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_94),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_89),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_99),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_103),
.A2(n_104),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.C(n_115),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_152),
.B(n_235),
.C(n_241),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_137),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_124),
.B(n_137),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_126),
.B(n_127),
.C(n_135),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_138),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_234),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_229),
.B(n_233),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_215),
.B(n_228),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_196),
.B(n_214),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_184),
.B(n_195),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_173),
.B(n_183),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_165),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_201),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_225),
.C(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);


endmodule