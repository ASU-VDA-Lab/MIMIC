module fake_jpeg_13148_n_359 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_13),
.B(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_53),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_39),
.B1(n_27),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_74),
.B1(n_16),
.B2(n_35),
.Y(n_106)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_16),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_72),
.B1(n_75),
.B2(n_22),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_29),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_26),
.B1(n_16),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_21),
.B1(n_30),
.B2(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_33),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_40),
.B(n_29),
.CON(n_79),
.SN(n_79)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_81),
.B(n_22),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_25),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_51),
.B1(n_26),
.B2(n_33),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_84),
.A2(n_97),
.B(n_101),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_89),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_81),
.B1(n_66),
.B2(n_41),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_117),
.B1(n_32),
.B2(n_23),
.Y(n_140)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_29),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_103),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_109),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_20),
.B1(n_25),
.B2(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_57),
.B1(n_80),
.B2(n_71),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_13),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_45),
.B1(n_38),
.B2(n_58),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_22),
.B(n_58),
.C(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_17),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_49),
.B1(n_47),
.B2(n_45),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_19),
.B1(n_32),
.B2(n_35),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_80),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_106),
.B1(n_84),
.B2(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_135),
.B1(n_146),
.B2(n_148),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_69),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_63),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_63),
.C(n_73),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_73),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_151),
.B(n_105),
.C(n_116),
.D(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_98),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_113),
.B(n_100),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_85),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_34),
.B1(n_23),
.B2(n_17),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_71),
.B1(n_80),
.B2(n_19),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_19),
.B1(n_34),
.B2(n_32),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_35),
.C(n_34),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_101),
.B1(n_115),
.B2(n_88),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_157),
.B1(n_175),
.B2(n_178),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_155),
.B(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_156),
.B(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_102),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_166),
.Y(n_188)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_124),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_126),
.B1(n_146),
.B2(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_147),
.B1(n_135),
.B2(n_133),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_105),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_91),
.B1(n_90),
.B2(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_104),
.B1(n_96),
.B2(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_103),
.B1(n_17),
.B2(n_31),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_0),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_12),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_12),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_103),
.B(n_1),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_103),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_132),
.B1(n_137),
.B2(n_143),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_203),
.B1(n_222),
.B2(n_181),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_200),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_131),
.B1(n_130),
.B2(n_148),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_131),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_129),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_213),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_141),
.B1(n_129),
.B2(n_120),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_141),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_120),
.C(n_1),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_209),
.B(n_199),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_152),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_3),
.C(n_4),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_165),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_154),
.B1(n_155),
.B2(n_162),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_234),
.B1(n_245),
.B2(n_242),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_239),
.B(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_241),
.C(n_212),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_219),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_180),
.B1(n_178),
.B2(n_175),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_169),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_186),
.B(n_172),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_156),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_184),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_187),
.B1(n_179),
.B2(n_176),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_251),
.B1(n_222),
.B2(n_196),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_205),
.A2(n_174),
.B(n_153),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_157),
.B1(n_168),
.B2(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_198),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_246),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_194),
.B(n_163),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_197),
.B1(n_221),
.B2(n_206),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_204),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_252),
.A2(n_258),
.B1(n_265),
.B2(n_275),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_200),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_228),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_212),
.CI(n_214),
.CON(n_261),
.SN(n_261)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_261),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_197),
.B(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_195),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_236),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_202),
.C(n_211),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_208),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_211),
.C(n_206),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.C(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_217),
.C(n_208),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_204),
.B1(n_208),
.B2(n_215),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_215),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_289),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_225),
.B1(n_234),
.B2(n_224),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_250),
.B1(n_233),
.B2(n_237),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_282),
.B1(n_284),
.B2(n_291),
.Y(n_299)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_233),
.B1(n_240),
.B2(n_243),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_239),
.B1(n_227),
.B2(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_294),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_287),
.B(n_10),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_238),
.C(n_229),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_290),
.C(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_5),
.C(n_6),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_256),
.B(n_7),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_298),
.B(n_302),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_259),
.C(n_253),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_271),
.B1(n_263),
.B2(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_295),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_261),
.A3(n_254),
.B1(n_266),
.B2(n_269),
.C(n_265),
.Y(n_307)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_269),
.C(n_8),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_290),
.C(n_289),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_7),
.B(n_9),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_279),
.B(n_10),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_9),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_10),
.Y(n_324)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_320),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_319),
.B(n_302),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_288),
.C(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_299),
.B(n_304),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_314),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_329),
.B(n_331),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_322),
.B(n_303),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_334),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_305),
.B(n_310),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g335 ( 
.A1(n_315),
.A2(n_317),
.B(n_318),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_335),
.A2(n_315),
.B1(n_300),
.B2(n_316),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_298),
.C(n_312),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_344),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_345),
.A2(n_340),
.B(n_323),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_312),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_333),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_349),
.A2(n_350),
.B(n_352),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_348),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_351),
.Y(n_355)
);

A2O1A1O1Ixp25_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_345),
.B(n_346),
.C(n_341),
.D(n_354),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_356),
.A2(n_321),
.B1(n_335),
.B2(n_319),
.Y(n_357)
);

AOI221xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_330),
.B1(n_334),
.B2(n_10),
.C(n_11),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_11),
.Y(n_359)
);


endmodule