module fake_netlist_5_287_n_134 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_134);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_134;

wire n_91;
wire n_82;
wire n_122;
wire n_124;
wire n_86;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_101;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_30;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_29;
wire n_79;
wire n_131;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_26;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_R g53 ( 
.A(n_29),
.B(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_30),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_41),
.B1(n_37),
.B2(n_35),
.Y(n_61)
);

OR2x6_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_27),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_44),
.B(n_52),
.C(n_50),
.Y(n_65)
);

AO31x2_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_55),
.A3(n_58),
.B(n_46),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_40),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_50),
.B(n_46),
.Y(n_70)
);

OAI21x1_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_51),
.B(n_48),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_62),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_19),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_20),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_56),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_12),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_65),
.B1(n_68),
.B2(n_56),
.Y(n_78)
);

AOI21x1_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_60),
.B(n_6),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_23),
.B(n_24),
.Y(n_80)
);

AOI21x1_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_60),
.B(n_8),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_3),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_8),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_77),
.B(n_74),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_78),
.B(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_74),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_88),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_97),
.C(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_103),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_84),
.B1(n_74),
.B2(n_93),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

OAI322xp33_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_75),
.A3(n_90),
.B1(n_87),
.B2(n_92),
.C1(n_9),
.C2(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_102),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_74),
.C(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_102),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_75),
.B1(n_113),
.B2(n_108),
.C(n_114),
.Y(n_120)
);

OAI211xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_99),
.B(n_106),
.C(n_96),
.Y(n_121)
);

OAI221xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_99),
.B1(n_89),
.B2(n_96),
.C(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_115),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_121),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_9),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_125),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_122),
.A3(n_118),
.B1(n_79),
.B2(n_81),
.C1(n_80),
.C2(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_96),
.B(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_130),
.B1(n_80),
.B2(n_79),
.Y(n_134)
);


endmodule