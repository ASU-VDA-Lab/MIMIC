module fake_jpeg_26825_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_4),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_0),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_66),
.C(n_70),
.Y(n_87)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_57),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_56),
.B1(n_76),
.B2(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_90),
.B1(n_53),
.B2(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_73),
.B1(n_49),
.B2(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_49),
.B1(n_60),
.B2(n_69),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_105),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_108),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_106),
.B1(n_83),
.B2(n_78),
.Y(n_112)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_57),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_81),
.B1(n_50),
.B2(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_90),
.B1(n_83),
.B2(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_118),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_65),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_51),
.A3(n_52),
.B1(n_61),
.B2(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_1),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_85),
.C(n_107),
.Y(n_128)
);

XOR2x1_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_64),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_111),
.B1(n_110),
.B2(n_98),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_131),
.Y(n_140)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_3),
.B(n_5),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_2),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_84),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_7),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_50),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_141),
.B(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_121),
.C(n_63),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.C(n_28),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_63),
.C(n_23),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_9),
.B(n_10),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_26),
.C(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_13),
.B(n_14),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_15),
.C(n_16),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_18),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B1(n_137),
.B2(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_159),
.C(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_138),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_160),
.B1(n_157),
.B2(n_30),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_144),
.CI(n_25),
.CON(n_167),
.SN(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_19),
.B(n_32),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_167),
.B(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_33),
.Y(n_170)
);

AO21x2_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_36),
.B(n_37),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_38),
.CI(n_39),
.CON(n_172),
.SN(n_172)
);


endmodule