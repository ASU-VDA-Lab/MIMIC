module real_aes_9665_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_2043;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_2014;
wire n_1314;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_2035;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_2040;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_2049;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_2004;
wire n_1201;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_2038;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_2041;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_2050;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_2012;
wire n_1018;
wire n_1563;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2045;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_2036;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_1971;
wire n_964;
wire n_731;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2039;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_2023;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_2052;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_2019;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_2042;
wire n_1066;
wire n_2046;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_2048;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_2053;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_2055;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1931;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_2037;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_2030;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_2044;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1584;
wire n_1277;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_2047;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_2010;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_2051;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_2054;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_0), .A2(n_338), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
INVx1_ASAP7_75t_L g1290 ( .A(n_0), .Y(n_1290) );
AOI22xp5_ASAP7_75t_L g1741 ( .A1(n_1), .A2(n_360), .B1(n_1727), .B2(n_1730), .Y(n_1741) );
INVx1_ASAP7_75t_L g1656 ( .A(n_2), .Y(n_1656) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_3), .A2(n_259), .B1(n_527), .B2(n_604), .C(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g635 ( .A(n_3), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_4), .A2(n_123), .B1(n_1411), .B2(n_1413), .Y(n_1463) );
INVx1_ASAP7_75t_L g1500 ( .A(n_4), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_5), .A2(n_330), .B1(n_456), .B2(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g540 ( .A(n_5), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g1259 ( .A(n_6), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_7), .A2(n_216), .B1(n_527), .B2(n_737), .C(n_738), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_7), .A2(n_332), .B1(n_460), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g1559 ( .A(n_8), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_8), .A2(n_130), .B1(n_1267), .B2(n_1577), .Y(n_1576) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_9), .A2(n_36), .B1(n_656), .B2(n_1137), .C(n_1139), .Y(n_1136) );
INVx1_ASAP7_75t_L g1174 ( .A(n_9), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1531 ( .A1(n_10), .A2(n_121), .B1(n_485), .B2(n_516), .Y(n_1531) );
AOI221xp5_ASAP7_75t_L g1537 ( .A1(n_10), .A2(n_121), .B1(n_1103), .B2(n_1365), .C(n_1538), .Y(n_1537) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_11), .A2(n_22), .B1(n_1013), .B2(n_1017), .Y(n_1016) );
INVxp67_ASAP7_75t_SL g1022 ( .A(n_11), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_12), .A2(n_137), .B1(n_1373), .B2(n_1567), .Y(n_1566) );
AOI22xp33_ASAP7_75t_SL g1573 ( .A1(n_12), .A2(n_137), .B1(n_1107), .B2(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1200 ( .A(n_13), .Y(n_1200) );
OAI211xp5_ASAP7_75t_SL g1224 ( .A1(n_13), .A2(n_516), .B(n_1225), .C(n_1234), .Y(n_1224) );
INVx1_ASAP7_75t_L g1083 ( .A(n_14), .Y(n_1083) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_14), .A2(n_299), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
INVx1_ASAP7_75t_L g425 ( .A(n_15), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_16), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_17), .A2(n_90), .B1(n_1411), .B2(n_1413), .Y(n_1410) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_17), .A2(n_202), .B1(n_390), .B2(n_1045), .Y(n_1420) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_18), .A2(n_42), .B1(n_609), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_18), .A2(n_42), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g2024 ( .A(n_19), .Y(n_2024) );
AOI22xp5_ASAP7_75t_L g1742 ( .A1(n_20), .A2(n_319), .B1(n_1720), .B2(n_1738), .Y(n_1742) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_21), .Y(n_595) );
INVxp33_ASAP7_75t_L g1043 ( .A(n_22), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_23), .Y(n_824) );
INVx1_ASAP7_75t_L g859 ( .A(n_24), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_24), .A2(n_235), .B1(n_668), .B2(n_926), .C(n_928), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_25), .A2(n_108), .B1(n_581), .B2(n_663), .Y(n_815) );
INVx1_ASAP7_75t_L g840 ( .A(n_25), .Y(n_840) );
CKINVDCx16_ASAP7_75t_R g1718 ( .A(n_26), .Y(n_1718) );
AOI22xp33_ASAP7_75t_SL g1568 ( .A1(n_27), .A2(n_116), .B1(n_1373), .B2(n_1569), .Y(n_1568) );
INVxp67_ASAP7_75t_SL g1592 ( .A(n_27), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_28), .A2(n_372), .B1(n_693), .B2(n_695), .Y(n_692) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_28), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_29), .A2(n_152), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx1_ASAP7_75t_L g1153 ( .A(n_29), .Y(n_1153) );
INVx1_ASAP7_75t_L g1405 ( .A(n_30), .Y(n_1405) );
OAI222xp33_ASAP7_75t_L g1417 ( .A1(n_30), .A2(n_247), .B1(n_345), .B2(n_1031), .C1(n_1418), .C2(n_1419), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_31), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_32), .A2(n_223), .B1(n_427), .B2(n_707), .Y(n_760) );
INVx1_ASAP7_75t_L g786 ( .A(n_32), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g1367 ( .A1(n_33), .A2(n_149), .B1(n_1095), .B2(n_1265), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_33), .A2(n_149), .B1(n_600), .B2(n_733), .Y(n_1379) );
OAI22xp5_ASAP7_75t_L g1942 ( .A1(n_34), .A2(n_355), .B1(n_1943), .B2(n_1944), .Y(n_1942) );
INVxp67_ASAP7_75t_SL g1994 ( .A(n_34), .Y(n_1994) );
INVx1_ASAP7_75t_L g618 ( .A(n_35), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_35), .A2(n_320), .B1(n_668), .B2(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g1169 ( .A(n_36), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_37), .A2(n_91), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g638 ( .A(n_37), .Y(n_638) );
INVx1_ASAP7_75t_L g610 ( .A(n_38), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_38), .A2(n_187), .B1(n_660), .B2(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g1352 ( .A(n_39), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_39), .A2(n_348), .B1(n_609), .B2(n_737), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1462 ( .A(n_40), .B(n_1409), .Y(n_1462) );
INVx1_ASAP7_75t_L g1498 ( .A(n_40), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_41), .Y(n_1197) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_43), .Y(n_1065) );
INVx1_ASAP7_75t_L g381 ( .A(n_44), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_45), .A2(n_135), .B1(n_546), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g652 ( .A(n_45), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_46), .A2(n_136), .B1(n_1408), .B2(n_1409), .Y(n_1407) );
AOI22xp33_ASAP7_75t_SL g1428 ( .A1(n_46), .A2(n_136), .B1(n_600), .B2(n_1375), .Y(n_1428) );
INVx1_ASAP7_75t_L g1659 ( .A(n_47), .Y(n_1659) );
OAI211xp5_ASAP7_75t_SL g1682 ( .A1(n_47), .A2(n_516), .B(n_1683), .C(n_1687), .Y(n_1682) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_48), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_49), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_50), .A2(n_177), .B1(n_1727), .B2(n_1730), .Y(n_1726) );
XOR2xp5_ASAP7_75t_L g405 ( .A(n_51), .B(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g1822 ( .A1(n_51), .A2(n_238), .B1(n_1714), .B2(n_1781), .Y(n_1822) );
INVxp67_ASAP7_75t_SL g1560 ( .A(n_52), .Y(n_1560) );
OAI22xp33_ASAP7_75t_L g1584 ( .A1(n_52), .A2(n_196), .B1(n_1355), .B2(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1950 ( .A(n_53), .Y(n_1950) );
OAI221xp5_ASAP7_75t_L g1970 ( .A1(n_53), .A2(n_325), .B1(n_1971), .B2(n_1973), .C(n_1975), .Y(n_1970) );
INVx1_ASAP7_75t_L g1599 ( .A(n_54), .Y(n_1599) );
AOI22xp33_ASAP7_75t_L g1629 ( .A1(n_54), .A2(n_234), .B1(n_737), .B2(n_1316), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_55), .A2(n_307), .B1(n_693), .B2(n_695), .Y(n_765) );
INVx1_ASAP7_75t_L g799 ( .A(n_55), .Y(n_799) );
INVx1_ASAP7_75t_L g1306 ( .A(n_56), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_56), .A2(n_302), .B1(n_849), .B2(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1422 ( .A(n_57), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_57), .A2(n_243), .B1(n_693), .B2(n_695), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1625 ( .A1(n_58), .A2(n_170), .B1(n_1282), .B2(n_1316), .Y(n_1625) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_58), .A2(n_170), .B1(n_1100), .B2(n_1365), .Y(n_1632) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_59), .A2(n_262), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
INVx1_ASAP7_75t_L g1287 ( .A(n_59), .Y(n_1287) );
AOI22x1_ASAP7_75t_SL g1397 ( .A1(n_60), .A2(n_1398), .B1(n_1437), .B2(n_1438), .Y(n_1397) );
INVx1_ASAP7_75t_L g1437 ( .A(n_60), .Y(n_1437) );
AO221x2_ASAP7_75t_L g1744 ( .A1(n_60), .A2(n_275), .B1(n_1720), .B2(n_1738), .C(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g826 ( .A(n_61), .Y(n_826) );
CKINVDCx16_ASAP7_75t_R g1721 ( .A(n_62), .Y(n_1721) );
AOI22xp33_ASAP7_75t_L g2000 ( .A1(n_62), .A2(n_2001), .B1(n_2005), .B2(n_2048), .Y(n_2000) );
AOI22xp5_ASAP7_75t_L g1736 ( .A1(n_63), .A2(n_154), .B1(n_1727), .B2(n_1730), .Y(n_1736) );
INVx1_ASAP7_75t_L g1116 ( .A(n_64), .Y(n_1116) );
XNOR2xp5_ASAP7_75t_L g1182 ( .A(n_65), .B(n_1183), .Y(n_1182) );
AOI22xp5_ASAP7_75t_SL g1758 ( .A1(n_65), .A2(n_251), .B1(n_1714), .B2(n_1720), .Y(n_1758) );
OAI22xp33_ASAP7_75t_L g1667 ( .A1(n_66), .A2(n_260), .B1(n_456), .B2(n_460), .Y(n_1667) );
INVx1_ASAP7_75t_L g1685 ( .A(n_66), .Y(n_1685) );
INVx1_ASAP7_75t_L g823 ( .A(n_67), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_67), .A2(n_215), .B1(n_604), .B2(n_781), .C(n_782), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_68), .A2(n_80), .B1(n_999), .B2(n_1001), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_68), .A2(n_80), .B1(n_704), .B2(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g509 ( .A(n_69), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_69), .A2(n_245), .B1(n_568), .B2(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g688 ( .A(n_70), .Y(n_688) );
INVx1_ASAP7_75t_L g1360 ( .A(n_71), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_71), .A2(n_200), .B1(n_1373), .B2(n_1375), .Y(n_1372) );
INVx1_ASAP7_75t_L g892 ( .A(n_72), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_72), .A2(n_191), .B1(n_668), .B2(n_938), .C(n_940), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_73), .A2(n_249), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_73), .A2(n_249), .B1(n_656), .B2(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g2039 ( .A(n_74), .Y(n_2039) );
OAI22xp33_ASAP7_75t_L g2045 ( .A1(n_74), .A2(n_150), .B1(n_460), .B2(n_745), .Y(n_2045) );
INVx1_ASAP7_75t_L g1324 ( .A(n_75), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_75), .A2(n_293), .B1(n_693), .B2(n_695), .Y(n_1346) );
INVxp33_ASAP7_75t_L g976 ( .A(n_76), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_76), .A2(n_161), .B1(n_601), .B2(n_999), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_77), .A2(n_359), .B1(n_587), .B2(n_770), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_77), .A2(n_359), .B1(n_549), .B2(n_554), .Y(n_800) );
INVx1_ASAP7_75t_L g1326 ( .A(n_78), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_78), .A2(n_328), .B1(n_581), .B2(n_663), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g2015 ( .A1(n_79), .A2(n_374), .B1(n_577), .B2(n_693), .Y(n_2015) );
INVx1_ASAP7_75t_L g2030 ( .A(n_79), .Y(n_2030) );
CKINVDCx14_ASAP7_75t_R g1786 ( .A(n_81), .Y(n_1786) );
AOI22xp33_ASAP7_75t_L g1961 ( .A1(n_82), .A2(n_224), .B1(n_814), .B2(n_1962), .Y(n_1961) );
AOI22xp33_ASAP7_75t_L g1982 ( .A1(n_82), .A2(n_224), .B1(n_1333), .B2(n_1983), .Y(n_1982) );
INVx1_ASAP7_75t_L g496 ( .A(n_83), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_83), .A2(n_211), .B1(n_574), .B2(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g1514 ( .A(n_84), .Y(n_1514) );
AOI221xp5_ASAP7_75t_L g1533 ( .A1(n_84), .A2(n_268), .B1(n_1365), .B2(n_1534), .C(n_1536), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_85), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_86), .A2(n_336), .B1(n_549), .B2(n_554), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_86), .A2(n_336), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_L g1312 ( .A(n_87), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_87), .A2(n_346), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
INVx1_ASAP7_75t_L g768 ( .A(n_88), .Y(n_768) );
OAI211xp5_ASAP7_75t_SL g774 ( .A1(n_88), .A2(n_516), .B(n_775), .C(n_783), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1623 ( .A1(n_89), .A2(n_212), .B1(n_1373), .B2(n_1624), .Y(n_1623) );
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_89), .A2(n_212), .B1(n_658), .B2(n_1574), .Y(n_1631) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_90), .A2(n_166), .B1(n_1316), .B2(n_1333), .Y(n_1429) );
INVx1_ASAP7_75t_L g636 ( .A(n_91), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_92), .A2(n_311), .B1(n_451), .B2(n_582), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_92), .A2(n_485), .B1(n_725), .B2(n_838), .C(n_844), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g1820 ( .A1(n_93), .A2(n_226), .B1(n_1727), .B2(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g466 ( .A(n_94), .Y(n_466) );
INVx1_ASAP7_75t_L g972 ( .A(n_95), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_96), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_97), .Y(n_1252) );
AOI22xp33_ASAP7_75t_SL g1426 ( .A1(n_98), .A2(n_173), .B1(n_1233), .B2(n_1316), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_98), .A2(n_173), .B1(n_581), .B2(n_582), .Y(n_1432) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_99), .A2(n_361), .B1(n_708), .B2(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1236 ( .A(n_99), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_100), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_101), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_102), .A2(n_264), .B1(n_1132), .B2(n_1133), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_102), .A2(n_264), .B1(n_878), .B2(n_881), .C(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1664 ( .A(n_103), .Y(n_1664) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_103), .A2(n_242), .B1(n_711), .B2(n_712), .Y(n_1672) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_104), .A2(n_366), .B1(n_1103), .B2(n_1268), .Y(n_1269) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_104), .A2(n_485), .B1(n_725), .B2(n_1286), .C(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1600 ( .A(n_105), .Y(n_1600) );
AOI22xp33_ASAP7_75t_L g1627 ( .A1(n_105), .A2(n_188), .B1(n_1373), .B2(n_1628), .Y(n_1627) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_106), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g2014 ( .A(n_107), .Y(n_2014) );
INVx1_ASAP7_75t_L g843 ( .A(n_108), .Y(n_843) );
INVxp33_ASAP7_75t_SL g1966 ( .A(n_109), .Y(n_1966) );
AOI22xp33_ASAP7_75t_L g1987 ( .A1(n_109), .A2(n_353), .B1(n_1983), .B2(n_1985), .Y(n_1987) );
INVx1_ASAP7_75t_L g1206 ( .A(n_110), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_110), .A2(n_312), .B1(n_711), .B2(n_712), .Y(n_1214) );
CKINVDCx14_ASAP7_75t_R g1746 ( .A(n_111), .Y(n_1746) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_112), .Y(n_678) );
XNOR2x2_ASAP7_75t_L g1505 ( .A(n_113), .B(n_1506), .Y(n_1505) );
INVxp67_ASAP7_75t_SL g1554 ( .A(n_114), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_114), .A2(n_273), .B1(n_1574), .B2(n_1580), .Y(n_1579) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_115), .Y(n_1524) );
INVxp33_ASAP7_75t_L g1591 ( .A(n_116), .Y(n_1591) );
INVx1_ASAP7_75t_L g424 ( .A(n_117), .Y(n_424) );
BUFx2_ASAP7_75t_L g469 ( .A(n_117), .Y(n_469) );
BUFx2_ASAP7_75t_L g474 ( .A(n_117), .Y(n_474) );
OR2x2_ASAP7_75t_L g877 ( .A(n_117), .B(n_479), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_118), .A2(n_254), .B1(n_626), .B2(n_1375), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_118), .A2(n_254), .B1(n_669), .B2(n_813), .Y(n_1431) );
INVx1_ASAP7_75t_L g777 ( .A(n_119), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_119), .A2(n_208), .B1(n_747), .B2(n_749), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_120), .A2(n_356), .B1(n_1100), .B2(n_1365), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_120), .A2(n_356), .B1(n_737), .B2(n_1381), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_122), .A2(n_370), .B1(n_626), .B2(n_627), .Y(n_1335) );
AOI22xp33_ASAP7_75t_SL g1343 ( .A1(n_122), .A2(n_370), .B1(n_770), .B2(n_814), .Y(n_1343) );
INVx1_ASAP7_75t_L g1455 ( .A(n_123), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_124), .A2(n_179), .B1(n_1311), .B2(n_1355), .Y(n_1354) );
OAI22xp33_ASAP7_75t_L g1390 ( .A1(n_124), .A2(n_179), .B1(n_1029), .B2(n_1321), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_125), .Y(n_1512) );
INVx1_ASAP7_75t_L g1255 ( .A(n_126), .Y(n_1255) );
AOI221xp5_ASAP7_75t_L g1280 ( .A1(n_126), .A2(n_306), .B1(n_527), .B2(n_1281), .C(n_1282), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_127), .A2(n_203), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_127), .A2(n_203), .B1(n_660), .B2(n_663), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_128), .A2(n_220), .B1(n_737), .B2(n_780), .Y(n_1570) );
INVxp67_ASAP7_75t_SL g1583 ( .A(n_128), .Y(n_1583) );
INVx1_ASAP7_75t_L g1308 ( .A(n_129), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_129), .A2(n_145), .B1(n_622), .B2(n_1340), .Y(n_1339) );
INVxp33_ASAP7_75t_L g1556 ( .A(n_130), .Y(n_1556) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_131), .A2(n_485), .B1(n_490), .B2(n_502), .C(n_512), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_131), .A2(n_279), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_132), .A2(n_285), .B1(n_581), .B2(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1175 ( .A(n_132), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_133), .A2(n_208), .B1(n_737), .B2(n_780), .C(n_782), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_133), .A2(n_256), .B1(n_460), .B2(n_745), .Y(n_802) );
INVxp67_ASAP7_75t_SL g979 ( .A(n_134), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g1006 ( .A1(n_134), .A2(n_228), .B1(n_607), .B2(n_1004), .Y(n_1006) );
INVx1_ASAP7_75t_L g651 ( .A(n_135), .Y(n_651) );
XNOR2x2_ASAP7_75t_L g1297 ( .A(n_138), .B(n_1298), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_139), .A2(n_231), .B1(n_693), .B2(n_695), .Y(n_1019) );
INVxp33_ASAP7_75t_SL g1036 ( .A(n_139), .Y(n_1036) );
INVx1_ASAP7_75t_L g1658 ( .A(n_140), .Y(n_1658) );
OAI221xp5_ASAP7_75t_L g1673 ( .A1(n_140), .A2(n_485), .B1(n_725), .B2(n_1674), .C(n_1678), .Y(n_1673) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_141), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_142), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_143), .A2(n_169), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g845 ( .A(n_143), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g2021 ( .A1(n_144), .A2(n_210), .B1(n_427), .B2(n_2022), .Y(n_2021) );
INVx1_ASAP7_75t_L g2043 ( .A(n_144), .Y(n_2043) );
INVx1_ASAP7_75t_L g1301 ( .A(n_145), .Y(n_1301) );
OA22x2_ASAP7_75t_L g1443 ( .A1(n_146), .A2(n_1444), .B1(n_1503), .B2(n_1504), .Y(n_1443) );
INVxp67_ASAP7_75t_SL g1504 ( .A(n_146), .Y(n_1504) );
INVx1_ASAP7_75t_L g731 ( .A(n_147), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_147), .A2(n_216), .B1(n_747), .B2(n_749), .Y(n_746) );
XNOR2xp5_ASAP7_75t_L g1246 ( .A(n_148), .B(n_1247), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g2040 ( .A1(n_150), .A2(n_321), .B1(n_737), .B2(n_738), .C(n_1522), .Y(n_2040) );
CKINVDCx5p33_ASAP7_75t_R g1070 ( .A(n_151), .Y(n_1070) );
INVx1_ASAP7_75t_L g1158 ( .A(n_152), .Y(n_1158) );
INVx1_ASAP7_75t_L g700 ( .A(n_153), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_153), .A2(n_485), .B1(n_714), .B2(n_721), .C(n_725), .Y(n_713) );
INVx1_ASAP7_75t_L g454 ( .A(n_155), .Y(n_454) );
INVx1_ASAP7_75t_L g1615 ( .A(n_156), .Y(n_1615) );
AOI22xp33_ASAP7_75t_SL g1634 ( .A1(n_156), .A2(n_331), .B1(n_1365), .B2(n_1635), .Y(n_1634) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_157), .A2(n_181), .B1(n_1271), .B2(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1392 ( .A(n_157), .Y(n_1392) );
CKINVDCx5p33_ASAP7_75t_R g1518 ( .A(n_158), .Y(n_1518) );
AOI221xp5_ASAP7_75t_L g1957 ( .A1(n_159), .A2(n_329), .B1(n_1264), .B2(n_1958), .C(n_1959), .Y(n_1957) );
AOI22xp33_ASAP7_75t_L g1984 ( .A1(n_159), .A2(n_329), .B1(n_1985), .B2(n_1986), .Y(n_1984) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_160), .A2(n_303), .B1(n_549), .B2(n_554), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_160), .A2(n_303), .B1(n_584), .B2(n_587), .Y(n_583) );
INVxp33_ASAP7_75t_SL g967 ( .A(n_161), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_162), .A2(n_214), .B1(n_1095), .B2(n_1271), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1293 ( .A1(n_162), .A2(n_214), .B1(n_549), .B2(n_554), .Y(n_1293) );
INVx1_ASAP7_75t_L g1079 ( .A(n_163), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_163), .A2(n_304), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g1256 ( .A(n_164), .Y(n_1256) );
INVx1_ASAP7_75t_L g2038 ( .A(n_165), .Y(n_2038) );
OAI22xp33_ASAP7_75t_L g2046 ( .A1(n_165), .A2(n_321), .B1(n_747), .B2(n_749), .Y(n_2046) );
INVx1_ASAP7_75t_L g1402 ( .A(n_166), .Y(n_1402) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_167), .Y(n_1456) );
AOI22xp5_ASAP7_75t_SL g1757 ( .A1(n_168), .A2(n_185), .B1(n_1727), .B2(n_1730), .Y(n_1757) );
INVx1_ASAP7_75t_L g847 ( .A(n_169), .Y(n_847) );
INVxp33_ASAP7_75t_SL g1965 ( .A(n_171), .Y(n_1965) );
AOI22xp33_ASAP7_75t_L g1988 ( .A1(n_171), .A2(n_313), .B1(n_1333), .B2(n_1986), .Y(n_1988) );
INVx1_ASAP7_75t_L g1704 ( .A(n_172), .Y(n_1704) );
INVx1_ASAP7_75t_L g1610 ( .A(n_174), .Y(n_1610) );
AOI22xp33_ASAP7_75t_L g1636 ( .A1(n_174), .A2(n_209), .B1(n_442), .B2(n_658), .Y(n_1636) );
CKINVDCx16_ASAP7_75t_R g1711 ( .A(n_175), .Y(n_1711) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_176), .A2(n_296), .B1(n_693), .B2(n_695), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_176), .A2(n_296), .B1(n_549), .B2(n_712), .Y(n_850) );
INVx1_ASAP7_75t_L g1088 ( .A(n_178), .Y(n_1088) );
INVx1_ASAP7_75t_L g1557 ( .A(n_180), .Y(n_1557) );
INVx1_ASAP7_75t_L g1394 ( .A(n_181), .Y(n_1394) );
INVx1_ASAP7_75t_L g1651 ( .A(n_182), .Y(n_1651) );
INVx1_ASAP7_75t_L g1705 ( .A(n_183), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_183), .B(n_1703), .Y(n_1710) );
INVx1_ASAP7_75t_L g980 ( .A(n_184), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_184), .A2(n_365), .B1(n_1029), .B2(n_1031), .Y(n_1028) );
INVx2_ASAP7_75t_L g393 ( .A(n_186), .Y(n_393) );
INVx1_ASAP7_75t_L g629 ( .A(n_187), .Y(n_629) );
INVx1_ASAP7_75t_L g1603 ( .A(n_188), .Y(n_1603) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_189), .A2(n_222), .B1(n_707), .B2(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g740 ( .A(n_189), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g1476 ( .A(n_190), .Y(n_1476) );
INVx1_ASAP7_75t_L g894 ( .A(n_191), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g2019 ( .A1(n_192), .A2(n_367), .B1(n_658), .B2(n_2020), .Y(n_2019) );
OAI22xp5_ASAP7_75t_L g2026 ( .A1(n_192), .A2(n_367), .B1(n_549), .B2(n_554), .Y(n_2026) );
BUFx3_ASAP7_75t_L g432 ( .A(n_193), .Y(n_432) );
INVx1_ASAP7_75t_L g459 ( .A(n_193), .Y(n_459) );
INVx1_ASAP7_75t_L g897 ( .A(n_194), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_194), .A2(n_217), .B1(n_942), .B2(n_945), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_195), .Y(n_1469) );
INVx1_ASAP7_75t_L g1562 ( .A(n_196), .Y(n_1562) );
CKINVDCx5p33_ASAP7_75t_R g1460 ( .A(n_197), .Y(n_1460) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_198), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g1530 ( .A1(n_199), .A2(n_340), .B1(n_711), .B2(n_712), .Y(n_1530) );
INVx1_ASAP7_75t_L g1540 ( .A(n_199), .Y(n_1540) );
INVx1_ASAP7_75t_L g1361 ( .A(n_200), .Y(n_1361) );
OAI221xp5_ASAP7_75t_L g1604 ( .A1(n_201), .A2(n_267), .B1(n_1355), .B2(n_1605), .C(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1613 ( .A(n_201), .Y(n_1613) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_202), .A2(n_247), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
INVx1_ASAP7_75t_L g702 ( .A(n_204), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g726 ( .A1(n_204), .A2(n_516), .B(n_727), .C(n_739), .Y(n_726) );
XNOR2xp5_ASAP7_75t_L g804 ( .A(n_205), .B(n_805), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_206), .A2(n_218), .B1(n_1123), .B2(n_1124), .C(n_1125), .Y(n_1122) );
INVx1_ASAP7_75t_L g1157 ( .A(n_206), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_207), .A2(n_373), .B1(n_527), .B2(n_609), .C(n_1233), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_207), .A2(n_305), .B1(n_747), .B2(n_749), .Y(n_1239) );
INVx1_ASAP7_75t_L g1611 ( .A(n_209), .Y(n_1611) );
INVx1_ASAP7_75t_L g2042 ( .A(n_210), .Y(n_2042) );
INVx1_ASAP7_75t_L g501 ( .A(n_211), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_213), .Y(n_1066) );
INVx1_ASAP7_75t_L g821 ( .A(n_215), .Y(n_821) );
INVx1_ASAP7_75t_L g889 ( .A(n_217), .Y(n_889) );
INVx1_ASAP7_75t_L g1155 ( .A(n_218), .Y(n_1155) );
INVx1_ASAP7_75t_L g420 ( .A(n_219), .Y(n_420) );
INVx1_ASAP7_75t_L g566 ( .A(n_219), .Y(n_566) );
INVxp33_ASAP7_75t_L g1589 ( .A(n_220), .Y(n_1589) );
OAI22xp33_ASAP7_75t_L g1668 ( .A1(n_221), .A2(n_290), .B1(n_747), .B2(n_749), .Y(n_1668) );
AOI221xp5_ASAP7_75t_L g1686 ( .A1(n_221), .A2(n_260), .B1(n_606), .B2(n_865), .C(n_1522), .Y(n_1686) );
INVx1_ASAP7_75t_L g741 ( .A(n_222), .Y(n_741) );
INVx1_ASAP7_75t_L g784 ( .A(n_223), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g1480 ( .A(n_225), .Y(n_1480) );
CKINVDCx20_ASAP7_75t_R g1784 ( .A(n_227), .Y(n_1784) );
INVxp33_ASAP7_75t_SL g962 ( .A(n_228), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_229), .Y(n_1072) );
XOR2x2_ASAP7_75t_L g1057 ( .A(n_230), .B(n_1058), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1040 ( .A(n_231), .Y(n_1040) );
INVx1_ASAP7_75t_L g1199 ( .A(n_232), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_232), .A2(n_485), .B1(n_512), .B2(n_1216), .C(n_1223), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_233), .Y(n_1358) );
INVx1_ASAP7_75t_L g1607 ( .A(n_234), .Y(n_1607) );
INVx1_ASAP7_75t_L g869 ( .A(n_235), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_236), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_237), .Y(n_1528) );
OAI221xp5_ASAP7_75t_L g1541 ( .A1(n_237), .A2(n_410), .B1(n_427), .B2(n_647), .C(n_1542), .Y(n_1541) );
CKINVDCx14_ASAP7_75t_R g1747 ( .A(n_239), .Y(n_1747) );
INVx1_ASAP7_75t_L g449 ( .A(n_240), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g1653 ( .A(n_241), .Y(n_1653) );
INVx1_ASAP7_75t_L g1661 ( .A(n_242), .Y(n_1661) );
INVx1_ASAP7_75t_L g1423 ( .A(n_243), .Y(n_1423) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_244), .Y(n_1069) );
INVx1_ASAP7_75t_L g507 ( .A(n_245), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_246), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g1602 ( .A(n_248), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_250), .A2(n_337), .B1(n_607), .B2(n_1333), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1344 ( .A1(n_250), .A2(n_337), .B1(n_568), .B2(n_663), .Y(n_1344) );
INVx1_ASAP7_75t_L g2018 ( .A(n_252), .Y(n_2018) );
OAI211xp5_ASAP7_75t_SL g2036 ( .A1(n_252), .A2(n_516), .B(n_2037), .C(n_2041), .Y(n_2036) );
CKINVDCx16_ASAP7_75t_R g1548 ( .A(n_253), .Y(n_1548) );
INVx1_ASAP7_75t_L g772 ( .A(n_255), .Y(n_772) );
INVx1_ASAP7_75t_L g778 ( .A(n_256), .Y(n_778) );
INVx1_ASAP7_75t_L g2017 ( .A(n_257), .Y(n_2017) );
OAI221xp5_ASAP7_75t_L g2027 ( .A1(n_257), .A2(n_485), .B1(n_512), .B2(n_2028), .C(n_2035), .Y(n_2027) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_258), .Y(n_763) );
INVx1_ASAP7_75t_L g640 ( .A(n_259), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g854 ( .A(n_261), .B(n_855), .Y(n_854) );
XNOR2x1_ASAP7_75t_L g1050 ( .A(n_261), .B(n_855), .Y(n_1050) );
INVx1_ASAP7_75t_L g1288 ( .A(n_262), .Y(n_1288) );
INVx1_ASAP7_75t_L g1650 ( .A(n_263), .Y(n_1650) );
CKINVDCx5p33_ASAP7_75t_R g1520 ( .A(n_265), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_266), .A2(n_283), .B1(n_1448), .B2(n_1450), .Y(n_1447) );
INVx1_ASAP7_75t_L g1490 ( .A(n_266), .Y(n_1490) );
INVx1_ASAP7_75t_L g1614 ( .A(n_267), .Y(n_1614) );
AOI21xp33_ASAP7_75t_L g1515 ( .A1(n_268), .A2(n_480), .B(n_623), .Y(n_1515) );
CKINVDCx5p33_ASAP7_75t_R g2013 ( .A(n_269), .Y(n_2013) );
OAI221xp5_ASAP7_75t_L g1061 ( .A1(n_270), .A2(n_516), .B1(n_1062), .B2(n_1067), .C(n_1071), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_270), .A2(n_344), .B1(n_1101), .B2(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1148 ( .A(n_271), .Y(n_1148) );
OAI211xp5_ASAP7_75t_L g1451 ( .A1(n_272), .A2(n_789), .B(n_1452), .C(n_1453), .Y(n_1451) );
INVx1_ASAP7_75t_L g1487 ( .A(n_272), .Y(n_1487) );
INVx1_ASAP7_75t_L g1553 ( .A(n_273), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_274), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g872 ( .A1(n_276), .A2(n_364), .B1(n_873), .B2(n_878), .C(n_881), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_276), .A2(n_364), .B1(n_920), .B2(n_923), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g1706 ( .A(n_277), .Y(n_1706) );
BUFx3_ASAP7_75t_L g415 ( .A(n_278), .Y(n_415) );
INVx1_ASAP7_75t_L g445 ( .A(n_278), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_279), .A2(n_516), .B1(n_523), .B2(n_532), .C(n_541), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g757 ( .A(n_280), .B(n_758), .Y(n_757) );
AO221x2_ASAP7_75t_L g1780 ( .A1(n_280), .A2(n_349), .B1(n_1781), .B2(n_1782), .C(n_1783), .Y(n_1780) );
INVx1_ASAP7_75t_L g1670 ( .A(n_281), .Y(n_1670) );
AO22x2_ASAP7_75t_L g1595 ( .A1(n_282), .A2(n_1596), .B1(n_1637), .B2(n_1638), .Y(n_1595) );
INVxp67_ASAP7_75t_L g1637 ( .A(n_282), .Y(n_1637) );
AOI22xp5_ASAP7_75t_L g1737 ( .A1(n_282), .A2(n_288), .B1(n_1720), .B2(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1489 ( .A(n_283), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_284), .Y(n_905) );
INVx1_ASAP7_75t_L g1167 ( .A(n_285), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_286), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_286), .B(n_350), .Y(n_479) );
AND2x2_ASAP7_75t_L g487 ( .A(n_286), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g531 ( .A(n_286), .Y(n_531) );
XNOR2xp5_ASAP7_75t_L g1644 ( .A(n_287), .B(n_1645), .Y(n_1644) );
AOI21xp5_ASAP7_75t_L g1951 ( .A1(n_289), .A2(n_1125), .B(n_1952), .Y(n_1951) );
INVx1_ASAP7_75t_L g1978 ( .A(n_289), .Y(n_1978) );
INVx1_ASAP7_75t_L g1684 ( .A(n_290), .Y(n_1684) );
AO22x2_ASAP7_75t_L g957 ( .A1(n_291), .A2(n_958), .B1(n_959), .B2(n_1047), .Y(n_957) );
INVxp67_ASAP7_75t_SL g958 ( .A(n_291), .Y(n_958) );
AOI21xp33_ASAP7_75t_L g1521 ( .A1(n_292), .A2(n_1334), .B(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1544 ( .A(n_292), .Y(n_1544) );
INVx1_ASAP7_75t_L g1323 ( .A(n_293), .Y(n_1323) );
XNOR2xp5_ASAP7_75t_L g1348 ( .A(n_294), .B(n_1349), .Y(n_1348) );
INVx2_ASAP7_75t_L g422 ( .A(n_295), .Y(n_422) );
OR2x2_ASAP7_75t_L g448 ( .A(n_295), .B(n_420), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_297), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_298), .Y(n_1190) );
INVx1_ASAP7_75t_L g1086 ( .A(n_299), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_300), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g1474 ( .A(n_301), .Y(n_1474) );
INVx1_ASAP7_75t_L g1303 ( .A(n_302), .Y(n_1303) );
INVx1_ASAP7_75t_L g1076 ( .A(n_304), .Y(n_1076) );
INVx1_ASAP7_75t_L g1228 ( .A(n_305), .Y(n_1228) );
INVx1_ASAP7_75t_L g1253 ( .A(n_306), .Y(n_1253) );
INVx1_ASAP7_75t_L g795 ( .A(n_307), .Y(n_795) );
INVx1_ASAP7_75t_L g1231 ( .A(n_308), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_308), .A2(n_373), .B1(n_456), .B2(n_460), .Y(n_1238) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_309), .Y(n_1517) );
AOI22xp5_ASAP7_75t_SL g1732 ( .A1(n_310), .A2(n_315), .B1(n_1714), .B2(n_1720), .Y(n_1732) );
OAI211xp5_ASAP7_75t_SL g828 ( .A1(n_311), .A2(n_516), .B(n_829), .C(n_836), .Y(n_828) );
INVx1_ASAP7_75t_L g1203 ( .A(n_312), .Y(n_1203) );
INVxp67_ASAP7_75t_SL g1956 ( .A(n_313), .Y(n_1956) );
AOI22xp5_ASAP7_75t_L g2006 ( .A1(n_314), .A2(n_2007), .B1(n_2008), .B2(n_2047), .Y(n_2006) );
CKINVDCx5p33_ASAP7_75t_R g2007 ( .A(n_314), .Y(n_2007) );
AOI221xp5_ASAP7_75t_L g1946 ( .A1(n_316), .A2(n_325), .B1(n_814), .B2(n_1264), .C(n_1947), .Y(n_1946) );
INVxp33_ASAP7_75t_L g1976 ( .A(n_316), .Y(n_1976) );
CKINVDCx5p33_ASAP7_75t_R g1482 ( .A(n_317), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_318), .A2(n_339), .B1(n_1365), .B2(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1396 ( .A(n_318), .Y(n_1396) );
INVx1_ASAP7_75t_L g617 ( .A(n_320), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_322), .A2(n_351), .B1(n_587), .B2(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_322), .A2(n_351), .B1(n_711), .B2(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g675 ( .A(n_323), .Y(n_675) );
INVx1_ASAP7_75t_L g767 ( .A(n_324), .Y(n_767) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_324), .A2(n_485), .B1(n_725), .B2(n_788), .C(n_791), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_326), .A2(n_371), .B1(n_737), .B2(n_738), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_326), .A2(n_371), .B1(n_1015), .B2(n_1100), .Y(n_1575) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_327), .Y(n_1260) );
INVx1_ASAP7_75t_L g1318 ( .A(n_328), .Y(n_1318) );
INVx1_ASAP7_75t_L g525 ( .A(n_330), .Y(n_525) );
INVx1_ASAP7_75t_L g1620 ( .A(n_331), .Y(n_1620) );
INVx1_ASAP7_75t_L g735 ( .A(n_332), .Y(n_735) );
INVx1_ASAP7_75t_L g433 ( .A(n_333), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_334), .Y(n_1305) );
OAI22xp33_ASAP7_75t_L g1665 ( .A1(n_335), .A2(n_354), .B1(n_708), .B2(n_1209), .Y(n_1665) );
INVx1_ASAP7_75t_L g1689 ( .A(n_335), .Y(n_1689) );
INVx1_ASAP7_75t_L g1291 ( .A(n_338), .Y(n_1291) );
INVx1_ASAP7_75t_L g1389 ( .A(n_339), .Y(n_1389) );
INVx1_ASAP7_75t_L g1539 ( .A(n_340), .Y(n_1539) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_341), .B(n_381), .Y(n_1701) );
AND3x2_ASAP7_75t_L g1717 ( .A(n_341), .B(n_381), .C(n_1704), .Y(n_1717) );
CKINVDCx5p33_ASAP7_75t_R g1212 ( .A(n_342), .Y(n_1212) );
INVx2_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_344), .A2(n_485), .B1(n_512), .B2(n_1075), .C(n_1080), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_345), .Y(n_1404) );
INVx1_ASAP7_75t_L g1309 ( .A(n_346), .Y(n_1309) );
INVx1_ASAP7_75t_L g1273 ( .A(n_347), .Y(n_1273) );
INVx1_ASAP7_75t_L g1357 ( .A(n_348), .Y(n_1357) );
INVx1_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
INVx2_ASAP7_75t_L g488 ( .A(n_350), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_352), .Y(n_1446) );
INVxp67_ASAP7_75t_SL g1939 ( .A(n_353), .Y(n_1939) );
INVx1_ASAP7_75t_L g1688 ( .A(n_354), .Y(n_1688) );
INVxp67_ASAP7_75t_SL g1992 ( .A(n_355), .Y(n_1992) );
INVx1_ASAP7_75t_L g1527 ( .A(n_357), .Y(n_1527) );
HB1xp67_ASAP7_75t_L g1542 ( .A(n_357), .Y(n_1542) );
OAI211xp5_ASAP7_75t_L g1464 ( .A1(n_358), .A2(n_1406), .B(n_1465), .C(n_1467), .Y(n_1464) );
INVx1_ASAP7_75t_L g1502 ( .A(n_358), .Y(n_1502) );
INVx1_ASAP7_75t_L g1235 ( .A(n_361), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1936 ( .A(n_362), .Y(n_1936) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_363), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g984 ( .A(n_365), .Y(n_984) );
OAI211xp5_ASAP7_75t_SL g1275 ( .A1(n_366), .A2(n_516), .B(n_1276), .C(n_1284), .Y(n_1275) );
INVx1_ASAP7_75t_L g687 ( .A(n_368), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_369), .Y(n_1073) );
INVxp33_ASAP7_75t_SL g723 ( .A(n_372), .Y(n_723) );
INVx1_ASAP7_75t_L g2034 ( .A(n_374), .Y(n_2034) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_397), .B(n_1691), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1999 ( .A(n_379), .B(n_385), .Y(n_1999) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g2004 ( .A(n_380), .Y(n_2004) );
NAND2xp5_ASAP7_75t_L g2055 ( .A(n_380), .B(n_382), .Y(n_2055) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g2003 ( .A(n_382), .B(n_2004), .Y(n_2003) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_387), .B(n_469), .Y(n_1046) );
OR2x6_ASAP7_75t_L g1328 ( .A(n_387), .B(n_469), .Y(n_1328) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g511 ( .A(n_388), .B(n_396), .Y(n_511) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g623 ( .A(n_389), .B(n_624), .Y(n_623) );
INVx8_ASAP7_75t_L g1042 ( .A(n_390), .Y(n_1042) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_391), .Y(n_508) );
INVx1_ASAP7_75t_L g842 ( .A(n_391), .Y(n_842) );
INVx2_ASAP7_75t_SL g888 ( .A(n_391), .Y(n_888) );
OR2x2_ASAP7_75t_L g912 ( .A(n_391), .B(n_877), .Y(n_912) );
OR2x6_ASAP7_75t_L g1045 ( .A(n_391), .B(n_1035), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1681 ( .A(n_391), .Y(n_1681) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g482 ( .A(n_393), .B(n_394), .Y(n_482) );
INVx2_ASAP7_75t_L g495 ( .A(n_393), .Y(n_495) );
AND2x4_ASAP7_75t_L g499 ( .A(n_393), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_393), .Y(n_506) );
INVx1_ASAP7_75t_L g522 ( .A(n_393), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_394), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g500 ( .A(n_394), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_394), .Y(n_505) );
INVx1_ASAP7_75t_L g544 ( .A(n_394), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_394), .Y(n_553) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_395), .B(n_544), .Y(n_1030) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_396), .B(n_1032), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_396), .B(n_1032), .Y(n_1321) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_1241), .Y(n_397) );
XOR2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_753), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_672), .B1(n_673), .B2(n_751), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_403), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_593), .B2(n_594), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND4xp75_ASAP7_75t_SL g406 ( .A(n_407), .B(n_465), .C(n_483), .D(n_561), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_440), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_425), .B1(n_426), .B2(n_433), .C(n_434), .Y(n_408) );
INVx1_ASAP7_75t_L g707 ( .A(n_409), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_409), .A2(n_426), .B1(n_809), .B2(n_810), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_409), .A2(n_426), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g650 ( .A(n_410), .Y(n_650) );
INVx1_ASAP7_75t_L g1092 ( .A(n_410), .Y(n_1092) );
INVx2_ASAP7_75t_L g1210 ( .A(n_410), .Y(n_1210) );
HB1xp67_ASAP7_75t_L g2022 ( .A(n_410), .Y(n_2022) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_416), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g922 ( .A(n_412), .Y(n_922) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g983 ( .A(n_413), .Y(n_983) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g453 ( .A(n_414), .B(n_431), .Y(n_453) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g438 ( .A(n_415), .B(n_432), .Y(n_438) );
AND2x4_ASAP7_75t_L g458 ( .A(n_415), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OR2x6_ASAP7_75t_L g427 ( .A(n_417), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
OR2x2_ASAP7_75t_L g708 ( .A(n_417), .B(n_428), .Y(n_708) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_453), .Y(n_470) );
AND2x4_ASAP7_75t_L g921 ( .A(n_418), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g924 ( .A(n_418), .Y(n_924) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_418), .B(n_429), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1945 ( .A(n_418), .B(n_429), .Y(n_1945) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g592 ( .A(n_421), .B(n_566), .Y(n_592) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g565 ( .A(n_422), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g965 ( .A(n_422), .Y(n_965) );
INVx1_ASAP7_75t_L g970 ( .A(n_422), .Y(n_970) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_422), .Y(n_975) );
OR2x6_ASAP7_75t_L g908 ( .A(n_423), .B(n_529), .Y(n_908) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g447 ( .A(n_424), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g862 ( .A(n_424), .B(n_487), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_425), .A2(n_433), .B1(n_542), .B2(n_545), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_426), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_426), .A2(n_1072), .B1(n_1073), .B2(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g923 ( .A(n_428), .B(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x6_ASAP7_75t_L g985 ( .A(n_430), .B(n_970), .Y(n_985) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g444 ( .A(n_432), .B(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g680 ( .A(n_434), .Y(n_680) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_434), .Y(n_1185) );
NOR3xp33_ASAP7_75t_SL g1646 ( .A(n_434), .B(n_1647), .C(n_1665), .Y(n_1646) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g1123 ( .A(n_436), .Y(n_1123) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_437), .Y(n_948) );
AND2x4_ASAP7_75t_L g987 ( .A(n_437), .B(n_988), .Y(n_987) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_437), .Y(n_1015) );
INVx2_ASAP7_75t_L g1366 ( .A(n_437), .Y(n_1366) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_438), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_439), .B(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_449), .B1(n_450), .B2(n_454), .C(n_455), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_441), .A2(n_450), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_441), .A2(n_450), .B1(n_823), .B2(n_824), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_441), .A2(n_450), .B1(n_1066), .B2(n_1069), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_441), .A2(n_450), .B1(n_1255), .B2(n_1256), .Y(n_1254) );
AOI222xp33_ASAP7_75t_L g1543 ( .A1(n_441), .A2(n_450), .B1(n_468), .B2(n_1517), .C1(n_1524), .C2(n_1544), .Y(n_1543) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g1386 ( .A(n_443), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g1488 ( .A1(n_443), .A2(n_1489), .B1(n_1490), .B2(n_1491), .Y(n_1488) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_444), .Y(n_576) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_444), .Y(n_586) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_444), .Y(n_657) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_444), .Y(n_694) );
BUFx3_ASAP7_75t_L g705 ( .A(n_444), .Y(n_705) );
AND2x6_ASAP7_75t_L g968 ( .A(n_444), .B(n_969), .Y(n_968) );
BUFx2_ASAP7_75t_L g1264 ( .A(n_444), .Y(n_1264) );
BUFx2_ASAP7_75t_L g1574 ( .A(n_444), .Y(n_1574) );
INVx1_ASAP7_75t_L g464 ( .A(n_445), .Y(n_464) );
AND2x2_ASAP7_75t_L g450 ( .A(n_446), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g456 ( .A(n_447), .B(n_457), .Y(n_456) );
OR2x6_ASAP7_75t_L g460 ( .A(n_447), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g745 ( .A(n_447), .B(n_457), .Y(n_745) );
OR2x2_ASAP7_75t_L g747 ( .A(n_447), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g749 ( .A(n_447), .B(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g918 ( .A(n_448), .Y(n_918) );
OR2x2_ASAP7_75t_L g951 ( .A(n_448), .B(n_686), .Y(n_951) );
OR2x2_ASAP7_75t_L g953 ( .A(n_448), .B(n_954), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_449), .A2(n_533), .B1(n_536), .B2(n_540), .Y(n_532) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_451), .Y(n_1013) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g581 ( .A(n_452), .Y(n_581) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_L g570 ( .A(n_453), .Y(n_570) );
AND2x4_ASAP7_75t_L g973 ( .A(n_453), .B(n_974), .Y(n_973) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_453), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_454), .A2(n_508), .B1(n_524), .B2(n_525), .C(n_526), .Y(n_523) );
CKINVDCx6p67_ASAP7_75t_R g639 ( .A(n_456), .Y(n_639) );
INVx2_ASAP7_75t_L g945 ( .A(n_457), .Y(n_945) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_458), .Y(n_579) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_458), .Y(n_589) );
INVx1_ASAP7_75t_L g670 ( .A(n_458), .Y(n_670) );
INVx2_ASAP7_75t_L g954 ( .A(n_458), .Y(n_954) );
INVx1_ASAP7_75t_L g463 ( .A(n_459), .Y(n_463) );
CKINVDCx6p67_ASAP7_75t_R g641 ( .A(n_460), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_461), .A2(n_683), .B1(n_763), .B2(n_764), .C(n_765), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g1198 ( .A1(n_461), .A2(n_684), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
BUFx3_ASAP7_75t_L g1486 ( .A(n_461), .Y(n_1486) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx4f_ASAP7_75t_L g691 ( .A(n_462), .Y(n_691) );
INVx1_ASAP7_75t_L g1196 ( .A(n_462), .Y(n_1196) );
INVx1_ASAP7_75t_L g1484 ( .A(n_462), .Y(n_1484) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OR2x2_ASAP7_75t_L g686 ( .A(n_463), .B(n_464), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g643 ( .A(n_467), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_467), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_467), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_467), .B(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_467), .B(n_1088), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_467), .B(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_467), .B(n_1273), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_467), .B(n_1670), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g2023 ( .A(n_467), .B(n_2024), .Y(n_2023) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .Y(n_467) );
INVx2_ASAP7_75t_L g913 ( .A(n_468), .Y(n_913) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
AND2x4_ASAP7_75t_L g591 ( .A(n_469), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g1110 ( .A(n_469), .B(n_592), .Y(n_1110) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx2_ASAP7_75t_L g742 ( .A(n_472), .Y(n_742) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x6_ASAP7_75t_L g563 ( .A(n_473), .B(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g632 ( .A(n_473), .Y(n_632) );
AND2x4_ASAP7_75t_L g997 ( .A(n_473), .B(n_511), .Y(n_997) );
OAI31xp33_ASAP7_75t_L g1059 ( .A1(n_473), .A2(n_1060), .A3(n_1061), .B(n_1074), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_473), .B(n_564), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_473), .B(n_1370), .Y(n_1369) );
AND2x4_ASAP7_75t_L g1425 ( .A(n_473), .B(n_511), .Y(n_1425) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g560 ( .A(n_474), .Y(n_560) );
OR2x6_ASAP7_75t_L g884 ( .A(n_474), .B(n_623), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
AND2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g785 ( .A(n_476), .B(n_543), .Y(n_785) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g512 ( .A(n_477), .B(n_513), .Y(n_512) );
OR2x6_ASAP7_75t_L g546 ( .A(n_477), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g615 ( .A(n_477), .Y(n_615) );
OR2x2_ASAP7_75t_L g725 ( .A(n_477), .B(n_513), .Y(n_725) );
INVx1_ASAP7_75t_L g1529 ( .A(n_477), .Y(n_1529) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g737 ( .A(n_480), .Y(n_737) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g606 ( .A(n_481), .Y(n_606) );
INVx2_ASAP7_75t_L g1334 ( .A(n_481), .Y(n_1334) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_482), .Y(n_489) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_515), .A3(n_548), .B(n_558), .Y(n_483) );
CKINVDCx6p67_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_486), .A2(n_620), .B1(n_625), .B2(n_629), .C(n_630), .Y(n_619) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_487), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g530 ( .A(n_488), .Y(n_530) );
INVx1_ASAP7_75t_L g624 ( .A(n_488), .Y(n_624) );
BUFx6f_ASAP7_75t_L g1233 ( .A(n_489), .Y(n_1233) );
INVx3_ASAP7_75t_L g1283 ( .A(n_489), .Y(n_1283) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_496), .B1(n_497), .B2(n_501), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_491), .A2(n_1469), .B1(n_1496), .B2(n_1498), .Y(n_1495) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g846 ( .A(n_492), .Y(n_846) );
INVx2_ASAP7_75t_L g1173 ( .A(n_492), .Y(n_1173) );
INVx2_ASAP7_75t_L g1675 ( .A(n_492), .Y(n_1675) );
BUFx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g730 ( .A(n_493), .Y(n_730) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
BUFx2_ASAP7_75t_L g896 ( .A(n_494), .Y(n_896) );
INVx1_ASAP7_75t_L g547 ( .A(n_495), .Y(n_547) );
AND2x4_ASAP7_75t_L g551 ( .A(n_495), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g602 ( .A(n_498), .Y(n_602) );
INVx4_ASAP7_75t_L g628 ( .A(n_498), .Y(n_628) );
BUFx3_ASAP7_75t_L g849 ( .A(n_498), .Y(n_849) );
INVx2_ASAP7_75t_SL g898 ( .A(n_498), .Y(n_898) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g539 ( .A(n_499), .Y(n_539) );
INVx1_ASAP7_75t_L g557 ( .A(n_499), .Y(n_557) );
INVx1_ASAP7_75t_L g1039 ( .A(n_499), .Y(n_1039) );
AND2x4_ASAP7_75t_L g521 ( .A(n_500), .B(n_522), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_507), .B1(n_508), .B2(n_509), .C(n_510), .Y(n_502) );
INVx2_ASAP7_75t_L g1064 ( .A(n_503), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1178 ( .A(n_503), .Y(n_1178) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_503), .A2(n_508), .B1(n_719), .B2(n_1194), .C(n_1197), .Y(n_1223) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g514 ( .A(n_505), .B(n_506), .Y(n_514) );
INVx1_ASAP7_75t_L g1032 ( .A(n_506), .Y(n_1032) );
INVx1_ASAP7_75t_L g718 ( .A(n_508), .Y(n_718) );
BUFx2_ASAP7_75t_L g790 ( .A(n_508), .Y(n_790) );
INVx1_ASAP7_75t_L g1085 ( .A(n_508), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_508), .A2(n_1081), .B1(n_1480), .B2(n_1482), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_508), .A2(n_1500), .B1(n_1501), .B2(n_1502), .Y(n_1499) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_510), .A2(n_763), .B1(n_764), .B2(n_789), .C(n_790), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_510), .A2(n_839), .B1(n_840), .B2(n_841), .C(n_843), .Y(n_838) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g720 ( .A(n_511), .Y(n_720) );
INVx2_ASAP7_75t_L g630 ( .A(n_512), .Y(n_630) );
INVx1_ASAP7_75t_L g1082 ( .A(n_513), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_513), .B(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g524 ( .A(n_514), .Y(n_524) );
BUFx2_ASAP7_75t_L g716 ( .A(n_514), .Y(n_716) );
INVx2_ASAP7_75t_L g1419 ( .A(n_514), .Y(n_1419) );
INVx8_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_517), .A2(n_599), .B1(n_603), .B2(n_610), .C(n_611), .Y(n_598) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g555 ( .A(n_518), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1024 ( .A(n_520), .Y(n_1024) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_521), .Y(n_609) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_521), .Y(n_781) );
BUFx3_ASAP7_75t_L g865 ( .A(n_521), .Y(n_865) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_521), .B(n_1026), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1618 ( .A(n_521), .Y(n_1618) );
BUFx2_ASAP7_75t_L g839 ( .A(n_524), .Y(n_839) );
INVx1_ASAP7_75t_L g891 ( .A(n_524), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g1513 ( .A1(n_524), .A2(n_1514), .B(n_1515), .Y(n_1513) );
OAI221xp5_ASAP7_75t_L g1678 ( .A1(n_524), .A2(n_719), .B1(n_1653), .B2(n_1656), .C(n_1679), .Y(n_1678) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_526), .A2(n_717), .B1(n_1063), .B2(n_1065), .C(n_1066), .Y(n_1062) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g782 ( .A(n_528), .Y(n_782) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g1522 ( .A(n_529), .Y(n_1522) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g1027 ( .A(n_530), .Y(n_1027) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g1277 ( .A(n_534), .Y(n_1277) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g722 ( .A(n_535), .Y(n_722) );
INVx1_ASAP7_75t_L g794 ( .A(n_535), .Y(n_794) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_535), .Y(n_1218) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g1002 ( .A(n_538), .Y(n_1002) );
INVx2_ASAP7_75t_L g1078 ( .A(n_538), .Y(n_1078) );
INVx2_ASAP7_75t_L g1230 ( .A(n_538), .Y(n_1230) );
INVx2_ASAP7_75t_SL g1497 ( .A(n_538), .Y(n_1497) );
INVx2_ASAP7_75t_L g1628 ( .A(n_538), .Y(n_1628) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g798 ( .A(n_539), .Y(n_798) );
INVx3_ASAP7_75t_L g1222 ( .A(n_539), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_542), .A2(n_545), .B1(n_740), .B2(n_741), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_542), .A2(n_545), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_542), .A2(n_545), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_542), .A2(n_545), .B1(n_1259), .B2(n_1260), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g2041 ( .A1(n_542), .A2(n_545), .B1(n_2042), .B2(n_2043), .Y(n_2041) );
AND2x4_ASAP7_75t_L g1991 ( .A(n_543), .B(n_876), .Y(n_1991) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g614 ( .A(n_544), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g1526 ( .A1(n_544), .A2(n_880), .B1(n_1527), .B2(n_1528), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_545), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_545), .A2(n_785), .B1(n_809), .B2(n_810), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1687 ( .A1(n_545), .A2(n_785), .B1(n_1688), .B2(n_1689), .Y(n_1687) );
CKINVDCx11_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g880 ( .A(n_547), .Y(n_880) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_550), .A2(n_555), .B1(n_617), .B2(n_618), .Y(n_616) );
INVx3_ASAP7_75t_L g711 ( .A(n_550), .Y(n_711) );
BUFx2_ASAP7_75t_L g600 ( .A(n_551), .Y(n_600) );
BUFx2_ASAP7_75t_L g626 ( .A(n_551), .Y(n_626) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_551), .Y(n_871) );
BUFx6f_ASAP7_75t_L g1000 ( .A(n_551), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_551), .B(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1374 ( .A(n_551), .Y(n_1374) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g712 ( .A(n_555), .Y(n_712) );
INVx1_ASAP7_75t_L g734 ( .A(n_556), .Y(n_734) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g834 ( .A(n_557), .Y(n_834) );
OAI31xp33_ASAP7_75t_L g827 ( .A1(n_558), .A2(n_828), .A3(n_837), .B(n_850), .Y(n_827) );
INVx5_ASAP7_75t_L g1968 ( .A(n_558), .Y(n_1968) );
BUFx8_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g1119 ( .A(n_559), .Y(n_1119) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g956 ( .A(n_560), .Y(n_956) );
AND2x4_ASAP7_75t_L g991 ( .A(n_560), .B(n_992), .Y(n_991) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_560), .B(n_992), .Y(n_1414) );
AOI33xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_567), .A3(n_573), .B1(n_580), .B2(n_583), .B3(n_590), .Y(n_561) );
AOI33xp33_ASAP7_75t_L g1093 ( .A1(n_562), .A2(n_1094), .A3(n_1099), .B1(n_1102), .B2(n_1105), .B3(n_1108), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_563), .Y(n_654) );
OAI22xp5_ASAP7_75t_SL g681 ( .A1(n_563), .A2(n_682), .B1(n_696), .B2(n_697), .Y(n_681) );
OAI22xp5_ASAP7_75t_SL g761 ( .A1(n_563), .A2(n_696), .B1(n_762), .B2(n_766), .Y(n_761) );
INVx2_ASAP7_75t_L g1262 ( .A(n_563), .Y(n_1262) );
OAI22xp5_ASAP7_75t_SL g2011 ( .A1(n_563), .A2(n_1207), .B1(n_2012), .B2(n_2016), .Y(n_2011) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_SL g940 ( .A(n_565), .Y(n_940) );
INVx1_ASAP7_75t_L g1370 ( .A(n_565), .Y(n_1370) );
BUFx3_ASAP7_75t_L g1960 ( .A(n_565), .Y(n_1960) );
INVx1_ASAP7_75t_L g992 ( .A(n_566), .Y(n_992) );
BUFx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g1434 ( .A(n_569), .Y(n_1434) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g662 ( .A(n_570), .Y(n_662) );
INVx2_ASAP7_75t_L g944 ( .A(n_570), .Y(n_944) );
INVx2_ASAP7_75t_L g966 ( .A(n_570), .Y(n_966) );
BUFx6f_ASAP7_75t_L g1104 ( .A(n_570), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_570), .Y(n_1535) );
INVx1_ASAP7_75t_L g1635 ( .A(n_570), .Y(n_1635) );
AOI222xp33_ASAP7_75t_L g1307 ( .A1(n_571), .A2(n_985), .B1(n_1308), .B2(n_1309), .C1(n_1310), .C2(n_1312), .Y(n_1307) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g582 ( .A(n_572), .Y(n_582) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_572), .Y(n_648) );
INVx2_ASAP7_75t_SL g664 ( .A(n_572), .Y(n_664) );
AND2x4_ASAP7_75t_L g936 ( .A(n_572), .B(n_918), .Y(n_936) );
INVx1_ASAP7_75t_L g939 ( .A(n_572), .Y(n_939) );
INVx1_ASAP7_75t_L g1578 ( .A(n_572), .Y(n_1578) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g813 ( .A(n_575), .Y(n_813) );
INVx1_ASAP7_75t_L g1127 ( .A(n_575), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1536 ( .A1(n_575), .A2(n_670), .B1(n_1510), .B2(n_1512), .Y(n_1536) );
OAI22xp5_ASAP7_75t_L g1660 ( .A1(n_575), .A2(n_1661), .B1(n_1662), .B2(n_1664), .Y(n_1660) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
BUFx3_ASAP7_75t_L g668 ( .A(n_576), .Y(n_668) );
AND2x4_ASAP7_75t_L g917 ( .A(n_576), .B(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
INVx1_ASAP7_75t_L g927 ( .A(n_579), .Y(n_927) );
BUFx3_ASAP7_75t_L g1142 ( .A(n_579), .Y(n_1142) );
AOI222xp33_ASAP7_75t_L g978 ( .A1(n_582), .A2(n_979), .B1(n_980), .B2(n_981), .C1(n_984), .C2(n_985), .Y(n_978) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g1106 ( .A(n_585), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1538 ( .A1(n_585), .A2(n_1097), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g1467 ( .A1(n_586), .A2(n_985), .A3(n_1456), .B1(n_1460), .B2(n_1468), .C1(n_1469), .C2(n_1470), .Y(n_1467) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g814 ( .A(n_588), .Y(n_814) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x6_ASAP7_75t_L g977 ( .A(n_589), .B(n_964), .Y(n_977) );
INVx1_ASAP7_75t_L g1011 ( .A(n_589), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_589), .Y(n_1107) );
INVx1_ASAP7_75t_L g1491 ( .A(n_589), .Y(n_1491) );
BUFx6f_ASAP7_75t_L g1580 ( .A(n_589), .Y(n_1580) );
BUFx6f_ASAP7_75t_L g1663 ( .A(n_589), .Y(n_1663) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_590), .Y(n_696) );
BUFx4f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx4f_ASAP7_75t_L g671 ( .A(n_591), .Y(n_671) );
AOI33xp33_ASAP7_75t_L g1008 ( .A1(n_591), .A2(n_654), .A3(n_1009), .B1(n_1012), .B2(n_1016), .B3(n_1019), .Y(n_1008) );
INVx4_ASAP7_75t_L g1207 ( .A(n_591), .Y(n_1207) );
AOI33xp33_ASAP7_75t_L g1430 ( .A1(n_591), .A2(n_654), .A3(n_1431), .B1(n_1432), .B2(n_1433), .B3(n_1436), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1532 ( .A1(n_591), .A2(n_1262), .B1(n_1533), .B2(n_1537), .C(n_1541), .Y(n_1532) );
INVx2_ASAP7_75t_L g932 ( .A(n_592), .Y(n_932) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NOR4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_633), .C(n_642), .D(n_644), .Y(n_596) );
AOI31xp33_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_616), .A3(n_619), .B(n_631), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_602), .A2(n_895), .B1(n_900), .B2(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g621 ( .A(n_606), .Y(n_621) );
AND2x4_ASAP7_75t_L g868 ( .A(n_606), .B(n_862), .Y(n_868) );
BUFx3_ASAP7_75t_L g1004 ( .A(n_606), .Y(n_1004) );
AOI211xp5_ASAP7_75t_L g1388 ( .A1(n_607), .A2(n_1025), .B(n_1389), .C(n_1390), .Y(n_1388) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g622 ( .A(n_608), .Y(n_622) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_609), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2x1_ASAP7_75t_SL g875 ( .A(n_613), .B(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g1558 ( .A1(n_622), .A2(n_1457), .B1(n_1559), .B2(n_1560), .C1(n_1561), .C2(n_1562), .Y(n_1558) );
INVx1_ASAP7_75t_L g1035 ( .A(n_624), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1985 ( .A(n_626), .Y(n_1985) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_628), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_628), .A2(n_1130), .B1(n_1147), .B2(n_1171), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1683 ( .A1(n_628), .A2(n_846), .B1(n_1684), .B2(n_1685), .C(n_1686), .Y(n_1683) );
INVx2_ASAP7_75t_L g1983 ( .A(n_628), .Y(n_1983) );
INVx2_ASAP7_75t_L g1294 ( .A(n_631), .Y(n_1294) );
CKINVDCx8_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g773 ( .A1(n_632), .A2(n_774), .A3(n_787), .B(n_800), .Y(n_773) );
OAI31xp33_ASAP7_75t_SL g2025 ( .A1(n_632), .A2(n_2026), .A3(n_2027), .B(n_2036), .Y(n_2025) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_639), .A2(n_641), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_639), .A2(n_641), .B1(n_1065), .B2(n_1070), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_639), .A2(n_641), .B1(n_1252), .B2(n_1253), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_639), .A2(n_641), .B1(n_1518), .B2(n_1520), .Y(n_1545) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_649), .C(n_653), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g1090 ( .A(n_645), .B(n_1091), .C(n_1093), .Y(n_1090) );
NAND3xp33_ASAP7_75t_L g1257 ( .A(n_645), .B(n_1258), .C(n_1261), .Y(n_1257) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g807 ( .A(n_647), .B(n_808), .C(n_811), .Y(n_807) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_648), .Y(n_666) );
INVx1_ASAP7_75t_L g1018 ( .A(n_648), .Y(n_1018) );
AOI33xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .A3(n_659), .B1(n_665), .B2(n_667), .B3(n_671), .Y(n_653) );
AOI33xp33_ASAP7_75t_L g811 ( .A1(n_654), .A2(n_671), .A3(n_812), .B1(n_815), .B2(n_816), .B3(n_817), .Y(n_811) );
AOI33xp33_ASAP7_75t_L g1342 ( .A1(n_654), .A2(n_671), .A3(n_1343), .B1(n_1344), .B2(n_1345), .B3(n_1346), .Y(n_1342) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx3_ASAP7_75t_L g770 ( .A(n_657), .Y(n_770) );
INVx1_ASAP7_75t_L g1202 ( .A(n_657), .Y(n_1202) );
INVx1_ASAP7_75t_L g1649 ( .A(n_657), .Y(n_1649) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_663), .B(n_1402), .Y(n_1401) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1101 ( .A(n_664), .Y(n_1101) );
INVx1_ASAP7_75t_L g1268 ( .A(n_664), .Y(n_1268) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g695 ( .A(n_670), .Y(n_695) );
INVx1_ASAP7_75t_L g1205 ( .A(n_670), .Y(n_1205) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AND4x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .C(n_709), .D(n_743), .Y(n_676) );
NOR3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_681), .C(n_706), .Y(n_679) );
NOR3xp33_ASAP7_75t_SL g759 ( .A(n_680), .B(n_760), .C(n_761), .Y(n_759) );
NOR3xp33_ASAP7_75t_SL g2010 ( .A(n_680), .B(n_2011), .C(n_2021), .Y(n_2010) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_688), .B2(n_689), .C(n_692), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g2012 ( .A1(n_683), .A2(n_689), .B1(n_2013), .B2(n_2014), .C(n_2015), .Y(n_2012) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g699 ( .A(n_686), .Y(n_699) );
BUFx2_ASAP7_75t_L g930 ( .A(n_686), .Y(n_930) );
OR2x2_ASAP7_75t_L g1411 ( .A(n_686), .B(n_1412), .Y(n_1411) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_687), .A2(n_688), .B1(n_715), .B2(n_717), .C(n_719), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_689), .A2(n_698), .B1(n_767), .B2(n_768), .C(n_769), .Y(n_766) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g701 ( .A(n_691), .Y(n_701) );
INVx1_ASAP7_75t_L g929 ( .A(n_691), .Y(n_929) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g750 ( .A(n_694), .Y(n_750) );
BUFx4f_ASAP7_75t_L g1095 ( .A(n_694), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_701), .B2(n_702), .C(n_703), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g2016 ( .A1(n_698), .A2(n_1654), .B1(n_2017), .B2(n_2018), .C(n_2019), .Y(n_2016) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g748 ( .A(n_699), .Y(n_748) );
INVx2_ASAP7_75t_L g1481 ( .A(n_699), .Y(n_1481) );
HB1xp67_ASAP7_75t_L g1949 ( .A(n_699), .Y(n_1949) );
OAI22xp33_ASAP7_75t_L g1657 ( .A1(n_701), .A2(n_1481), .B1(n_1658), .B2(n_1659), .Y(n_1657) );
BUFx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_705), .Y(n_1189) );
OAI31xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .A3(n_726), .B(n_742), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g789 ( .A(n_716), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g1286 ( .A1(n_717), .A2(n_719), .B1(n_789), .B2(n_1287), .C(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_719), .A2(n_1081), .B1(n_1083), .B2(n_1084), .C(n_1086), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g2035 ( .A1(n_719), .A2(n_790), .B1(n_1419), .B2(n_2013), .C(n_2014), .Y(n_2035) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_722), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_722), .A2(n_1290), .B1(n_1291), .B2(n_1292), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_722), .A2(n_1510), .B1(n_1511), .B2(n_1512), .Y(n_1509) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_722), .A2(n_1376), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_731), .B1(n_732), .B2(n_735), .C(n_736), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g2037 ( .A1(n_728), .A2(n_831), .B1(n_2038), .B2(n_2039), .C(n_2040), .Y(n_2037) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g776 ( .A(n_729), .Y(n_776) );
INVx2_ASAP7_75t_L g2029 ( .A(n_729), .Y(n_2029) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g830 ( .A(n_730), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_732), .A2(n_776), .B1(n_777), .B2(n_778), .C(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1279 ( .A(n_734), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1494 ( .A1(n_734), .A2(n_1226), .B1(n_1474), .B2(n_1476), .Y(n_1494) );
OAI31xp33_ASAP7_75t_L g1213 ( .A1(n_742), .A2(n_1214), .A3(n_1215), .B(n_1224), .Y(n_1213) );
OAI31xp33_ASAP7_75t_L g1507 ( .A1(n_742), .A2(n_1508), .A3(n_1530), .B(n_1531), .Y(n_1507) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AO22x2_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_1052), .B1(n_1053), .B2(n_1240), .Y(n_753) );
INVx2_ASAP7_75t_SL g1240 ( .A(n_754), .Y(n_1240) );
AO22x2_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_853), .B2(n_1051), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AO22x1_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_804), .B1(n_851), .B2(n_852), .Y(n_756) );
INVx1_ASAP7_75t_L g852 ( .A(n_757), .Y(n_852) );
AND4x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_771), .C(n_773), .D(n_801), .Y(n_758) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_SL g1317 ( .A(n_781), .Y(n_1317) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_781), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_795), .B1(n_796), .B2(n_799), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
BUFx3_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g861 ( .A(n_798), .B(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g851 ( .A(n_804), .Y(n_851) );
AND3x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_825), .C(n_827), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_818), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_820), .A2(n_824), .B1(n_830), .B2(n_831), .C(n_835), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_830), .A2(n_1076), .B1(n_1077), .B2(n_1079), .Y(n_1075) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g1166 ( .A(n_842), .Y(n_1166) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1051 ( .A(n_853), .Y(n_1051) );
AOI22x1_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_957), .B1(n_1048), .B2(n_1049), .Y(n_853) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_909), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_872), .C(n_883), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_866), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_863), .B2(n_864), .Y(n_858) );
BUFx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_861), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1977 ( .A(n_861), .Y(n_1977) );
AND2x6_ASAP7_75t_L g864 ( .A(n_862), .B(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g870 ( .A(n_862), .B(n_871), .Y(n_870) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_862), .B(n_871), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1974 ( .A(n_862), .B(n_871), .Y(n_1974) );
OAI221xp5_ASAP7_75t_L g928 ( .A1(n_863), .A2(n_867), .B1(n_929), .B2(n_930), .C(n_931), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_864), .A2(n_1153), .B1(n_1154), .B2(n_1155), .Y(n_1152) );
BUFx2_ASAP7_75t_L g1979 ( .A(n_864), .Y(n_1979) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_865), .B(n_876), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_868), .A2(n_1157), .B1(n_1158), .B2(n_1159), .Y(n_1156) );
BUFx2_ASAP7_75t_L g1972 ( .A(n_868), .Y(n_1972) );
INVx2_ASAP7_75t_SL g1338 ( .A(n_871), .Y(n_1338) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_874), .Y(n_1161) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND2x1p5_ASAP7_75t_L g879 ( .A(n_876), .B(n_880), .Y(n_879) );
AND2x4_ASAP7_75t_L g1993 ( .A(n_876), .B(n_1458), .Y(n_1993) );
AND2x4_ASAP7_75t_L g1995 ( .A(n_876), .B(n_1618), .Y(n_1995) );
INVx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
BUFx4f_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
OAI33xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .A3(n_893), .B1(n_899), .B2(n_902), .B3(n_906), .Y(n_883) );
INVx1_ASAP7_75t_L g1164 ( .A(n_884), .Y(n_1164) );
OAI33xp33_ASAP7_75t_L g1492 ( .A1(n_884), .A2(n_906), .A3(n_1493), .B1(n_1494), .B2(n_1495), .B3(n_1499), .Y(n_1492) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_889), .B1(n_890), .B2(n_892), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_886), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1177 ( .A1(n_886), .A2(n_1144), .B1(n_1146), .B2(n_1178), .Y(n_1177) );
BUFx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g904 ( .A(n_891), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_897), .B2(n_898), .Y(n_893) );
BUFx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g1227 ( .A(n_896), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_896), .B(n_1449), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_898), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_898), .A2(n_1171), .B1(n_1174), .B2(n_1175), .Y(n_1170) );
AOI211xp5_ASAP7_75t_L g916 ( .A1(n_900), .A2(n_917), .B(n_919), .C(n_925), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_901), .A2(n_903), .B1(n_950), .B2(n_952), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_905), .A2(n_934), .B1(n_937), .B2(n_941), .C(n_946), .Y(n_933) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AOI33xp33_ASAP7_75t_L g1330 ( .A1(n_907), .A2(n_1331), .A3(n_1332), .B1(n_1335), .B2(n_1336), .B3(n_1339), .Y(n_1330) );
AOI33xp33_ASAP7_75t_L g1424 ( .A1(n_907), .A2(n_1425), .A3(n_1426), .B1(n_1427), .B2(n_1428), .B3(n_1429), .Y(n_1424) );
AOI33xp33_ASAP7_75t_L g1564 ( .A1(n_907), .A2(n_1425), .A3(n_1565), .B1(n_1566), .B2(n_1568), .B3(n_1570), .Y(n_1564) );
INVx6_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx5_ASAP7_75t_L g1007 ( .A(n_908), .Y(n_1007) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_914), .B(n_915), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx5_ASAP7_75t_L g1149 ( .A(n_911), .Y(n_1149) );
INVx1_ASAP7_75t_L g1935 ( .A(n_911), .Y(n_1935) );
AND2x4_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
AOI31xp33_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_933), .A3(n_949), .B(n_955), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_917), .A2(n_1122), .B1(n_1126), .B2(n_1130), .C(n_1131), .Y(n_1121) );
INVx1_ASAP7_75t_L g1941 ( .A(n_917), .Y(n_1941) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g1132 ( .A(n_921), .Y(n_1132) );
INVx1_ASAP7_75t_L g1943 ( .A(n_921), .Y(n_1943) );
INVx1_ASAP7_75t_SL g947 ( .A(n_924), .Y(n_947) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g1648 ( .A1(n_927), .A2(n_1649), .B1(n_1650), .B2(n_1651), .Y(n_1648) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_930), .A2(n_1194), .B1(n_1195), .B2(n_1197), .Y(n_1193) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_932), .Y(n_1125) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
BUFx6f_ASAP7_75t_L g1143 ( .A(n_936), .Y(n_1143) );
INVx1_ASAP7_75t_L g1955 ( .A(n_936), .Y(n_1955) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1140 ( .A(n_940), .Y(n_1140) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_944), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1135 ( .A1(n_946), .A2(n_1136), .B1(n_1141), .B2(n_1143), .C(n_1144), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1963 ( .A(n_946), .Y(n_1963) );
AND2x4_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
INVx1_ASAP7_75t_L g1138 ( .A(n_948), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g1435 ( .A(n_948), .Y(n_1435) );
OAI21xp33_ASAP7_75t_L g1606 ( .A1(n_948), .A2(n_988), .B(n_1607), .Y(n_1606) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_950), .A2(n_952), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1964 ( .A1(n_950), .A2(n_952), .B1(n_1965), .B2(n_1966), .Y(n_1964) );
INVx6_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx4_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g1098 ( .A(n_954), .Y(n_1098) );
INVx1_ASAP7_75t_L g1478 ( .A(n_954), .Y(n_1478) );
INVx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_L g1048 ( .A(n_957), .Y(n_1048) );
INVx1_ASAP7_75t_L g1047 ( .A(n_959), .Y(n_1047) );
AOI211x1_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_989), .B(n_993), .C(n_1020), .Y(n_959) );
NAND4xp25_ASAP7_75t_L g960 ( .A(n_961), .B(n_971), .C(n_978), .D(n_986), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_963), .B1(n_967), .B2(n_968), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_963), .A2(n_973), .B1(n_1557), .B2(n_1589), .Y(n_1588) );
AND2x4_ASAP7_75t_L g963 ( .A(n_964), .B(n_966), .Y(n_963) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_964), .B(n_966), .Y(n_1302) );
INVx1_ASAP7_75t_SL g964 ( .A(n_965), .Y(n_964) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_965), .B(n_1587), .Y(n_1586) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_968), .A2(n_1301), .B1(n_1302), .B2(n_1303), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_968), .A2(n_977), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
CKINVDCx6p67_ASAP7_75t_R g1408 ( .A(n_968), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_968), .A2(n_977), .B1(n_1591), .B2(n_1592), .Y(n_1590) );
AOI221xp5_ASAP7_75t_L g1601 ( .A1(n_968), .A2(n_973), .B1(n_1602), .B2(n_1603), .C(n_1604), .Y(n_1601) );
INVx1_ASAP7_75t_L g988 ( .A(n_969), .Y(n_988) );
INVx1_ASAP7_75t_L g1412 ( .A(n_969), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_969), .B(n_1015), .Y(n_1466) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B1(n_976), .B2(n_977), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_972), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_973), .A2(n_977), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_973), .A2(n_1302), .B1(n_1357), .B2(n_1358), .Y(n_1356) );
INVx4_ASAP7_75t_L g1413 ( .A(n_973), .Y(n_1413) );
AND2x4_ASAP7_75t_L g981 ( .A(n_974), .B(n_982), .Y(n_981) );
AND2x2_ASAP7_75t_SL g1470 ( .A(n_974), .B(n_982), .Y(n_1470) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx4_ASAP7_75t_L g1409 ( .A(n_977), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_977), .A2(n_1302), .B1(n_1599), .B2(n_1600), .Y(n_1598) );
INVx1_ASAP7_75t_L g1311 ( .A(n_981), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_981), .A2(n_985), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g1587 ( .A(n_983), .Y(n_1587) );
INVx3_ASAP7_75t_L g1355 ( .A(n_985), .Y(n_1355) );
NAND4xp25_ASAP7_75t_SL g1299 ( .A(n_986), .B(n_1300), .C(n_1304), .D(n_1307), .Y(n_1299) );
INVx5_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
AOI211xp5_ASAP7_75t_L g1351 ( .A1(n_987), .A2(n_1352), .B(n_1353), .C(n_1354), .Y(n_1351) );
CKINVDCx8_ASAP7_75t_R g1406 ( .A(n_987), .Y(n_1406) );
AOI211xp5_ASAP7_75t_L g1582 ( .A1(n_987), .A2(n_1466), .B(n_1583), .C(n_1584), .Y(n_1582) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx6f_ASAP7_75t_L g1313 ( .A(n_991), .Y(n_1313) );
AO211x2_ASAP7_75t_L g1349 ( .A1(n_991), .A2(n_1350), .B(n_1362), .C(n_1387), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_1008), .Y(n_993) );
AOI33xp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_998), .A3(n_1003), .B1(n_1005), .B2(n_1006), .B3(n_1007), .Y(n_994) );
AOI33xp33_ASAP7_75t_L g1981 ( .A1(n_995), .A2(n_1982), .A3(n_1984), .B1(n_1987), .B2(n_1988), .B3(n_1989), .Y(n_1981) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_997), .Y(n_1331) );
NAND3xp33_ASAP7_75t_L g1378 ( .A(n_997), .B(n_1379), .C(n_1380), .Y(n_1378) );
BUFx3_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
CKINVDCx8_ASAP7_75t_R g1179 ( .A(n_1007), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1371 ( .A(n_1007), .B(n_1372), .C(n_1377), .Y(n_1371) );
NAND3xp33_ASAP7_75t_L g1626 ( .A(n_1007), .B(n_1627), .C(n_1629), .Y(n_1626) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_1015), .Y(n_1353) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
AOI31xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1033), .A3(n_1041), .B(n_1046), .Y(n_1020) );
AOI211xp5_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1023), .B(n_1025), .C(n_1028), .Y(n_1021) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1024), .Y(n_1281) );
AOI211xp5_ASAP7_75t_L g1315 ( .A1(n_1025), .A2(n_1316), .B(n_1318), .C(n_1319), .Y(n_1315) );
NOR3xp33_ASAP7_75t_L g1416 ( .A(n_1025), .B(n_1417), .C(n_1420), .Y(n_1416) );
CKINVDCx11_ASAP7_75t_R g1452 ( .A(n_1025), .Y(n_1452) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVxp67_ASAP7_75t_L g1459 ( .A(n_1027), .Y(n_1459) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1029), .Y(n_1561) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx2_ASAP7_75t_L g1320 ( .A(n_1030), .Y(n_1320) );
INVx2_ASAP7_75t_L g1418 ( .A(n_1030), .Y(n_1418) );
AOI322xp5_ASAP7_75t_L g1453 ( .A1(n_1030), .A2(n_1449), .A3(n_1454), .B1(n_1455), .B2(n_1456), .C1(n_1457), .C2(n_1460), .Y(n_1453) );
AOI222xp33_ASAP7_75t_L g1612 ( .A1(n_1030), .A2(n_1457), .B1(n_1613), .B2(n_1614), .C1(n_1615), .C2(n_1616), .Y(n_1612) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1032), .Y(n_1458) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_1034), .A2(n_1036), .B1(n_1037), .B2(n_1040), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_1034), .A2(n_1037), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
AOI22xp33_ASAP7_75t_SL g1391 ( .A1(n_1034), .A2(n_1392), .B1(n_1393), .B2(n_1394), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_1034), .A2(n_1393), .B1(n_1422), .B2(n_1423), .Y(n_1421) );
AOI22xp5_ASAP7_75t_L g1552 ( .A1(n_1034), .A2(n_1037), .B1(n_1553), .B2(n_1554), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g1609 ( .A1(n_1034), .A2(n_1037), .B1(n_1610), .B2(n_1611), .Y(n_1609) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_1035), .B(n_1038), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1393 ( .A(n_1035), .B(n_1038), .Y(n_1393) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1035), .Y(n_1449) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g1292 ( .A(n_1039), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_1042), .A2(n_1305), .B1(n_1326), .B2(n_1327), .Y(n_1325) );
AOI22xp33_ASAP7_75t_SL g1395 ( .A1(n_1042), .A2(n_1044), .B1(n_1358), .B2(n_1396), .Y(n_1395) );
AOI211xp5_ASAP7_75t_L g1445 ( .A1(n_1042), .A2(n_1446), .B(n_1447), .C(n_1451), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_1042), .A2(n_1327), .B1(n_1556), .B2(n_1557), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_1042), .A2(n_1327), .B1(n_1602), .B2(n_1620), .Y(n_1619) );
INVx5_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx4_ASAP7_75t_L g1327 ( .A(n_1045), .Y(n_1327) );
OAI211xp5_ASAP7_75t_L g1444 ( .A1(n_1046), .A2(n_1445), .B(n_1461), .C(n_1471), .Y(n_1444) );
INVx3_ASAP7_75t_SL g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
XOR2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1180), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
AOI22x1_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1057), .B1(n_1114), .B2(n_1115), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
NAND3xp33_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1087), .C(n_1089), .Y(n_1058) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1064), .Y(n_1168) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1064), .Y(n_1501) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NOR2xp33_ASAP7_75t_SL g1089 ( .A(n_1090), .B(n_1111), .Y(n_1089) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1096), .Y(n_1191) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1097), .Y(n_1265) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1097), .Y(n_1271) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_1098), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1962 ( .A(n_1100), .Y(n_1962) );
INVx4_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1104), .Y(n_1124) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1104), .Y(n_1384) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1106), .Y(n_1475) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AOI33xp33_ASAP7_75t_L g1261 ( .A1(n_1110), .A2(n_1262), .A3(n_1263), .B1(n_1266), .B2(n_1269), .B3(n_1270), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_1110), .B(n_1383), .C(n_1385), .Y(n_1382) );
AOI33xp33_ASAP7_75t_L g1571 ( .A1(n_1110), .A2(n_1572), .A3(n_1573), .B1(n_1575), .B2(n_1576), .B3(n_1579), .Y(n_1571) );
NAND3xp33_ASAP7_75t_L g1633 ( .A(n_1110), .B(n_1634), .C(n_1636), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
XNOR2x1_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1150), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1120), .B1(n_1148), .B2(n_1149), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1135), .C(n_1145), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NOR3xp33_ASAP7_75t_SL g1150 ( .A(n_1151), .B(n_1160), .C(n_1162), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1156), .Y(n_1151) );
OAI33xp33_ASAP7_75t_L g1162 ( .A1(n_1163), .A2(n_1165), .A3(n_1170), .B1(n_1176), .B2(n_1177), .B3(n_1179), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1167), .B1(n_1168), .B2(n_1169), .Y(n_1165) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1989 ( .A(n_1179), .Y(n_1989) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
AND4x1_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1211), .C(n_1213), .D(n_1237), .Y(n_1183) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .C(n_1208), .Y(n_1184) );
OAI33xp33_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1188), .A3(n_1193), .B1(n_1198), .B2(n_1201), .B3(n_1207), .Y(n_1186) );
OAI33xp33_ASAP7_75t_L g1472 ( .A1(n_1187), .A2(n_1207), .A3(n_1473), .B1(n_1479), .B2(n_1485), .B3(n_1488), .Y(n_1472) );
INVx1_ASAP7_75t_SL g1572 ( .A(n_1187), .Y(n_1572) );
OAI33xp33_ASAP7_75t_L g1647 ( .A1(n_1187), .A2(n_1207), .A3(n_1648), .B1(n_1652), .B2(n_1657), .B3(n_1660), .Y(n_1647) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1190), .A2(n_1192), .B1(n_1217), .B2(n_1219), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_1202), .A2(n_1203), .B1(n_1204), .B2(n_1206), .Y(n_1201) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1222), .Y(n_1376) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1222), .Y(n_1511) );
INVx1_ASAP7_75t_L g2033 ( .A(n_1222), .Y(n_2033) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1228), .B1(n_1229), .B2(n_1231), .C(n_1232), .Y(n_1225) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1233), .Y(n_1341) );
A2O1A1Ixp33_ASAP7_75t_L g1523 ( .A1(n_1233), .A2(n_1524), .B(n_1525), .C(n_1529), .Y(n_1523) );
NOR2xp33_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1243), .B1(n_1641), .B2(n_1690), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
AO22x2_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1439), .B1(n_1440), .B2(n_1640), .Y(n_1243) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1244), .Y(n_1640) );
XOR2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1295), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
NAND3xp33_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1272), .C(n_1274), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1257), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1254), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_1252), .A2(n_1256), .B1(n_1277), .B2(n_1278), .C(n_1280), .Y(n_1276) );
OAI31xp33_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1285), .A3(n_1293), .B(n_1294), .Y(n_1274) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1454 ( .A(n_1283), .Y(n_1454) );
OAI31xp33_ASAP7_75t_L g1671 ( .A1(n_1294), .A2(n_1672), .A3(n_1673), .B(n_1682), .Y(n_1671) );
XNOR2xp5_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1347), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AOI211x1_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1313), .B(n_1314), .C(n_1329), .Y(n_1298) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
AOI221x1_ASAP7_75t_L g1596 ( .A1(n_1313), .A2(n_1550), .B1(n_1597), .B2(n_1608), .C(n_1621), .Y(n_1596) );
AOI31xp33_ASAP7_75t_L g1314 ( .A1(n_1315), .A2(n_1322), .A3(n_1325), .B(n_1328), .Y(n_1314) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
AOI31xp33_ASAP7_75t_L g1387 ( .A1(n_1328), .A2(n_1388), .A3(n_1391), .B(n_1395), .Y(n_1387) );
AO21x1_ASAP7_75t_SL g1415 ( .A1(n_1328), .A2(n_1416), .B(n_1421), .Y(n_1415) );
CKINVDCx16_ASAP7_75t_R g1550 ( .A(n_1328), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1342), .Y(n_1329) );
BUFx3_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx3_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
XNOR2x1_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1397), .Y(n_1347) );
NAND3xp33_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1356), .C(n_1359), .Y(n_1350) );
NAND4xp25_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1371), .C(n_1378), .D(n_1382), .Y(n_1362) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1367), .C(n_1368), .Y(n_1363) );
INVx3_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1630 ( .A(n_1368), .B(n_1631), .C(n_1632), .Y(n_1630) );
INVx3_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1376), .Y(n_1567) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1376), .Y(n_1677) );
INVx5_ASAP7_75t_SL g1450 ( .A(n_1393), .Y(n_1450) );
AND4x1_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1415), .C(n_1424), .D(n_1430), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g1438 ( .A(n_1399), .B(n_1415), .C(n_1424), .D(n_1430), .Y(n_1438) );
OAI31xp33_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1407), .A3(n_1410), .B(n_1414), .Y(n_1399) );
NAND3xp33_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1403), .C(n_1406), .Y(n_1400) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1412), .Y(n_1468) );
OAI31xp33_ASAP7_75t_SL g1461 ( .A1(n_1414), .A2(n_1462), .A3(n_1463), .B(n_1464), .Y(n_1461) );
INVx1_ASAP7_75t_SL g1593 ( .A(n_1414), .Y(n_1593) );
OAI21xp33_ASAP7_75t_L g1519 ( .A1(n_1419), .A2(n_1520), .B(n_1521), .Y(n_1519) );
NAND3xp33_ASAP7_75t_L g1622 ( .A(n_1425), .B(n_1623), .C(n_1625), .Y(n_1622) );
HB1xp67_ASAP7_75t_L g1958 ( .A(n_1435), .Y(n_1958) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
XNOR2x1_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1546), .Y(n_1441) );
XNOR2x1_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1505), .Y(n_1442) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1444), .Y(n_1503) );
OAI22xp33_ASAP7_75t_L g1485 ( .A1(n_1446), .A2(n_1481), .B1(n_1486), .B2(n_1487), .Y(n_1485) );
NAND4xp25_ASAP7_75t_SL g1551 ( .A(n_1452), .B(n_1552), .C(n_1555), .D(n_1558), .Y(n_1551) );
NAND4xp25_ASAP7_75t_SL g1608 ( .A(n_1452), .B(n_1609), .C(n_1612), .D(n_1619), .Y(n_1608) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1459), .Y(n_1457) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1492), .Y(n_1471) );
OAI22xp5_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1475), .B1(n_1476), .B2(n_1477), .Y(n_1473) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
OAI22xp33_ASAP7_75t_SL g1479 ( .A1(n_1480), .A2(n_1481), .B1(n_1482), .B2(n_1483), .Y(n_1479) );
OAI22xp33_ASAP7_75t_L g1652 ( .A1(n_1481), .A2(n_1653), .B1(n_1654), .B2(n_1656), .Y(n_1652) );
INVx1_ASAP7_75t_L g1952 ( .A(n_1483), .Y(n_1952) );
BUFx2_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1484), .Y(n_1655) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
NAND4xp25_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1532), .C(n_1543), .D(n_1545), .Y(n_1506) );
OAI221xp5_ASAP7_75t_L g1508 ( .A1(n_1509), .A2(n_1513), .B1(n_1516), .B2(n_1519), .C(n_1523), .Y(n_1508) );
INVx2_ASAP7_75t_L g1569 ( .A(n_1511), .Y(n_1569) );
INVx2_ASAP7_75t_SL g1624 ( .A(n_1511), .Y(n_1624) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
OA22x2_ASAP7_75t_L g1546 ( .A1(n_1547), .A2(n_1594), .B1(n_1595), .B2(n_1639), .Y(n_1546) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1547), .Y(n_1639) );
XNOR2xp5_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
AOI211xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1551), .B(n_1563), .C(n_1581), .Y(n_1549) );
NAND2xp5_ASAP7_75t_SL g1563 ( .A(n_1564), .B(n_1571), .Y(n_1563) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
AOI31xp33_ASAP7_75t_SL g1581 ( .A1(n_1582), .A2(n_1588), .A3(n_1590), .B(n_1593), .Y(n_1581) );
INVx2_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1586), .Y(n_1605) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1596), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1601), .Y(n_1597) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
HB1xp67_ASAP7_75t_L g1986 ( .A(n_1618), .Y(n_1986) );
NAND4xp25_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1626), .C(n_1630), .D(n_1633), .Y(n_1621) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1641), .Y(n_1690) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
AND4x1_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1666), .C(n_1669), .D(n_1671), .Y(n_1645) );
INVx1_ASAP7_75t_L g2020 ( .A(n_1649), .Y(n_2020) );
OAI22xp5_ASAP7_75t_L g1674 ( .A1(n_1650), .A2(n_1651), .B1(n_1675), .B2(n_1676), .Y(n_1674) );
INVx2_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVx2_ASAP7_75t_SL g1662 ( .A(n_1663), .Y(n_1662) );
NOR2xp33_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1668), .Y(n_1666) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
INVx2_ASAP7_75t_SL g1679 ( .A(n_1680), .Y(n_1679) );
INVx2_ASAP7_75t_SL g1680 ( .A(n_1681), .Y(n_1680) );
OAI221xp5_ASAP7_75t_L g1691 ( .A1(n_1692), .A2(n_1929), .B1(n_1931), .B2(n_1996), .C(n_2000), .Y(n_1691) );
AOI311xp33_ASAP7_75t_L g1692 ( .A1(n_1693), .A2(n_1788), .A3(n_1816), .B(n_1823), .C(n_1895), .Y(n_1692) );
OAI211xp5_ASAP7_75t_L g1693 ( .A1(n_1694), .A2(n_1722), .B(n_1748), .C(n_1774), .Y(n_1693) );
A2O1A1Ixp33_ASAP7_75t_L g1748 ( .A1(n_1694), .A2(n_1749), .B(n_1753), .C(n_1759), .Y(n_1748) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1840 ( .A(n_1695), .B(n_1841), .Y(n_1840) );
AND2x2_ASAP7_75t_L g1922 ( .A(n_1695), .B(n_1817), .Y(n_1922) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx2_ASAP7_75t_SL g1764 ( .A(n_1696), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_1696), .B(n_1756), .Y(n_1799) );
AND2x4_ASAP7_75t_L g1813 ( .A(n_1696), .B(n_1755), .Y(n_1813) );
NAND2xp5_ASAP7_75t_L g1838 ( .A(n_1696), .B(n_1817), .Y(n_1838) );
AND2x2_ASAP7_75t_L g1844 ( .A(n_1696), .B(n_1845), .Y(n_1844) );
NOR2xp33_ASAP7_75t_L g1886 ( .A(n_1696), .B(n_1845), .Y(n_1886) );
HB1xp67_ASAP7_75t_L g1913 ( .A(n_1696), .Y(n_1913) );
CKINVDCx5p33_ASAP7_75t_R g1696 ( .A(n_1697), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1778 ( .A(n_1697), .B(n_1756), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1851 ( .A(n_1697), .B(n_1755), .Y(n_1851) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1712), .Y(n_1697) );
OAI22xp5_ASAP7_75t_L g1698 ( .A1(n_1699), .A2(n_1706), .B1(n_1707), .B2(n_1711), .Y(n_1698) );
BUFx3_ASAP7_75t_L g1785 ( .A(n_1699), .Y(n_1785) );
BUFx6f_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
OAI22xp5_ASAP7_75t_L g1745 ( .A1(n_1700), .A2(n_1709), .B1(n_1746), .B2(n_1747), .Y(n_1745) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1702), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1701), .B(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1701), .Y(n_1729) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1702), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1705), .Y(n_1702) );
HB1xp67_ASAP7_75t_L g2054 ( .A(n_1703), .Y(n_2054) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1705), .Y(n_1716) );
HB1xp67_ASAP7_75t_L g1787 ( .A(n_1707), .Y(n_1787) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1710), .Y(n_1731) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1713), .A2(n_1718), .B1(n_1719), .B2(n_1721), .Y(n_1712) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
BUFx3_ASAP7_75t_L g1782 ( .A(n_1714), .Y(n_1782) );
AND2x4_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1717), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1715), .B(n_1717), .Y(n_1738) );
HB1xp67_ASAP7_75t_L g2052 ( .A(n_1715), .Y(n_2052) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
AND2x4_ASAP7_75t_L g1720 ( .A(n_1716), .B(n_1717), .Y(n_1720) );
INVx2_ASAP7_75t_L g1781 ( .A(n_1719), .Y(n_1781) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1719), .Y(n_1930) );
INVx2_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
XNOR2x1_ASAP7_75t_L g1932 ( .A(n_1721), .B(n_1933), .Y(n_1932) );
OR2x2_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1733), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1750 ( .A(n_1723), .B(n_1751), .Y(n_1750) );
OAI321xp33_ASAP7_75t_SL g1836 ( .A1(n_1723), .A2(n_1837), .A3(n_1838), .B1(n_1839), .B2(n_1840), .C(n_1842), .Y(n_1836) );
NAND2xp5_ASAP7_75t_L g1848 ( .A(n_1723), .B(n_1766), .Y(n_1848) );
INVx2_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1835 ( .A(n_1724), .B(n_1739), .Y(n_1835) );
NAND2xp5_ASAP7_75t_SL g1870 ( .A(n_1724), .B(n_1871), .Y(n_1870) );
AND2x2_ASAP7_75t_L g1901 ( .A(n_1724), .B(n_1799), .Y(n_1901) );
BUFx2_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1762 ( .A(n_1725), .B(n_1763), .Y(n_1762) );
INVx2_ASAP7_75t_L g1770 ( .A(n_1725), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1725), .B(n_1792), .Y(n_1791) );
OR2x2_ASAP7_75t_L g1809 ( .A(n_1725), .B(n_1797), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1725), .B(n_1752), .Y(n_1828) );
INVx2_ASAP7_75t_L g1845 ( .A(n_1725), .Y(n_1845) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1732), .Y(n_1725) );
AND2x4_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1729), .Y(n_1727) );
AND2x4_ASAP7_75t_L g1730 ( .A(n_1729), .B(n_1731), .Y(n_1730) );
BUFx2_ASAP7_75t_L g1821 ( .A(n_1730), .Y(n_1821) );
INVx2_ASAP7_75t_L g1775 ( .A(n_1733), .Y(n_1775) );
NAND2xp5_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1739), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1734), .B(n_1762), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1734), .B(n_1772), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1734), .B(n_1767), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1734), .B(n_1777), .Y(n_1798) );
INVxp67_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
BUFx2_ASAP7_75t_L g1752 ( .A(n_1735), .Y(n_1752) );
BUFx3_ASAP7_75t_L g1797 ( .A(n_1735), .Y(n_1797) );
OR2x2_ASAP7_75t_L g1881 ( .A(n_1735), .B(n_1744), .Y(n_1881) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1736), .B(n_1737), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1739), .B(n_1797), .Y(n_1796) );
NOR2xp33_ASAP7_75t_L g1879 ( .A(n_1739), .B(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1739), .Y(n_1890) );
NAND3xp33_ASAP7_75t_SL g1908 ( .A(n_1739), .B(n_1769), .C(n_1832), .Y(n_1908) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1743), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1740), .B(n_1744), .Y(n_1763) );
INVx2_ASAP7_75t_L g1768 ( .A(n_1740), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1773 ( .A(n_1740), .B(n_1744), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1843 ( .A(n_1740), .B(n_1797), .Y(n_1843) );
NOR2xp33_ASAP7_75t_L g1871 ( .A(n_1740), .B(n_1797), .Y(n_1871) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1742), .Y(n_1740) );
NOR2x1_ASAP7_75t_L g1751 ( .A(n_1743), .B(n_1752), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1894 ( .A(n_1743), .B(n_1797), .Y(n_1894) );
INVx2_ASAP7_75t_SL g1743 ( .A(n_1744), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1744), .B(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
NOR2xp33_ASAP7_75t_L g1906 ( .A(n_1750), .B(n_1853), .Y(n_1906) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1751), .Y(n_1892) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1752), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1752), .B(n_1763), .Y(n_1815) );
A2O1A1Ixp33_ASAP7_75t_L g1759 ( .A1(n_1753), .A2(n_1760), .B(n_1764), .C(n_1765), .Y(n_1759) );
OAI221xp5_ASAP7_75t_L g1800 ( .A1(n_1753), .A2(n_1754), .B1(n_1801), .B2(n_1803), .C(n_1805), .Y(n_1800) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
AOI22xp33_ASAP7_75t_L g1910 ( .A1(n_1754), .A2(n_1789), .B1(n_1851), .B2(n_1911), .Y(n_1910) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1841 ( .A(n_1755), .B(n_1819), .Y(n_1841) );
OR2x2_ASAP7_75t_L g1853 ( .A(n_1755), .B(n_1854), .Y(n_1853) );
INVx3_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
OR2x2_ASAP7_75t_L g1877 ( .A(n_1756), .B(n_1819), .Y(n_1877) );
AND2x2_ASAP7_75t_L g1918 ( .A(n_1756), .B(n_1818), .Y(n_1918) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1757), .B(n_1758), .Y(n_1756) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1762), .Y(n_1839) );
O2A1O1Ixp33_ASAP7_75t_L g1896 ( .A1(n_1762), .A2(n_1897), .B(n_1898), .C(n_1899), .Y(n_1896) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1763), .Y(n_1802) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_1763), .B(n_1770), .Y(n_1804) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1764), .B(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1764), .Y(n_1790) );
NOR2xp33_ASAP7_75t_L g1807 ( .A(n_1764), .B(n_1808), .Y(n_1807) );
NOR2xp33_ASAP7_75t_L g1867 ( .A(n_1764), .B(n_1853), .Y(n_1867) );
INVx2_ASAP7_75t_L g1875 ( .A(n_1764), .Y(n_1875) );
AOI21xp33_ASAP7_75t_SL g1765 ( .A1(n_1766), .A2(n_1769), .B(n_1771), .Y(n_1765) );
OAI211xp5_ASAP7_75t_L g1864 ( .A1(n_1766), .A2(n_1845), .B(n_1851), .C(n_1865), .Y(n_1864) );
A2O1A1Ixp33_ASAP7_75t_SL g1909 ( .A1(n_1766), .A2(n_1883), .B(n_1910), .C(n_1915), .Y(n_1909) );
AND2x2_ASAP7_75t_L g1827 ( .A(n_1767), .B(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1767), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1837 ( .A(n_1768), .B(n_1797), .Y(n_1837) );
OAI321xp33_ASAP7_75t_L g1899 ( .A1(n_1768), .A2(n_1888), .A3(n_1900), .B1(n_1902), .B2(n_1903), .C(n_1905), .Y(n_1899) );
NOR2xp33_ASAP7_75t_L g1772 ( .A(n_1770), .B(n_1773), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1770), .B(n_1777), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1904 ( .A(n_1770), .B(n_1843), .Y(n_1904) );
INVx1_ASAP7_75t_L g1914 ( .A(n_1771), .Y(n_1914) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1773), .Y(n_1777) );
OR2x2_ASAP7_75t_L g1808 ( .A(n_1773), .B(n_1809), .Y(n_1808) );
NOR2xp33_ASAP7_75t_L g1849 ( .A(n_1773), .B(n_1850), .Y(n_1849) );
O2A1O1Ixp33_ASAP7_75t_L g1774 ( .A1(n_1775), .A2(n_1776), .B(n_1778), .C(n_1779), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1897 ( .A(n_1776), .B(n_1797), .Y(n_1897) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1777), .B(n_1828), .Y(n_1876) );
CKINVDCx5p33_ASAP7_75t_R g1833 ( .A(n_1778), .Y(n_1833) );
AOI211xp5_ASAP7_75t_SL g1846 ( .A1(n_1778), .A2(n_1847), .B(n_1849), .C(n_1852), .Y(n_1846) );
NAND4xp25_ASAP7_75t_L g1926 ( .A(n_1778), .B(n_1828), .C(n_1865), .D(n_1927), .Y(n_1926) );
INVx3_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
INVx3_ASAP7_75t_L g1805 ( .A(n_1780), .Y(n_1805) );
A2O1A1Ixp33_ASAP7_75t_SL g1823 ( .A1(n_1780), .A2(n_1824), .B(n_1846), .C(n_1862), .Y(n_1823) );
AND2x2_ASAP7_75t_L g1883 ( .A(n_1780), .B(n_1884), .Y(n_1883) );
OAI22xp33_ASAP7_75t_L g1783 ( .A1(n_1784), .A2(n_1785), .B1(n_1786), .B2(n_1787), .Y(n_1783) );
NAND4xp25_ASAP7_75t_L g1788 ( .A(n_1789), .B(n_1793), .C(n_1806), .D(n_1810), .Y(n_1788) );
OR2x2_ASAP7_75t_L g1789 ( .A(n_1790), .B(n_1791), .Y(n_1789) );
INVx1_ASAP7_75t_L g1917 ( .A(n_1791), .Y(n_1917) );
AOI21xp33_ASAP7_75t_L g1793 ( .A1(n_1794), .A2(n_1799), .B(n_1800), .Y(n_1793) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
NOR2xp33_ASAP7_75t_L g1795 ( .A(n_1796), .B(n_1798), .Y(n_1795) );
OR2x2_ASAP7_75t_L g1801 ( .A(n_1797), .B(n_1802), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1856 ( .A(n_1797), .B(n_1804), .Y(n_1856) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1798), .Y(n_1887) );
AOI221xp5_ASAP7_75t_L g1824 ( .A1(n_1799), .A2(n_1825), .B1(n_1829), .B2(n_1834), .C(n_1836), .Y(n_1824) );
AOI21xp5_ASAP7_75t_L g1915 ( .A1(n_1799), .A2(n_1813), .B(n_1855), .Y(n_1915) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1801), .Y(n_1872) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1816 ( .A(n_1805), .B(n_1817), .Y(n_1816) );
O2A1O1Ixp33_ASAP7_75t_L g1873 ( .A1(n_1805), .A2(n_1835), .B(n_1874), .C(n_1877), .Y(n_1873) );
OAI211xp5_ASAP7_75t_L g1895 ( .A1(n_1805), .A2(n_1896), .B(n_1909), .C(n_1916), .Y(n_1895) );
INVxp67_ASAP7_75t_SL g1806 ( .A(n_1807), .Y(n_1806) );
O2A1O1Ixp33_ASAP7_75t_L g1916 ( .A1(n_1807), .A2(n_1917), .B(n_1918), .C(n_1919), .Y(n_1916) );
NAND2xp5_ASAP7_75t_L g1825 ( .A(n_1808), .B(n_1826), .Y(n_1825) );
NOR2xp33_ASAP7_75t_L g1925 ( .A(n_1808), .B(n_1913), .Y(n_1925) );
OR2x2_ASAP7_75t_L g1889 ( .A(n_1809), .B(n_1890), .Y(n_1889) );
INVxp67_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
NOR2xp33_ASAP7_75t_L g1811 ( .A(n_1812), .B(n_1814), .Y(n_1811) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
AND2x2_ASAP7_75t_L g1861 ( .A(n_1813), .B(n_1817), .Y(n_1861) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
OAI332xp33_ASAP7_75t_L g1878 ( .A1(n_1816), .A2(n_1875), .A3(n_1879), .B1(n_1882), .B2(n_1885), .B3(n_1887), .C1(n_1888), .C2(n_1889), .Y(n_1878) );
INVx2_ASAP7_75t_L g1865 ( .A(n_1817), .Y(n_1865) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1818), .Y(n_1832) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1819), .Y(n_1854) );
INVx1_ASAP7_75t_L g1902 ( .A(n_1819), .Y(n_1902) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1820), .B(n_1822), .Y(n_1819) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1866 ( .A(n_1827), .B(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
OR2x2_ASAP7_75t_L g1830 ( .A(n_1831), .B(n_1833), .Y(n_1830) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1832), .Y(n_1884) );
AOI211xp5_ASAP7_75t_L g1891 ( .A1(n_1832), .A2(n_1850), .B(n_1892), .C(n_1893), .Y(n_1891) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1898 ( .A(n_1838), .Y(n_1898) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1841), .Y(n_1888) );
NAND2xp5_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1844), .Y(n_1842) );
NAND2xp5_ASAP7_75t_L g1850 ( .A(n_1845), .B(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
OAI21xp33_ASAP7_75t_L g1852 ( .A1(n_1853), .A2(n_1855), .B(n_1857), .Y(n_1852) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
INVxp33_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
NOR2xp33_ASAP7_75t_L g1858 ( .A(n_1859), .B(n_1860), .Y(n_1858) );
NAND2xp5_ASAP7_75t_L g1928 ( .A(n_1859), .B(n_1890), .Y(n_1928) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
OAI21xp5_ASAP7_75t_L g1868 ( .A1(n_1861), .A2(n_1869), .B(n_1872), .Y(n_1868) );
NOR4xp25_ASAP7_75t_L g1862 ( .A(n_1863), .B(n_1873), .C(n_1878), .D(n_1891), .Y(n_1862) );
NAND3xp33_ASAP7_75t_L g1863 ( .A(n_1864), .B(n_1866), .C(n_1868), .Y(n_1863) );
A2O1A1Ixp33_ASAP7_75t_L g1919 ( .A1(n_1865), .A2(n_1920), .B(n_1924), .C(n_1926), .Y(n_1919) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1875), .B(n_1876), .Y(n_1874) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1881), .Y(n_1880) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1883), .Y(n_1882) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVxp67_ASAP7_75t_L g1923 ( .A(n_1889), .Y(n_1923) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1894), .Y(n_1893) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1904), .Y(n_1903) );
NOR2xp33_ASAP7_75t_L g1905 ( .A(n_1906), .B(n_1907), .Y(n_1905) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
INVxp33_ASAP7_75t_L g1911 ( .A(n_1912), .Y(n_1911) );
NOR2xp33_ASAP7_75t_L g1912 ( .A(n_1913), .B(n_1914), .Y(n_1912) );
NAND2xp5_ASAP7_75t_L g1920 ( .A(n_1921), .B(n_1923), .Y(n_1920) );
INVx1_ASAP7_75t_L g1921 ( .A(n_1922), .Y(n_1921) );
INVx1_ASAP7_75t_L g1924 ( .A(n_1925), .Y(n_1924) );
INVx1_ASAP7_75t_L g1927 ( .A(n_1928), .Y(n_1927) );
INVx1_ASAP7_75t_L g1929 ( .A(n_1930), .Y(n_1929) );
INVx2_ASAP7_75t_SL g1931 ( .A(n_1932), .Y(n_1931) );
AND2x2_ASAP7_75t_L g1933 ( .A(n_1934), .B(n_1969), .Y(n_1933) );
AOI21xp5_ASAP7_75t_L g1934 ( .A1(n_1935), .A2(n_1936), .B(n_1937), .Y(n_1934) );
AOI31xp33_ASAP7_75t_L g1937 ( .A1(n_1938), .A2(n_1953), .A3(n_1964), .B(n_1967), .Y(n_1937) );
AOI211xp5_ASAP7_75t_SL g1938 ( .A1(n_1939), .A2(n_1940), .B(n_1942), .C(n_1946), .Y(n_1938) );
INVx1_ASAP7_75t_L g1940 ( .A(n_1941), .Y(n_1940) );
INVx3_ASAP7_75t_L g1944 ( .A(n_1945), .Y(n_1944) );
OAI21xp5_ASAP7_75t_SL g1947 ( .A1(n_1948), .A2(n_1950), .B(n_1951), .Y(n_1947) );
INVx1_ASAP7_75t_L g1948 ( .A(n_1949), .Y(n_1948) );
AOI221xp5_ASAP7_75t_L g1953 ( .A1(n_1954), .A2(n_1956), .B1(n_1957), .B2(n_1961), .C(n_1963), .Y(n_1953) );
CKINVDCx5p33_ASAP7_75t_R g1954 ( .A(n_1955), .Y(n_1954) );
INVx1_ASAP7_75t_L g1959 ( .A(n_1960), .Y(n_1959) );
INVx1_ASAP7_75t_SL g1967 ( .A(n_1968), .Y(n_1967) );
NOR2xp33_ASAP7_75t_L g1969 ( .A(n_1970), .B(n_1980), .Y(n_1969) );
INVx1_ASAP7_75t_L g1971 ( .A(n_1972), .Y(n_1971) );
INVx1_ASAP7_75t_L g1973 ( .A(n_1974), .Y(n_1973) );
AOI22xp33_ASAP7_75t_L g1975 ( .A1(n_1976), .A2(n_1977), .B1(n_1978), .B2(n_1979), .Y(n_1975) );
NAND2xp5_ASAP7_75t_SL g1980 ( .A(n_1981), .B(n_1990), .Y(n_1980) );
AOI221xp5_ASAP7_75t_L g1990 ( .A1(n_1991), .A2(n_1992), .B1(n_1993), .B2(n_1994), .C(n_1995), .Y(n_1990) );
INVx4_ASAP7_75t_SL g1996 ( .A(n_1997), .Y(n_1996) );
BUFx3_ASAP7_75t_L g1997 ( .A(n_1998), .Y(n_1997) );
BUFx2_ASAP7_75t_L g1998 ( .A(n_1999), .Y(n_1998) );
INVx1_ASAP7_75t_L g2001 ( .A(n_2002), .Y(n_2001) );
CKINVDCx5p33_ASAP7_75t_R g2002 ( .A(n_2003), .Y(n_2002) );
A2O1A1Ixp33_ASAP7_75t_L g2050 ( .A1(n_2004), .A2(n_2051), .B(n_2053), .C(n_2055), .Y(n_2050) );
INVxp33_ASAP7_75t_L g2005 ( .A(n_2006), .Y(n_2005) );
INVx1_ASAP7_75t_L g2047 ( .A(n_2008), .Y(n_2047) );
HB1xp67_ASAP7_75t_L g2008 ( .A(n_2009), .Y(n_2008) );
AND4x1_ASAP7_75t_L g2009 ( .A(n_2010), .B(n_2023), .C(n_2025), .D(n_2044), .Y(n_2009) );
OAI22xp5_ASAP7_75t_L g2028 ( .A1(n_2029), .A2(n_2030), .B1(n_2031), .B2(n_2034), .Y(n_2028) );
INVx1_ASAP7_75t_L g2031 ( .A(n_2032), .Y(n_2031) );
INVx1_ASAP7_75t_L g2032 ( .A(n_2033), .Y(n_2032) );
NOR2xp33_ASAP7_75t_L g2044 ( .A(n_2045), .B(n_2046), .Y(n_2044) );
BUFx2_ASAP7_75t_L g2048 ( .A(n_2049), .Y(n_2048) );
HB1xp67_ASAP7_75t_L g2049 ( .A(n_2050), .Y(n_2049) );
INVx1_ASAP7_75t_L g2051 ( .A(n_2052), .Y(n_2051) );
INVx1_ASAP7_75t_L g2053 ( .A(n_2054), .Y(n_2053) );
endmodule