module fake_jpeg_2010_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx13_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_82),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_1),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_56),
.B1(n_74),
.B2(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_76),
.B1(n_80),
.B2(n_68),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_83),
.B1(n_78),
.B2(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_108),
.B1(n_61),
.B2(n_73),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_75),
.B(n_51),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_54),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.C(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_63),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_62),
.B1(n_64),
.B2(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_73),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_64),
.B1(n_61),
.B2(n_71),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_70),
.B1(n_69),
.B2(n_67),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_52),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_51),
.B(n_55),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_59),
.B(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_53),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_1),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_117),
.C(n_111),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_158),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_65),
.B(n_59),
.Y(n_152)
);

OAI221xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_160),
.C(n_163),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_65),
.B(n_59),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_125),
.C(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_2),
.Y(n_160)
);

NOR4xp25_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_49),
.C(n_45),
.D(n_43),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_125),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_172),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_40),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_171),
.C(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_37),
.C(n_29),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_170),
.C(n_177),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_174),
.B1(n_176),
.B2(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_27),
.C(n_25),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_24),
.B(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_21),
.B(n_20),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_7),
.C(n_8),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_154),
.C(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_179),
.C(n_173),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_142),
.A3(n_157),
.B1(n_143),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_176),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_192),
.B1(n_197),
.B2(n_190),
.Y(n_198)
);

FAx1_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_181),
.CI(n_175),
.CON(n_192),
.SN(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.C(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_186),
.B1(n_183),
.B2(n_17),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_15),
.Y(n_197)
);

OAI211xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_199),
.B(n_200),
.C(n_192),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_192),
.A3(n_195),
.B(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_15),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_19),
.B(n_16),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_16),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_18),
.Y(n_208)
);


endmodule