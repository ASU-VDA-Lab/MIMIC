module real_aes_133_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_841, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_841;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g221 ( .A(n_0), .B(n_158), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_1), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_2), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g130 ( .A(n_3), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_4), .B(n_134), .Y(n_179) );
NAND2xp33_ASAP7_75t_SL g241 ( .A(n_5), .B(n_140), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_6), .A2(n_103), .B1(n_829), .B2(n_838), .Y(n_102) );
INVx1_ASAP7_75t_L g233 ( .A(n_7), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_8), .B(n_184), .Y(n_457) );
INVx1_ASAP7_75t_L g501 ( .A(n_9), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g836 ( .A(n_10), .Y(n_836) );
AND2x2_ASAP7_75t_L g177 ( .A(n_11), .B(n_163), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_12), .Y(n_493) );
INVx2_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_14), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g834 ( .A(n_14), .B(n_835), .C(n_837), .Y(n_834) );
INVx1_ASAP7_75t_L g466 ( .A(n_15), .Y(n_466) );
AOI221x1_ASAP7_75t_L g236 ( .A1(n_16), .A2(n_142), .B1(n_237), .B2(n_239), .C(n_240), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_17), .B(n_134), .Y(n_201) );
INVx1_ASAP7_75t_L g446 ( .A(n_18), .Y(n_446) );
INVx1_ASAP7_75t_L g464 ( .A(n_19), .Y(n_464) );
INVx1_ASAP7_75t_SL g560 ( .A(n_20), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_21), .B(n_135), .Y(n_534) );
AOI33xp33_ASAP7_75t_L g510 ( .A1(n_22), .A2(n_54), .A3(n_127), .B1(n_147), .B2(n_511), .B3(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_23), .A2(n_142), .B(n_181), .Y(n_180) );
AOI221xp5_ASAP7_75t_SL g210 ( .A1(n_24), .A2(n_41), .B1(n_134), .B2(n_142), .C(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_25), .B(n_158), .Y(n_182) );
INVx1_ASAP7_75t_L g487 ( .A(n_26), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_27), .Y(n_813) );
OAI22x1_ASAP7_75t_R g107 ( .A1(n_28), .A2(n_52), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_28), .Y(n_109) );
OA21x2_ASAP7_75t_L g121 ( .A1(n_29), .A2(n_91), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g164 ( .A(n_29), .B(n_91), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_156), .Y(n_205) );
INVxp67_ASAP7_75t_L g235 ( .A(n_31), .Y(n_235) );
AND2x2_ASAP7_75t_L g174 ( .A(n_32), .B(n_162), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_33), .B(n_125), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_34), .A2(n_142), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_35), .B(n_156), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_36), .A2(n_53), .B1(n_646), .B2(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_36), .Y(n_826) );
AND2x2_ASAP7_75t_L g132 ( .A(n_37), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g140 ( .A(n_37), .B(n_130), .Y(n_140) );
INVx1_ASAP7_75t_L g146 ( .A(n_37), .Y(n_146) );
OR2x6_ASAP7_75t_L g444 ( .A(n_38), .B(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g837 ( .A(n_38), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_39), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_40), .B(n_125), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_42), .A2(n_184), .B1(n_217), .B2(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_43), .B(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_44), .A2(n_83), .B1(n_142), .B2(n_144), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_45), .B(n_135), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_46), .B(n_158), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_47), .B(n_120), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_48), .B(n_135), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_49), .Y(n_531) );
AND2x2_ASAP7_75t_L g224 ( .A(n_50), .B(n_162), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_51), .B(n_162), .Y(n_214) );
INVx1_ASAP7_75t_L g108 ( .A(n_52), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_53), .Y(n_646) );
HB1xp67_ASAP7_75t_SL g717 ( .A(n_53), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_55), .B(n_135), .Y(n_479) );
OAI22x1_ASAP7_75t_R g824 ( .A1(n_56), .A2(n_825), .B1(n_827), .B2(n_828), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_56), .Y(n_828) );
INVx1_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
INVx1_ASAP7_75t_L g137 ( .A(n_57), .Y(n_137) );
AND2x2_ASAP7_75t_L g480 ( .A(n_58), .B(n_162), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_59), .A2(n_76), .B1(n_125), .B2(n_144), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_60), .B(n_125), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_61), .B(n_134), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_62), .B(n_217), .Y(n_495) );
AOI21xp5_ASAP7_75t_SL g520 ( .A1(n_63), .A2(n_144), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g165 ( .A(n_64), .B(n_162), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_65), .B(n_156), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_66), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_67), .B(n_163), .Y(n_206) );
INVx1_ASAP7_75t_L g460 ( .A(n_68), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_69), .A2(n_142), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g478 ( .A(n_70), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_71), .B(n_156), .Y(n_183) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_72), .B(n_120), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_73), .A2(n_144), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g133 ( .A(n_74), .Y(n_133) );
INVx1_ASAP7_75t_L g139 ( .A(n_74), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_75), .B(n_125), .Y(n_513) );
AND2x2_ASAP7_75t_L g562 ( .A(n_77), .B(n_239), .Y(n_562) );
INVx1_ASAP7_75t_L g462 ( .A(n_78), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_79), .A2(n_144), .B(n_559), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_80), .A2(n_119), .B(n_144), .C(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_81), .A2(n_86), .B1(n_125), .B2(n_134), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_82), .B(n_134), .Y(n_160) );
INVx1_ASAP7_75t_L g447 ( .A(n_84), .Y(n_447) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_85), .B(n_239), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_87), .A2(n_144), .B1(n_508), .B2(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_88), .B(n_158), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_89), .B(n_158), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_90), .A2(n_142), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g522 ( .A(n_92), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_93), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g514 ( .A(n_94), .B(n_239), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_95), .A2(n_485), .B(n_486), .C(n_488), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_96), .B(n_134), .Y(n_223) );
INVxp67_ASAP7_75t_L g238 ( .A(n_97), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_98), .B(n_156), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_99), .A2(n_142), .B(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g808 ( .A(n_100), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_101), .B(n_135), .Y(n_523) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_804), .B(n_814), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_799), .Y(n_104) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_110), .B(n_794), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp33_ASAP7_75t_L g799 ( .A(n_107), .B(n_800), .Y(n_799) );
OAI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_441), .B1(n_448), .B2(n_790), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g800 ( .A1(n_112), .A2(n_449), .B1(n_801), .B2(n_802), .Y(n_800) );
AND3x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_312), .C(n_386), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_254), .C(n_285), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_187), .B(n_196), .C(n_225), .Y(n_114) );
AOI21x1_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_166), .B(n_185), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_116), .A2(n_288), .B1(n_294), .B2(n_297), .Y(n_287) );
AND2x2_ASAP7_75t_L g421 ( .A(n_116), .B(n_189), .Y(n_421) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_150), .Y(n_116) );
BUFx2_ASAP7_75t_L g192 ( .A(n_117), .Y(n_192) );
AND2x2_ASAP7_75t_L g280 ( .A(n_117), .B(n_151), .Y(n_280) );
AND2x2_ASAP7_75t_L g351 ( .A(n_117), .B(n_195), .Y(n_351) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_118), .Y(n_245) );
AOI21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_149), .Y(n_118) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_119), .A2(n_506), .B(n_514), .Y(n_505) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_119), .A2(n_506), .B(n_514), .Y(n_577) );
INVx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_120), .A2(n_201), .B(n_202), .Y(n_200) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_120), .A2(n_499), .B(n_503), .Y(n_498) );
BUFx4f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g217 ( .A(n_121), .Y(n_217) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_122), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g184 ( .A(n_122), .B(n_164), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_141), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_125), .A2(n_144), .B1(n_232), .B2(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g496 ( .A(n_125), .Y(n_496) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
INVx1_ASAP7_75t_L g529 ( .A(n_126), .Y(n_529) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
OR2x6_ASAP7_75t_L g461 ( .A(n_127), .B(n_148), .Y(n_461) );
INVxp33_ASAP7_75t_L g511 ( .A(n_127), .Y(n_511) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g143 ( .A(n_128), .B(n_130), .Y(n_143) );
AND2x4_ASAP7_75t_L g156 ( .A(n_128), .B(n_138), .Y(n_156) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g530 ( .A(n_131), .Y(n_530) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x6_ASAP7_75t_L g142 ( .A(n_132), .B(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
AND2x6_ASAP7_75t_L g158 ( .A(n_133), .B(n_136), .Y(n_158) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
INVx1_ASAP7_75t_L g242 ( .A(n_135), .Y(n_242) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_140), .Y(n_488) );
AND2x4_ASAP7_75t_L g144 ( .A(n_143), .B(n_145), .Y(n_144) );
INVxp67_ASAP7_75t_L g494 ( .A(n_144), .Y(n_494) );
NOR2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g512 ( .A(n_147), .Y(n_512) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g244 ( .A(n_150), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g186 ( .A(n_151), .B(n_176), .Y(n_186) );
OR2x2_ASAP7_75t_L g194 ( .A(n_151), .B(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g249 ( .A(n_151), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g296 ( .A(n_151), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_151), .B(n_195), .Y(n_304) );
AND2x2_ASAP7_75t_L g341 ( .A(n_151), .B(n_245), .Y(n_341) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_151), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_151), .B(n_175), .Y(n_382) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_161), .B(n_165), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_160), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
INVxp67_ASAP7_75t_L g467 ( .A(n_156), .Y(n_467) );
INVxp67_ASAP7_75t_L g465 ( .A(n_158), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_159), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_159), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_159), .A2(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_159), .B(n_184), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_159), .A2(n_461), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_159), .A2(n_461), .B(n_501), .C(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g508 ( .A(n_159), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_159), .A2(n_461), .B(n_522), .C(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_159), .A2(n_534), .B(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_159), .A2(n_461), .B(n_560), .C(n_561), .Y(n_559) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_161), .A2(n_168), .B(n_174), .Y(n_167) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_168), .B(n_174), .Y(n_195) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_161), .A2(n_556), .B(n_562), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_162), .Y(n_161) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_162), .A2(n_210), .B(n_214), .Y(n_209) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g283 ( .A(n_166), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_166), .B(n_244), .Y(n_339) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_166), .Y(n_440) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_175), .Y(n_166) );
AND2x2_ASAP7_75t_L g185 ( .A(n_167), .B(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g265 ( .A(n_167), .B(n_176), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_167), .B(n_296), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_173), .Y(n_168) );
AND2x2_ASAP7_75t_L g332 ( .A(n_175), .B(n_249), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_175), .B(n_244), .Y(n_388) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g190 ( .A(n_176), .Y(n_190) );
AND2x2_ASAP7_75t_L g259 ( .A(n_176), .B(n_250), .Y(n_259) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
AND2x4_ASAP7_75t_L g286 ( .A(n_176), .B(n_195), .Y(n_286) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_176), .B(n_245), .Y(n_433) );
OR2x6_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_184), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_184), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_184), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_184), .B(n_238), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g240 ( .A(n_184), .B(n_241), .C(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_184), .A2(n_520), .B(n_524), .Y(n_519) );
INVx1_ASAP7_75t_L g412 ( .A(n_185), .Y(n_412) );
INVx1_ASAP7_75t_L g354 ( .A(n_186), .Y(n_354) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_191), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g276 ( .A(n_190), .B(n_194), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_190), .B(n_245), .Y(n_369) );
AND2x2_ASAP7_75t_L g371 ( .A(n_190), .B(n_193), .Y(n_371) );
AOI32xp33_ASAP7_75t_L g437 ( .A1(n_190), .A2(n_253), .A3(n_408), .B1(n_438), .B2(n_440), .Y(n_437) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
AND2x2_ASAP7_75t_L g263 ( .A(n_192), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g381 ( .A(n_192), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g404 ( .A(n_192), .B(n_265), .Y(n_404) );
AND2x2_ASAP7_75t_L g431 ( .A(n_192), .B(n_332), .Y(n_431) );
AND2x2_ASAP7_75t_L g357 ( .A(n_193), .B(n_245), .Y(n_357) );
AND2x2_ASAP7_75t_L g432 ( .A(n_193), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g290 ( .A(n_198), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g308 ( .A(n_198), .Y(n_308) );
OR2x2_ASAP7_75t_L g336 ( .A(n_198), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x4_ASAP7_75t_SL g253 ( .A(n_199), .B(n_230), .Y(n_253) );
AND2x4_ASAP7_75t_L g269 ( .A(n_199), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g272 ( .A(n_199), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g300 ( .A(n_199), .B(n_209), .Y(n_300) );
OR2x2_ASAP7_75t_L g325 ( .A(n_199), .B(n_274), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_199), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_199), .B(n_209), .Y(n_360) );
INVx2_ASAP7_75t_L g376 ( .A(n_199), .Y(n_376) );
AND2x2_ASAP7_75t_L g391 ( .A(n_199), .B(n_229), .Y(n_391) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_199), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_199), .Y(n_420) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_206), .Y(n_199) );
AND2x2_ASAP7_75t_L g284 ( .A(n_207), .B(n_269), .Y(n_284) );
AND2x2_ASAP7_75t_L g305 ( .A(n_207), .B(n_253), .Y(n_305) );
INVx1_ASAP7_75t_L g337 ( .A(n_207), .Y(n_337) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_215), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g228 ( .A(n_209), .Y(n_228) );
INVx2_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
BUFx3_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
AND2x2_ASAP7_75t_L g330 ( .A(n_209), .B(n_215), .Y(n_330) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_209), .Y(n_428) );
INVx2_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
INVx1_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
OR2x2_ASAP7_75t_L g273 ( .A(n_215), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g293 ( .A(n_215), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_215), .B(n_270), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_215), .B(n_376), .Y(n_375) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_224), .Y(n_216) );
INVx4_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_217), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_244), .B(n_246), .Y(n_225) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_227), .Y(n_436) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_228), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_228), .B(n_268), .Y(n_310) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_228), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_229), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g315 ( .A(n_229), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g366 ( .A(n_229), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_229), .A2(n_371), .B1(n_372), .B2(n_377), .C(n_380), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_229), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_243), .Y(n_229) );
INVx3_ASAP7_75t_L g270 ( .A(n_230), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_230), .B(n_274), .Y(n_374) );
AND2x2_ASAP7_75t_L g403 ( .A(n_230), .B(n_376), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_230), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_236), .Y(n_230) );
INVx3_ASAP7_75t_L g473 ( .A(n_239), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_239), .A2(n_473), .B1(n_484), .B2(n_489), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_242), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_242), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g311 ( .A(n_244), .B(n_286), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_244), .A2(n_264), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g248 ( .A(n_245), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g257 ( .A(n_245), .Y(n_257) );
OR2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_245), .B(n_286), .Y(n_395) );
OR2x2_ASAP7_75t_L g427 ( .A(n_245), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g439 ( .A(n_245), .B(n_345), .Y(n_439) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx2_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
INVx3_ASAP7_75t_SL g383 ( .A(n_249), .Y(n_383) );
INVxp67_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AOI322xp5_ASAP7_75t_L g255 ( .A1(n_253), .A2(n_256), .A3(n_260), .B1(n_263), .B2(n_266), .C1(n_271), .C2(n_275), .Y(n_255) );
INVx1_ASAP7_75t_SL g344 ( .A(n_253), .Y(n_344) );
AND2x4_ASAP7_75t_L g429 ( .A(n_253), .B(n_316), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_277), .Y(n_254) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OR2x2_ASAP7_75t_L g282 ( .A(n_257), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g378 ( .A(n_257), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g406 ( .A(n_257), .B(n_259), .Y(n_406) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_257), .A2(n_258), .A3(n_408), .B1(n_410), .B2(n_413), .Y(n_407) );
OR2x2_ASAP7_75t_L g411 ( .A(n_257), .B(n_304), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g367 ( .A(n_258), .B(n_283), .C(n_368), .Y(n_367) );
OAI22xp33_ASAP7_75t_SL g387 ( .A1(n_258), .A2(n_324), .B1(n_388), .B2(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g390 ( .A(n_261), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_265), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI322xp33_ASAP7_75t_L g313 ( .A1(n_269), .A2(n_273), .A3(n_282), .B1(n_314), .B2(n_317), .C1(n_318), .C2(n_319), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_269), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_269), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g324 ( .A(n_270), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_270), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g385 ( .A(n_273), .Y(n_385) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_284), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_280), .B(n_328), .Y(n_327) );
AOI322xp5_ASAP7_75t_SL g422 ( .A1(n_280), .A2(n_286), .A3(n_403), .B1(n_421), .B2(n_423), .C1(n_426), .C2(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_301), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_286), .B(n_296), .Y(n_318) );
INVx2_ASAP7_75t_SL g328 ( .A(n_286), .Y(n_328) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_SL g353 ( .A(n_292), .Y(n_353) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g398 ( .A(n_299), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_353), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_306), .B2(n_311), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR4xp75_ASAP7_75t_L g312 ( .A(n_313), .B(n_326), .C(n_346), .D(n_362), .Y(n_312) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_324), .A2(n_401), .B1(n_404), .B2(n_405), .Y(n_400) );
OR2x2_ASAP7_75t_L g365 ( .A(n_325), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g409 ( .A(n_325), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_334), .Y(n_326) );
INVx2_ASAP7_75t_L g345 ( .A(n_330), .Y(n_345) );
AND2x2_ASAP7_75t_L g402 ( .A(n_330), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .B1(n_340), .B2(n_342), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g397 ( .A(n_341), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_342), .A2(n_348), .B1(n_364), .B2(n_367), .Y(n_363) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_352), .B1(n_354), .B2(n_355), .C(n_841), .Y(n_346) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g414 ( .A(n_353), .B(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_370), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_384), .Y(n_380) );
NOR3xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_392), .C(n_416), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_407), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_398), .C(n_400), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g408 ( .A(n_399), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
NAND4xp25_ASAP7_75t_SL g416 ( .A(n_417), .B(n_422), .C(n_430), .D(n_437), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_432), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx11_ASAP7_75t_R g803 ( .A(n_441), .Y(n_803) );
OR2x6_ASAP7_75t_SL g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AND2x6_ASAP7_75t_SL g793 ( .A(n_442), .B(n_444), .Y(n_793) );
OR2x2_ASAP7_75t_L g798 ( .A(n_442), .B(n_444), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_442), .B(n_443), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g833 ( .A(n_445), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI211x1_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_646), .B(n_647), .C(n_787), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND4x1_ASAP7_75t_L g787 ( .A(n_451), .B(n_648), .C(n_788), .D(n_789), .Y(n_787) );
NAND3x1_ASAP7_75t_L g822 ( .A(n_451), .B(n_648), .C(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_614), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_537), .B(n_549), .C(n_590), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_469), .B(n_515), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_SL g537 ( .A1(n_455), .A2(n_538), .B(n_543), .C(n_548), .Y(n_537) );
NAND2x1_ASAP7_75t_L g667 ( .A(n_455), .B(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_455), .B(n_687), .Y(n_758) );
AND2x2_ASAP7_75t_L g777 ( .A(n_455), .B(n_517), .Y(n_777) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g554 ( .A(n_456), .Y(n_554) );
AND2x2_ASAP7_75t_L g625 ( .A(n_456), .B(n_555), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_456), .B(n_526), .Y(n_630) );
NOR2x1_ASAP7_75t_SL g746 ( .A(n_456), .B(n_517), .Y(n_746) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_463), .B(n_468), .Y(n_458) );
INVxp67_ASAP7_75t_L g485 ( .A(n_461), .Y(n_485) );
INVx2_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_463) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_497), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_471), .B(n_595), .Y(n_661) );
AND2x2_ASAP7_75t_L g778 ( .A(n_471), .B(n_619), .Y(n_778) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_472), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g567 ( .A(n_472), .Y(n_567) );
AND2x2_ASAP7_75t_L g575 ( .A(n_472), .B(n_576), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g713 ( .A(n_472), .B(n_481), .Y(n_713) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_480), .Y(n_472) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_473), .A2(n_474), .B(n_480), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x2_ASAP7_75t_L g665 ( .A(n_481), .B(n_505), .Y(n_665) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g541 ( .A(n_482), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g545 ( .A(n_482), .Y(n_545) );
INVx1_ASAP7_75t_L g565 ( .A(n_482), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_482), .B(n_598), .Y(n_622) );
AND2x2_ASAP7_75t_L g671 ( .A(n_482), .B(n_498), .Y(n_671) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_490), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g626 ( .A(n_497), .B(n_621), .Y(n_626) );
AND2x2_ASAP7_75t_L g682 ( .A(n_497), .B(n_565), .Y(n_682) );
AND2x2_ASAP7_75t_L g697 ( .A(n_497), .B(n_611), .Y(n_697) );
AND2x2_ASAP7_75t_L g734 ( .A(n_497), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g750 ( .A(n_497), .Y(n_750) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
INVx2_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
INVx1_ASAP7_75t_L g547 ( .A(n_498), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_498), .B(n_577), .Y(n_580) );
INVx1_ASAP7_75t_L g594 ( .A(n_498), .Y(n_594) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_498), .Y(n_604) );
INVxp67_ASAP7_75t_L g620 ( .A(n_498), .Y(n_620) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
AND2x4_ASAP7_75t_L g566 ( .A(n_505), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g548 ( .A(n_515), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_515), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_SL g569 ( .A(n_516), .B(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_516), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_516), .B(n_583), .Y(n_726) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_516), .Y(n_764) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
INVx2_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
AND2x2_ASAP7_75t_L g600 ( .A(n_517), .B(n_526), .Y(n_600) );
INVx4_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_517), .B(n_584), .Y(n_644) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_517), .Y(n_657) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x4_ASAP7_75t_L g635 ( .A(n_525), .B(n_608), .Y(n_635) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g586 ( .A(n_526), .B(n_554), .Y(n_586) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_526), .Y(n_607) );
INVx2_ASAP7_75t_L g656 ( .A(n_526), .Y(n_656) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .C(n_531), .Y(n_528) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_539), .B(n_544), .Y(n_645) );
NAND2x1_ASAP7_75t_SL g759 ( .A(n_539), .B(n_541), .Y(n_759) );
OR2x2_ASAP7_75t_L g638 ( .A(n_540), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g741 ( .A(n_540), .Y(n_741) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g631 ( .A(n_541), .B(n_566), .Y(n_631) );
AND2x2_ASAP7_75t_L g747 ( .A(n_541), .B(n_740), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_543), .A2(n_756), .B1(n_759), .B2(n_760), .C(n_762), .Y(n_755) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_544), .A2(n_700), .B1(n_702), .B2(n_704), .Y(n_699) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_545), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g613 ( .A(n_545), .Y(n_613) );
BUFx2_ASAP7_75t_L g694 ( .A(n_545), .Y(n_694) );
AND2x2_ASAP7_75t_L g664 ( .A(n_546), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_568), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_563), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g637 ( .A(n_553), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g762 ( .A(n_553), .B(n_763), .C(n_764), .D(n_765), .Y(n_762) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
AND2x2_ASAP7_75t_L g655 ( .A(n_554), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx2_ASAP7_75t_L g585 ( .A(n_555), .Y(n_585) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_555), .Y(n_612) );
INVx1_ASAP7_75t_L g629 ( .A(n_555), .Y(n_629) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_555), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g776 ( .A(n_564), .Y(n_776) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g574 ( .A(n_565), .Y(n_574) );
AND2x2_ASAP7_75t_L g670 ( .A(n_566), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g770 ( .A(n_566), .B(n_771), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_573), .B1(n_578), .B2(n_581), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_570), .B(n_635), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_570), .B(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g751 ( .A(n_570), .B(n_729), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_570), .A2(n_606), .B(n_728), .Y(n_781) );
AND2x4_ASAP7_75t_SL g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_571), .B(n_655), .Y(n_692) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_571), .Y(n_708) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_574), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g595 ( .A(n_576), .Y(n_595) );
AND2x2_ASAP7_75t_L g619 ( .A(n_576), .B(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g740 ( .A(n_576), .B(n_597), .Y(n_740) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_577), .B(n_598), .Y(n_639) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g715 ( .A(n_580), .B(n_622), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .Y(n_581) );
INVx1_ASAP7_75t_L g696 ( .A(n_582), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_583), .B(n_592), .C(n_596), .Y(n_591) );
AND2x2_ASAP7_75t_L g634 ( .A(n_583), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g663 ( .A(n_583), .B(n_606), .Y(n_663) );
AND2x2_ASAP7_75t_L g745 ( .A(n_583), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g771 ( .A(n_583), .Y(n_771) );
INVx1_ASAP7_75t_L g785 ( .A(n_583), .Y(n_785) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g588 ( .A(n_586), .B(n_589), .Y(n_588) );
INVx4_ASAP7_75t_L g744 ( .A(n_586), .Y(n_744) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g784 ( .A(n_588), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
AO22x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_599), .B1(n_601), .B2(n_609), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_593), .B(n_597), .Y(n_677) );
INVx3_ASAP7_75t_L g711 ( .A(n_593), .Y(n_711) );
BUFx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g611 ( .A(n_597), .Y(n_611) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g689 ( .A(n_598), .B(n_604), .Y(n_689) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_598), .Y(n_736) );
AOI31xp33_ASAP7_75t_L g640 ( .A1(n_599), .A2(n_641), .A3(n_643), .B(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_600), .A2(n_617), .B1(n_623), .B2(n_626), .Y(n_616) );
AND2x2_ASAP7_75t_L g700 ( .A(n_600), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_600), .B(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_606), .B(n_761), .Y(n_760) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g636 ( .A(n_608), .B(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_608), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g731 ( .A(n_611), .B(n_671), .Y(n_731) );
INVx1_ASAP7_75t_L g766 ( .A(n_611), .Y(n_766) );
AND2x2_ASAP7_75t_L g716 ( .A(n_612), .B(n_655), .Y(n_716) );
BUFx2_ASAP7_75t_L g761 ( .A(n_612), .Y(n_761) );
AND2x2_ASAP7_75t_L g704 ( .A(n_613), .B(n_705), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_632), .C(n_640), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_627), .Y(n_615) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g693 ( .A(n_619), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_625), .B(n_635), .Y(n_658) );
AND2x2_ASAP7_75t_L g680 ( .A(n_625), .B(n_657), .Y(n_680) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_625), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
AND2x2_ASAP7_75t_L g783 ( .A(n_628), .B(n_657), .Y(n_783) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x2_ASAP7_75t_L g757 ( .A(n_629), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g674 ( .A(n_630), .Y(n_674) );
AND2x2_ASAP7_75t_L g774 ( .A(n_630), .B(n_657), .Y(n_774) );
AOI21xp33_ASAP7_75t_R g632 ( .A1(n_633), .A2(n_636), .B(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_634), .B(n_738), .Y(n_737) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_635), .Y(n_642) );
INVx1_ASAP7_75t_L g705 ( .A(n_639), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_641), .A2(n_659), .B1(n_673), .B2(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g673 ( .A(n_644), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_646), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_646), .B(n_753), .Y(n_752) );
NOR2xp67_ASAP7_75t_SL g788 ( .A(n_646), .B(n_719), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_717), .B(n_718), .C(n_752), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_683), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .C(n_678), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_659), .B(n_662), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_658), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_654), .A2(n_693), .B1(n_696), .B2(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g730 ( .A(n_656), .Y(n_730) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g722 ( .A(n_661), .B(n_711), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_670), .Y(n_662) );
INVx1_ASAP7_75t_L g676 ( .A(n_665), .Y(n_676) );
AND2x4_ASAP7_75t_L g688 ( .A(n_665), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g724 ( .A(n_667), .Y(n_724) );
INVx1_ASAP7_75t_L g701 ( .A(n_668), .Y(n_701) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_670), .A2(n_680), .B1(n_728), .B2(n_731), .Y(n_727) );
INVxp67_ASAP7_75t_L g772 ( .A(n_671), .Y(n_772) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_674), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVxp33_ASAP7_75t_L g786 ( .A(n_677), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_698), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_695), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_690), .B2(n_693), .Y(n_685) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_699), .B(n_706), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_714), .B2(n_716), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g763 ( .A(n_711), .Y(n_763) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g823 ( .A(n_720), .B(n_754), .Y(n_823) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_732), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_727), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND4xp25_ASAP7_75t_SL g732 ( .A(n_733), .B(n_737), .C(n_742), .D(n_748), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g775 ( .A(n_740), .B(n_776), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .B(n_747), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g789 ( .A(n_753), .Y(n_789) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR3x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_767), .C(n_779), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_772), .B(n_773), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_773) );
INVx1_ASAP7_75t_L g780 ( .A(n_778), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B(n_782), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B(n_786), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
CKINVDCx6p67_ASAP7_75t_R g801 ( .A(n_791), .Y(n_801) );
INVx3_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_808), .Y(n_815) );
INVxp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_810), .A2(n_817), .B(n_820), .Y(n_816) );
NOR2xp33_ASAP7_75t_SL g810 ( .A(n_811), .B(n_813), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g819 ( .A(n_812), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_825), .Y(n_827) );
BUFx3_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g839 ( .A(n_831), .Y(n_839) );
INVx2_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_SL g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
endmodule