module fake_jpeg_11207_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_54),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_16),
.C(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_42),
.C(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_64),
.B1(n_50),
.B2(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_46),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_51),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_69),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_35),
.B(n_39),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_60),
.B1(n_64),
.B2(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_0),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_1),
.B(n_3),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_79),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_20),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_88),
.B1(n_10),
.B2(n_13),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_22),
.C(n_32),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_15),
.C(n_21),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_4),
.C(n_5),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_96)
);

AOI21x1_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_102),
.B(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.C(n_104),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_23),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_90),
.C(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.C(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_89),
.B1(n_101),
.B2(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

AOI211xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_111),
.B(n_110),
.C(n_109),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_106),
.CON(n_118),
.SN(n_118)
);


endmodule