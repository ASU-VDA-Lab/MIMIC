module real_jpeg_14028_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_255)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_57),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_6),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_6),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_7),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_122),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_122),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_122),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_69),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_30),
.C(n_45),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_78),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_113),
.B(n_166),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_59),
.B(n_77),
.C(n_193),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_11),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_11),
.B(n_54),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_162),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_162),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_40),
.B1(n_42),
.B2(n_80),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_80),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_15),
.B(n_60),
.Y(n_251)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_323),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_310),
.B(n_322),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_138),
.B(n_307),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_125),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_100),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_22),
.B(n_100),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_70),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_23),
.B(n_71),
.C(n_86),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_52),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_24),
.A2(n_25),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_26),
.A2(n_27),
.B1(n_52),
.B2(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_28),
.A2(n_32),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_167),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_28),
.A2(n_32),
.B1(n_112),
.B2(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_29),
.B(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_32),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_34),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_51),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_38),
.A2(n_43),
.B1(n_51),
.B2(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_42),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_40),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_42),
.A2(n_76),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_43),
.A2(n_51),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_43),
.B(n_152),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_43),
.A2(n_51),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_43),
.A2(n_51),
.B1(n_117),
.B2(n_244),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_49),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_47),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_47),
.B(n_150),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_47),
.A2(n_163),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_51),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_58),
.B1(n_65),
.B2(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_55),
.A2(n_65),
.B(n_150),
.C(n_237),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_55),
.A2(n_59),
.A3(n_62),
.B1(n_238),
.B2(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_68),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_65),
.B1(n_89),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_58),
.A2(n_63),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_58),
.A2(n_65),
.B1(n_121),
.B2(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_64),
.A2(n_218),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_64),
.A2(n_218),
.B1(n_317),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_86),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_72),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_79),
.B1(n_81),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_73),
.A2(n_81),
.B1(n_94),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_73),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_73),
.A2(n_81),
.B1(n_213),
.B2(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_73),
.A2(n_199),
.B(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_78),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_74),
.B(n_200),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_74),
.A2(n_78),
.B(n_314),
.Y(n_313)
);

NOR2x1_ASAP7_75t_R g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_78),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_81),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_81),
.A2(n_119),
.B(n_214),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_84),
.A2(n_151),
.B(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g136 ( 
.A(n_88),
.B(n_91),
.C(n_96),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_88),
.B(n_129),
.C(n_136),
.Y(n_321)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_96),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_96),
.B(n_130),
.C(n_134),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_107),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_106),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_107),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.C(n_120),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_108),
.A2(n_109),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_110),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_113),
.A2(n_114),
.B1(n_195),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_113),
.A2(n_114),
.B1(n_221),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_114),
.A2(n_172),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_150),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_180),
.B(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_118),
.B(n_120),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_124),
.B(n_236),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_125),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_126),
.B(n_137),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_131),
.Y(n_316)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_135),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_301),
.B(n_306),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_289),
.B(n_300),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_257),
.A3(n_282),
.B1(n_287),
.B2(n_288),
.C(n_332),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_230),
.B(n_256),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_207),
.B(n_229),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_188),
.B(n_206),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_168),
.B(n_187),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_176),
.B(n_186),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_174),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_185),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_201),
.C(n_205),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_222),
.B2(n_223),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_225),
.C(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_216),
.C(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_247),
.C(n_248),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_245),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_240),
.C(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_272),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.C(n_271),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_260),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_266),
.C(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_271),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_281),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_276),
.C(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_299),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.C(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_321),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_325),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);


endmodule