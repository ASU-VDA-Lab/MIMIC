module fake_jpeg_11549_n_505 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_505);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_505;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_3),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_49),
.B(n_61),
.Y(n_115)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_52),
.B(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_8),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_14),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_7),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_0),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_89),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_15),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_105),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_25),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_59),
.B(n_21),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_114),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_129),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_63),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_48),
.Y(n_135)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_69),
.B(n_25),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_46),
.B(n_18),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_81),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_64),
.B(n_21),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_173),
.Y(n_219)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_65),
.B1(n_91),
.B2(n_90),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_162),
.B1(n_167),
.B2(n_171),
.Y(n_220)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_161),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_115),
.B1(n_104),
.B2(n_152),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_98),
.A2(n_94),
.B1(n_85),
.B2(n_83),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_163),
.A2(n_187),
.B1(n_123),
.B2(n_86),
.Y(n_208)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_74),
.B1(n_82),
.B2(n_53),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_73),
.B1(n_68),
.B2(n_57),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_42),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_182),
.Y(n_214)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_88),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_42),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_127),
.A2(n_21),
.B(n_27),
.C(n_20),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_58),
.B1(n_66),
.B2(n_28),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_198),
.B1(n_27),
.B2(n_43),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_111),
.A2(n_54),
.B1(n_43),
.B2(n_93),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_16),
.B(n_18),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_110),
.B(n_123),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_196),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_119),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_24),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_228),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_208),
.B1(n_153),
.B2(n_175),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_232),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_227),
.B(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_160),
.A2(n_142),
.B1(n_149),
.B2(n_99),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_163),
.B1(n_187),
.B2(n_192),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_158),
.A2(n_103),
.B(n_101),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_185),
.B(n_150),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_119),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_150),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_183),
.B1(n_155),
.B2(n_191),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_261),
.Y(n_285)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_221),
.B(n_228),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_248),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_218),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_254),
.B1(n_260),
.B2(n_266),
.Y(n_283)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_170),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_256),
.B(n_222),
.Y(n_295)
);

BUFx12_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_253),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_206),
.B1(n_226),
.B2(n_232),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_178),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_219),
.Y(n_276)
);

NAND2x1p5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_178),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_259),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_165),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_220),
.A2(n_193),
.B1(n_133),
.B2(n_164),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_172),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

OR2x2_ASAP7_75t_SL g263 ( 
.A(n_235),
.B(n_156),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_210),
.C(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_265),
.A2(n_267),
.B1(n_166),
.B2(n_211),
.Y(n_289)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_269),
.A2(n_273),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_214),
.C(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_270),
.B(n_272),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_223),
.C(n_219),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_240),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_255),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_210),
.C(n_229),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_260),
.B(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_225),
.B1(n_217),
.B2(n_207),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_222),
.B1(n_233),
.B2(n_112),
.Y(n_330)
);

CKINVDCx10_ASAP7_75t_R g317 ( 
.A(n_289),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_256),
.C(n_259),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_290),
.A2(n_292),
.B(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_210),
.B1(n_202),
.B2(n_224),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_249),
.B1(n_263),
.B2(n_240),
.Y(n_300)
);

AOI32xp33_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_216),
.A3(n_233),
.B1(n_229),
.B2(n_204),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_209),
.C(n_213),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_209),
.C(n_213),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_306),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_302),
.B1(n_308),
.B2(n_315),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_251),
.B1(n_240),
.B2(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_305),
.B(n_270),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_251),
.B1(n_243),
.B2(n_239),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_244),
.B(n_242),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_313),
.A2(n_325),
.B(n_137),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_280),
.A2(n_261),
.B1(n_237),
.B2(n_202),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

CKINVDCx12_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_319),
.Y(n_337)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_286),
.Y(n_320)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_257),
.B1(n_241),
.B2(n_179),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_327),
.B1(n_274),
.B2(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_323),
.Y(n_353)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_288),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_234),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_283),
.A2(n_264),
.B1(n_168),
.B2(n_159),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_277),
.B(n_216),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_329),
.B(n_272),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_192),
.B1(n_130),
.B2(n_113),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_307),
.A2(n_278),
.B(n_276),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_331),
.A2(n_358),
.B(n_330),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_273),
.B(n_271),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

NAND2x1_ASAP7_75t_SL g373 ( 
.A(n_336),
.B(n_329),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_312),
.B1(n_316),
.B2(n_322),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_293),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_313),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_288),
.C(n_282),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_352),
.C(n_362),
.Y(n_371)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_211),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_346),
.B(n_347),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_211),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_350),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_309),
.B(n_275),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_357),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_321),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_275),
.Y(n_351)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_282),
.C(n_189),
.Y(n_352)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_328),
.B(n_231),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_300),
.A2(n_113),
.B1(n_133),
.B2(n_130),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_359),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_360),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_231),
.C(n_197),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_302),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_364),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_349),
.B(n_359),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_315),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_373),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_367),
.A2(n_370),
.B1(n_380),
.B2(n_360),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_325),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_381),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_374),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_324),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_326),
.C(n_323),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_385),
.C(n_390),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_334),
.A2(n_317),
.B1(n_327),
.B2(n_320),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_317),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_265),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_387),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_332),
.C(n_337),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_334),
.B(n_161),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_169),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_389),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_353),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_199),
.C(n_253),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_365),
.A2(n_348),
.B(n_338),
.C(n_358),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_379),
.Y(n_396)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_401),
.Y(n_420)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_391),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_404),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_369),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_361),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_406),
.Y(n_430)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_362),
.C(n_353),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_408),
.B(n_415),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_212),
.B(n_107),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_373),
.B(n_363),
.CI(n_376),
.CON(n_410),
.SN(n_410)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_356),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_350),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_411),
.A2(n_416),
.B(n_177),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_339),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_188),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_383),
.A2(n_376),
.B1(n_377),
.B2(n_375),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_413),
.A2(n_381),
.B1(n_380),
.B2(n_366),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_414),
.A2(n_387),
.B1(n_345),
.B2(n_340),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_377),
.A2(n_361),
.B1(n_340),
.B2(n_355),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_368),
.A2(n_355),
.B(n_345),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_395),
.B(n_364),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_431),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_423),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_421),
.A2(n_393),
.B1(n_410),
.B2(n_149),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_408),
.C(n_412),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g425 ( 
.A(n_399),
.Y(n_425)
);

BUFx24_ASAP7_75t_SL g453 ( 
.A(n_425),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_390),
.C(n_367),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_429),
.Y(n_454)
);

AOI21x1_ASAP7_75t_SL g444 ( 
.A1(n_427),
.A2(n_433),
.B(n_434),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_413),
.A2(n_354),
.B1(n_356),
.B2(n_250),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_428),
.A2(n_414),
.B1(n_393),
.B2(n_398),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_354),
.C(n_253),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_253),
.C(n_250),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_190),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_436),
.B(n_398),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_196),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_392),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_447),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_440),
.A2(n_432),
.B1(n_429),
.B2(n_431),
.Y(n_460)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_402),
.C(n_395),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_448),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_452),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_410),
.B(n_393),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_435),
.B(n_434),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_450),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_99),
.B1(n_131),
.B2(n_120),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_131),
.C(n_114),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_SL g462 ( 
.A(n_451),
.B(n_455),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_196),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_435),
.B(n_428),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_457),
.B(n_468),
.Y(n_478)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_454),
.A2(n_424),
.B1(n_35),
.B2(n_32),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_23),
.B1(n_69),
.B2(n_20),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_442),
.B(n_194),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_466),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_100),
.C(n_194),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_444),
.A2(n_451),
.B(n_446),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_455),
.C(n_452),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_470),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_22),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_461),
.C(n_468),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_19),
.C(n_4),
.Y(n_488)
);

AOI31xp67_ASAP7_75t_L g472 ( 
.A1(n_458),
.A2(n_444),
.A3(n_100),
.B(n_12),
.Y(n_472)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_464),
.B(n_15),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_479),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_SL g475 ( 
.A1(n_456),
.A2(n_14),
.B(n_10),
.C(n_9),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_480),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_467),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_482),
.B(n_466),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_469),
.A2(n_23),
.B1(n_19),
.B2(n_93),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_10),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_485),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_461),
.C(n_462),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_45),
.A3(n_20),
.B1(n_10),
.B2(n_13),
.C1(n_4),
.C2(n_7),
.Y(n_486)
);

OAI321xp33_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_474),
.A3(n_475),
.B1(n_10),
.B2(n_4),
.C(n_13),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_19),
.C(n_7),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_487),
.A2(n_491),
.B(n_483),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_4),
.B(n_14),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_495),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_489),
.A2(n_475),
.B(n_1),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_0),
.C(n_2),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_493),
.A2(n_490),
.B1(n_483),
.B2(n_19),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_498),
.A2(n_494),
.B(n_2),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_499),
.A2(n_2),
.B1(n_3),
.B2(n_497),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_500),
.B(n_501),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_502),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_3),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_3),
.Y(n_505)
);


endmodule