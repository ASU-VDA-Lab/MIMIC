module fake_ariane_779_n_1868 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1868);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1868;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_206;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1759;
wire n_1557;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_66),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_17),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_2),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_116),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_98),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_62),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_28),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_20),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_18),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_69),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_77),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_56),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_12),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_38),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_57),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_38),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_72),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_68),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_85),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_32),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_62),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_80),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_59),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_50),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_155),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_60),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_130),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_31),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_109),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_44),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_153),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_149),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_159),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_122),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_131),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_163),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_49),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_20),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_64),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_55),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_147),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_117),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_54),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_120),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_146),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_71),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_138),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_34),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_156),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_65),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_167),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_86),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_128),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_21),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_100),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_124),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_42),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_91),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_70),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_56),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_59),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_57),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_67),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_46),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_10),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_1),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_55),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_76),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_111),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_162),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_23),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_63),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_89),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_93),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_15),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_107),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_29),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_152),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_151),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_36),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_54),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_63),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_64),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_27),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_43),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_1),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_7),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_7),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_36),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_25),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_110),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_129),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_78),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_19),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_140),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_104),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_43),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_96),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_127),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_37),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_65),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_286),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_198),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_198),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_255),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_181),
.B(n_0),
.Y(n_345)
);

BUFx2_ASAP7_75t_SL g346 ( 
.A(n_170),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_242),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_0),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_172),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_181),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_182),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_218),
.Y(n_359)
);

BUFx2_ASAP7_75t_SL g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_221),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_174),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_3),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_182),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_184),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_265),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_184),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_213),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_191),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_191),
.B(n_3),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_255),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_180),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_194),
.B(n_5),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_311),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_336),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_188),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_213),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_232),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_193),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_197),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_212),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_219),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_219),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_195),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_224),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_224),
.Y(n_391)
);

BUFx2_ASAP7_75t_SL g392 ( 
.A(n_250),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_232),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_230),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_196),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_230),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_200),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_237),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_329),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_243),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_207),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_243),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_215),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_256),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_256),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_227),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_232),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_229),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_234),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_244),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_247),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_259),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_248),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_273),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_273),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_255),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_259),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_343),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_369),
.B(n_177),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_343),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_357),
.B(n_292),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_353),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_358),
.B(n_292),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_261),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_364),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_261),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_368),
.B(n_292),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_337),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_363),
.A2(n_210),
.B1(n_217),
.B2(n_183),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_370),
.B(n_262),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_377),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_377),
.A2(n_267),
.B(n_262),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_267),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_385),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_386),
.B(n_274),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_387),
.B(n_274),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_345),
.B(n_177),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_391),
.B(n_313),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_391),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_347),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_394),
.B(n_313),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_394),
.A2(n_291),
.B(n_250),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_396),
.B(n_313),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_323),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_323),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_473),
.A2(n_379),
.B1(n_346),
.B2(n_360),
.Y(n_493)
);

OA22x2_ASAP7_75t_L g494 ( 
.A1(n_456),
.A2(n_342),
.B1(n_404),
.B2(n_402),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_452),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_404),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_452),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_452),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_434),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_434),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_474),
.B(n_352),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_438),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_455),
.B(n_381),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_434),
.A2(n_393),
.B1(n_409),
.B2(n_382),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

BUFx8_ASAP7_75t_SL g515 ( 
.A(n_455),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_449),
.B(n_360),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_177),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_440),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_474),
.B(n_362),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_250),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_474),
.B(n_373),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_406),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_434),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_449),
.B(n_348),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_463),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_434),
.A2(n_340),
.B1(n_399),
.B2(n_365),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_463),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_474),
.B(n_378),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_440),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_463),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_434),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_474),
.B(n_383),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_434),
.A2(n_371),
.B1(n_374),
.B2(n_201),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_463),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_474),
.B(n_389),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_430),
.B(n_395),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_463),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_482),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_456),
.A2(n_415),
.B1(n_407),
.B2(n_406),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_456),
.A2(n_415),
.B1(n_407),
.B2(n_321),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_463),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_425),
.B(n_321),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_425),
.Y(n_553)
);

NOR2x1p5_ASAP7_75t_L g554 ( 
.A(n_453),
.B(n_339),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_446),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_474),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_487),
.B(n_397),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_446),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_419),
.B(n_437),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_403),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_442),
.Y(n_564)
);

INVx6_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_447),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_419),
.B(n_411),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_474),
.B(n_408),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_474),
.B(n_410),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_482),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_450),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_439),
.B(n_412),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_447),
.A2(n_249),
.B1(n_254),
.B2(n_253),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_468),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_468),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_421),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_468),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_439),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_414),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_443),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_473),
.A2(n_302),
.B(n_278),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_419),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_443),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_468),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_448),
.B(n_416),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_446),
.B(n_323),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_448),
.B(n_273),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_448),
.B(n_273),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_481),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_446),
.B(n_185),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_426),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_448),
.B(n_413),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_462),
.B(n_291),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_476),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_476),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_476),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_437),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_450),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_451),
.B(n_291),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_426),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_450),
.B(n_458),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_417),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g619 ( 
.A(n_451),
.B(n_418),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_426),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_426),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_476),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_421),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_426),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_421),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_462),
.A2(n_454),
.B1(n_479),
.B2(n_446),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_450),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_429),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_451),
.B(n_278),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_428),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_450),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_450),
.Y(n_634)
);

AND3x1_ASAP7_75t_L g635 ( 
.A(n_437),
.B(n_187),
.C(n_185),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_437),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_429),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_458),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_457),
.A2(n_258),
.B1(n_268),
.B2(n_260),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_458),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_429),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_428),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_575),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_599),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_553),
.B(n_458),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_629),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_629),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_553),
.B(n_567),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_583),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_567),
.A2(n_459),
.B1(n_479),
.B2(n_454),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_496),
.B(n_458),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_597),
.B(n_422),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_542),
.A2(n_459),
.B1(n_479),
.B2(n_454),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_496),
.B(n_475),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_575),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_634),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_597),
.B(n_422),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_641),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_641),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_496),
.B(n_517),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_496),
.B(n_475),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_528),
.B(n_584),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_494),
.A2(n_321),
.B1(n_187),
.B2(n_203),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_498),
.Y(n_668)
);

OR2x2_ASAP7_75t_SL g669 ( 
.A(n_515),
.B(n_359),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_597),
.B(n_574),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_526),
.B(n_475),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_565),
.Y(n_673)
);

NOR2x1p5_ASAP7_75t_L g674 ( 
.A(n_568),
.B(n_453),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_498),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_556),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_520),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_526),
.B(n_475),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_529),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_601),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_534),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_558),
.A2(n_459),
.B1(n_479),
.B2(n_454),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_574),
.B(n_422),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_539),
.A2(n_475),
.B1(n_461),
.B2(n_464),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_587),
.B(n_475),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_587),
.B(n_457),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_494),
.A2(n_462),
.B1(n_479),
.B2(n_454),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_574),
.B(n_423),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_611),
.B(n_457),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_594),
.B(n_461),
.Y(n_692)
);

AO221x1_ASAP7_75t_L g693 ( 
.A1(n_493),
.A2(n_177),
.B1(n_241),
.B2(n_223),
.C(n_314),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_561),
.B(n_485),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_574),
.B(n_423),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_561),
.B(n_485),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_556),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_529),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_613),
.B(n_423),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_606),
.B(n_485),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_611),
.B(n_636),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_534),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_534),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_461),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_613),
.B(n_464),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_613),
.B(n_424),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_633),
.B(n_464),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_613),
.B(n_424),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_604),
.B(n_465),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_562),
.B(n_465),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_601),
.B(n_504),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_504),
.B(n_465),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_508),
.B(n_361),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_536),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_505),
.B(n_466),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_505),
.B(n_466),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_527),
.B(n_466),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_527),
.B(n_537),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_552),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_537),
.B(n_470),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_638),
.B(n_470),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_576),
.B(n_460),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_605),
.B(n_424),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_494),
.A2(n_462),
.B1(n_483),
.B2(n_454),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_638),
.B(n_470),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_638),
.B(n_639),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_605),
.B(n_436),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_638),
.B(n_639),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_639),
.B(n_471),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_573),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_536),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_536),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_639),
.B(n_471),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_551),
.B(n_471),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_565),
.B(n_477),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_551),
.B(n_477),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_556),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_551),
.A2(n_539),
.B1(n_493),
.B2(n_523),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_551),
.B(n_477),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_565),
.B(n_478),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_551),
.B(n_478),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_605),
.B(n_436),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_579),
.B(n_478),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_523),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_555),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_620),
.B(n_436),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_510),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_579),
.B(n_480),
.Y(n_755)
);

AND2x6_ASAP7_75t_SL g756 ( 
.A(n_601),
.B(n_199),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_601),
.B(n_485),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_624),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_556),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_554),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_624),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_624),
.B(n_480),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_531),
.B(n_486),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_493),
.A2(n_479),
.B1(n_483),
.B2(n_490),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_627),
.B(n_480),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_620),
.B(n_441),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_576),
.A2(n_467),
.B1(n_469),
.B2(n_472),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_627),
.B(n_490),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_617),
.A2(n_444),
.B(n_441),
.C(n_445),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_619),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_569),
.B(n_490),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_523),
.B(n_492),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_565),
.B(n_492),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_523),
.B(n_492),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_603),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_580),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_640),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_580),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_580),
.B(n_441),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_523),
.B(n_547),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_596),
.B(n_444),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_493),
.A2(n_483),
.B1(n_491),
.B2(n_486),
.Y(n_784)
);

NOR2x1p5_ASAP7_75t_L g785 ( 
.A(n_595),
.B(n_460),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_554),
.B(n_486),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_523),
.B(n_483),
.Y(n_787)
);

OAI22x1_ASAP7_75t_SL g788 ( 
.A1(n_635),
.A2(n_367),
.B1(n_375),
.B2(n_376),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_523),
.B(n_483),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_608),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_559),
.B(n_203),
.C(n_199),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_595),
.B(n_483),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_628),
.A2(n_462),
.B1(n_429),
.B2(n_486),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_555),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_595),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_631),
.A2(n_429),
.B1(n_491),
.B2(n_488),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_595),
.B(n_491),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_548),
.B(n_491),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_635),
.B(n_467),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_608),
.B(n_444),
.Y(n_800)
);

OAI221xp5_ASAP7_75t_L g801 ( 
.A1(n_598),
.A2(n_289),
.B1(n_241),
.B2(n_236),
.C(n_276),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_580),
.B(n_469),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_622),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_621),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_622),
.B(n_445),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_637),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_637),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_615),
.B(n_445),
.C(n_472),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_642),
.B(n_488),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_564),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_642),
.B(n_488),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_631),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_564),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_615),
.B(n_488),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_719),
.A2(n_728),
.B1(n_712),
.B2(n_714),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_773),
.A2(n_670),
.B(n_660),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_670),
.A2(n_570),
.B(n_522),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_654),
.A2(n_660),
.B(n_708),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_665),
.B(n_631),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_665),
.B(n_631),
.Y(n_820)
);

OAI321xp33_ASAP7_75t_L g821 ( 
.A1(n_745),
.A2(n_289),
.A3(n_228),
.B1(n_314),
.B2(n_208),
.C(n_223),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_737),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_712),
.B(n_631),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_713),
.B(n_631),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_631),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_799),
.B(n_768),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_802),
.B(n_564),
.Y(n_827)
);

O2A1O1Ixp5_ASAP7_75t_L g828 ( 
.A1(n_692),
.A2(n_525),
.B(n_533),
.C(n_506),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_695),
.B(n_499),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_723),
.B(n_615),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_692),
.A2(n_541),
.B(n_538),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_669),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_654),
.A2(n_557),
.B(n_518),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_644),
.B(n_489),
.Y(n_834)
);

OAI21xp33_ASAP7_75t_L g835 ( 
.A1(n_646),
.A2(n_277),
.B(n_272),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_795),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_648),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_695),
.B(n_499),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_708),
.A2(n_557),
.B(n_503),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_695),
.B(n_697),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_684),
.A2(n_630),
.B1(n_625),
.B2(n_503),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_697),
.B(n_500),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_730),
.A2(n_501),
.B(n_497),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_730),
.A2(n_749),
.B(n_734),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_734),
.A2(n_557),
.B(n_507),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_742),
.A2(n_630),
.B1(n_625),
.B2(n_507),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_666),
.A2(n_614),
.B1(n_586),
.B2(n_500),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_697),
.B(n_757),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_674),
.B(n_509),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_649),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_742),
.A2(n_630),
.B1(n_625),
.B2(n_511),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_779),
.B(n_509),
.Y(n_853)
);

OAI321xp33_ASAP7_75t_L g854 ( 
.A1(n_801),
.A2(n_276),
.A3(n_236),
.B1(n_228),
.B2(n_208),
.C(n_280),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_749),
.A2(n_557),
.B(n_512),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_655),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_659),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_645),
.B(n_280),
.C(n_190),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_668),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_685),
.A2(n_512),
.B(n_511),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_672),
.A2(n_489),
.B(n_550),
.C(n_519),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_685),
.A2(n_696),
.B(n_690),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_774),
.A2(n_501),
.B(n_497),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_690),
.A2(n_550),
.B(n_519),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_696),
.A2(n_582),
.B(n_572),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_663),
.B(n_572),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_744),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_646),
.A2(n_282),
.B(n_281),
.Y(n_868)
);

AOI33xp33_ASAP7_75t_L g869 ( 
.A1(n_658),
.A2(n_786),
.A3(n_761),
.B1(n_190),
.B2(n_757),
.B3(n_489),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_744),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_757),
.B(n_582),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_733),
.A2(n_589),
.B(n_585),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_798),
.B(n_585),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_704),
.B(n_589),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_797),
.B(n_590),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_714),
.B(n_590),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_736),
.A2(n_484),
.B(n_489),
.C(n_592),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_681),
.B(n_592),
.Y(n_878)
);

AO21x1_ASAP7_75t_L g879 ( 
.A1(n_753),
.A2(n_325),
.B(n_302),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_733),
.A2(n_513),
.B(n_502),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_614),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_679),
.B(n_614),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_698),
.B(n_546),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_744),
.B(n_780),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_702),
.A2(n_513),
.B(n_502),
.Y(n_885)
);

INVxp33_ASAP7_75t_L g886 ( 
.A(n_651),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_702),
.A2(n_516),
.B(n_514),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_666),
.A2(n_614),
.B1(n_586),
.B2(n_429),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_661),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_716),
.B(n_614),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_662),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_709),
.A2(n_516),
.B(n_514),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_795),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_647),
.A2(n_588),
.B(n_609),
.C(n_532),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_682),
.A2(n_614),
.B1(n_626),
.B2(n_623),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_735),
.A2(n_530),
.B(n_521),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_700),
.B(n_284),
.C(n_283),
.Y(n_897)
);

BUFx4f_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_736),
.B(n_747),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_747),
.B(n_614),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_744),
.B(n_524),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_764),
.B(n_495),
.Y(n_902)
);

BUFx8_ASAP7_75t_L g903 ( 
.A(n_682),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_780),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_709),
.A2(n_530),
.B(n_521),
.Y(n_905)
);

AOI21x1_ASAP7_75t_L g906 ( 
.A1(n_776),
.A2(n_535),
.B(n_532),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_754),
.B(n_586),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_775),
.B(n_495),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_780),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_675),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_775),
.B(n_495),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_711),
.A2(n_540),
.B(n_535),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_711),
.A2(n_543),
.B(n_540),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_803),
.A2(n_732),
.B(n_727),
.Y(n_914)
);

CKINVDCx10_ASAP7_75t_R g915 ( 
.A(n_788),
.Y(n_915)
);

CKINVDCx10_ASAP7_75t_R g916 ( 
.A(n_756),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_653),
.B(n_495),
.Y(n_917)
);

BUFx8_ASAP7_75t_L g918 ( 
.A(n_772),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_780),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_687),
.A2(n_577),
.B(n_626),
.C(n_623),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_792),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_688),
.A2(n_577),
.B(n_610),
.C(n_609),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_740),
.A2(n_545),
.B(n_543),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_785),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_657),
.B(n_549),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_664),
.B(n_549),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_741),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_667),
.B(n_549),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_721),
.B(n_549),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_698),
.B(n_571),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_753),
.A2(n_767),
.B(n_808),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_767),
.A2(n_560),
.B(n_545),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_783),
.A2(n_484),
.B(n_325),
.C(n_327),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_673),
.B(n_524),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_790),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_800),
.A2(n_566),
.B(n_560),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_787),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_721),
.B(n_571),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_812),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_691),
.B(n_571),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_789),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_783),
.A2(n_484),
.B(n_327),
.C(n_593),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_707),
.B(n_571),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_804),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_770),
.A2(n_578),
.B(n_566),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_652),
.B(n_612),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_671),
.A2(n_296),
.B(n_285),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_673),
.B(n_524),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_678),
.A2(n_298),
.B(n_297),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_806),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_673),
.A2(n_612),
.B1(n_588),
.B2(n_616),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_591),
.B(n_578),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_677),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_683),
.A2(n_706),
.B(n_705),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_683),
.A2(n_593),
.B(n_591),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_705),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_676),
.B(n_760),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_805),
.A2(n_607),
.B(n_602),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_710),
.B(n_612),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_656),
.A2(n_484),
.B(n_616),
.C(n_610),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_760),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_686),
.A2(n_602),
.B(n_607),
.C(n_612),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_706),
.A2(n_738),
.B(n_717),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_781),
.A2(n_563),
.B(n_524),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_781),
.A2(n_563),
.B(n_524),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_676),
.B(n_524),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_717),
.A2(n_600),
.B(n_546),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_812),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_750),
.A2(n_581),
.B(n_563),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_778),
.B(n_563),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_755),
.A2(n_581),
.B(n_563),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_812),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_738),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_778),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_763),
.A2(n_220),
.B(n_333),
.C(n_264),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_793),
.B(n_766),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_769),
.A2(n_581),
.B(n_563),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_715),
.A2(n_186),
.B(n_231),
.C(n_275),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_751),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_784),
.A2(n_319),
.B(n_299),
.C(n_303),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_782),
.A2(n_433),
.B(n_427),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_680),
.B(n_581),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_743),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_739),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_694),
.B(n_581),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_666),
.Y(n_987)
);

OAI321xp33_ASAP7_75t_L g988 ( 
.A1(n_746),
.A2(n_177),
.A3(n_225),
.B1(n_294),
.B2(n_432),
.C(n_433),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_699),
.B(n_581),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_701),
.B(n_304),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_720),
.B(n_546),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_725),
.B(n_546),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_739),
.Y(n_993)
);

AOI33xp33_ASAP7_75t_L g994 ( 
.A1(n_796),
.A2(n_305),
.A3(n_306),
.B1(n_308),
.B2(n_312),
.B3(n_316),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_729),
.B(n_546),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_759),
.B(n_317),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_751),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_791),
.B(n_318),
.C(n_324),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_748),
.A2(n_320),
.B(n_322),
.C(n_328),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_752),
.A2(n_335),
.B(n_177),
.C(n_334),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_762),
.B(n_546),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_814),
.A2(n_600),
.B(n_643),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_718),
.A2(n_600),
.B(n_643),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_898),
.A2(n_751),
.B1(n_724),
.B2(n_771),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_826),
.A2(n_722),
.B(n_726),
.C(n_807),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_898),
.B(n_689),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_899),
.A2(n_724),
.B(n_811),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_L g1008 ( 
.A1(n_831),
.A2(n_809),
.B(n_810),
.C(n_813),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_836),
.B(n_758),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_822),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_853),
.B(n_902),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_SL g1012 ( 
.A(n_867),
.B(n_600),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_837),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_940),
.B(n_794),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_850),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_853),
.B(n_794),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_886),
.B(n_810),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_902),
.B(n_813),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_867),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_867),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_823),
.A2(n_731),
.B1(n_600),
.B2(n_693),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_927),
.B(n_600),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_903),
.B(n_918),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_848),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_890),
.B(n_836),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_848),
.B(n_295),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_SL g1027 ( 
.A1(n_832),
.A2(n_326),
.B1(n_331),
.B2(n_330),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_998),
.A2(n_924),
.B1(n_942),
.B2(n_938),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_984),
.B(n_643),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_834),
.B(n_878),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_998),
.A2(n_245),
.B1(n_171),
.B2(n_173),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_859),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_910),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_819),
.A2(n_643),
.B(n_632),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_938),
.B(n_942),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_820),
.A2(n_643),
.B1(n_632),
.B2(n_315),
.Y(n_1036)
);

BUFx8_ASAP7_75t_L g1037 ( 
.A(n_940),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_824),
.A2(n_643),
.B1(n_632),
.B2(n_310),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_903),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_921),
.B(n_6),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_940),
.B(n_632),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_851),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_914),
.A2(n_816),
.B(n_929),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_939),
.A2(n_632),
.B(n_433),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_856),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_867),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_840),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_908),
.A2(n_632),
.B(n_433),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_911),
.A2(n_432),
.B(n_427),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_843),
.A2(n_432),
.B(n_427),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_900),
.A2(n_432),
.B(n_427),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_907),
.B(n_9),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_924),
.B(n_169),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_817),
.A2(n_238),
.B(n_176),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_818),
.A2(n_239),
.B(n_178),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_979),
.A2(n_931),
.B(n_976),
.C(n_825),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_918),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_987),
.A2(n_240),
.B1(n_179),
.B2(n_309),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_857),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_893),
.B(n_175),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_960),
.A2(n_246),
.B(n_192),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_940),
.B(n_9),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_969),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_933),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_830),
.A2(n_251),
.B(n_202),
.C(n_307),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_904),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_954),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_873),
.B(n_11),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_916),
.B(n_189),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_977),
.B(n_11),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_968),
.A2(n_252),
.B(n_205),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_830),
.A2(n_257),
.B(n_206),
.C(n_301),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_866),
.B(n_13),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_835),
.B(n_204),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_844),
.B(n_13),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_962),
.B(n_209),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_858),
.A2(n_266),
.B1(n_214),
.B2(n_300),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_999),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_904),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_969),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_858),
.A2(n_263),
.B1(n_216),
.B2(n_222),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_868),
.B(n_211),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_897),
.B(n_226),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_904),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_881),
.A2(n_271),
.B1(n_233),
.B2(n_235),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_849),
.B(n_269),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_880),
.A2(n_287),
.B(n_279),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_962),
.B(n_270),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_999),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_957),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_982),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_969),
.B(n_225),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_974),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_990),
.B(n_83),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_990),
.B(n_24),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_981),
.A2(n_294),
.B(n_225),
.C(n_431),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_969),
.B(n_225),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_889),
.B(n_26),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_975),
.B(n_431),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_891),
.B(n_29),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_970),
.A2(n_428),
.B(n_431),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_827),
.B(n_30),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_973),
.B(n_997),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_973),
.B(n_294),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_981),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_871),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_915),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_904),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_996),
.B(n_869),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_863),
.A2(n_431),
.B(n_428),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_946),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_973),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_975),
.B(n_431),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_919),
.Y(n_1114)
);

CKINVDCx6p67_ASAP7_75t_R g1115 ( 
.A(n_919),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_996),
.A2(n_294),
.B1(n_41),
.B2(n_42),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_948),
.B(n_40),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_829),
.B(n_45),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_919),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_R g1120 ( 
.A(n_973),
.B(n_919),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_985),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_961),
.A2(n_431),
.B(n_428),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_980),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_47),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_972),
.A2(n_428),
.B(n_431),
.Y(n_1125)
);

O2A1O1Ixp5_ASAP7_75t_L g1126 ( 
.A1(n_828),
.A2(n_935),
.B(n_949),
.C(n_901),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_936),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_838),
.B(n_47),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_906),
.A2(n_294),
.B(n_431),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_961),
.A2(n_842),
.B1(n_947),
.B2(n_934),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_978),
.A2(n_431),
.B(n_428),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_950),
.A2(n_48),
.B(n_49),
.C(n_51),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_935),
.A2(n_949),
.B(n_901),
.C(n_884),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_993),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_945),
.B(n_51),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_854),
.A2(n_294),
.B1(n_53),
.B2(n_58),
.C(n_60),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_839),
.A2(n_428),
.B(n_119),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_951),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_876),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_884),
.A2(n_52),
.B(n_53),
.C(n_428),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_874),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_870),
.B(n_73),
.Y(n_1142)
);

CKINVDCx8_ASAP7_75t_R g1143 ( 
.A(n_928),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_928),
.A2(n_79),
.B(n_84),
.C(n_88),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_870),
.B(n_92),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_821),
.B(n_97),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_994),
.B(n_101),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1002),
.A2(n_105),
.B(n_108),
.Y(n_1148)
);

CKINVDCx8_ASAP7_75t_R g1149 ( 
.A(n_1001),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_883),
.B(n_121),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_877),
.A2(n_123),
.B(n_126),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_909),
.B(n_132),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_875),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_934),
.A2(n_141),
.B1(n_154),
.B2(n_158),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_909),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_983),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_958),
.B(n_160),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1025),
.B(n_883),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1011),
.B(n_847),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1116),
.B(n_1000),
.C(n_953),
.Y(n_1160)
);

OA21x2_ASAP7_75t_L g1161 ( 
.A1(n_1122),
.A2(n_877),
.B(n_943),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1011),
.B(n_847),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1043),
.A2(n_896),
.B(n_956),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1122),
.A2(n_1003),
.B(n_943),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1129),
.A2(n_964),
.B(n_955),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1064),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1110),
.A2(n_959),
.B(n_937),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1026),
.A2(n_895),
.B1(n_958),
.B2(n_971),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1095),
.A2(n_1006),
.B1(n_1024),
.B2(n_1028),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1130),
.A2(n_963),
.B(n_882),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1005),
.A2(n_872),
.B(n_922),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1130),
.A2(n_879),
.A3(n_1000),
.B(n_1001),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1153),
.B(n_888),
.Y(n_1173)
);

AND2x6_ASAP7_75t_SL g1174 ( 
.A(n_1023),
.B(n_989),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1050),
.A2(n_923),
.B(n_965),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1150),
.B(n_1009),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1007),
.A2(n_1034),
.B(n_1137),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1016),
.A2(n_941),
.B(n_944),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1024),
.B(n_980),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1114),
.B(n_930),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1016),
.A2(n_966),
.B(n_846),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1101),
.A2(n_865),
.B(n_864),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1009),
.B(n_1030),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1141),
.B(n_888),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1021),
.A2(n_841),
.A3(n_852),
.B(n_952),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1018),
.A2(n_894),
.B(n_920),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1126),
.A2(n_988),
.B(n_932),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1021),
.A2(n_855),
.A3(n_845),
.B(n_995),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1052),
.B(n_917),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1096),
.A2(n_992),
.A3(n_860),
.B(n_833),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1154),
.A2(n_986),
.A3(n_925),
.B(n_926),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1125),
.A2(n_892),
.B(n_913),
.Y(n_1192)
);

NAND3x1_ASAP7_75t_L g1193 ( 
.A(n_1117),
.B(n_1040),
.C(n_1017),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1104),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1094),
.A2(n_861),
.B(n_862),
.C(n_971),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1056),
.A2(n_991),
.B(n_967),
.C(n_885),
.Y(n_1196)
);

AOI31xp67_ASAP7_75t_L g1197 ( 
.A1(n_1075),
.A2(n_967),
.A3(n_991),
.B(n_887),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1035),
.B(n_905),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1131),
.A2(n_912),
.B(n_164),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1154),
.A2(n_165),
.A3(n_1038),
.B(n_1036),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1136),
.A2(n_1105),
.B1(n_1078),
.B2(n_1089),
.C(n_1132),
.Y(n_1201)
);

BUFx12f_ASAP7_75t_L g1202 ( 
.A(n_1057),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1111),
.A2(n_1109),
.B(n_1075),
.C(n_1065),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1018),
.A2(n_1036),
.B(n_1038),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1070),
.A2(n_1008),
.B(n_1133),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_1044),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1032),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1070),
.A2(n_1156),
.A3(n_1146),
.B(n_1048),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1073),
.A2(n_1068),
.B(n_1102),
.Y(n_1209)
);

NAND3x1_ASAP7_75t_L g1210 ( 
.A(n_1031),
.B(n_1074),
.C(n_1082),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1035),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_L g1212 ( 
.A(n_1091),
.B(n_1143),
.C(n_1087),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1124),
.A2(n_1086),
.B1(n_1033),
.B2(n_1090),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1013),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1039),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1077),
.A2(n_1135),
.B1(n_1047),
.B2(n_1025),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1073),
.A2(n_1068),
.B(n_1102),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1012),
.B(n_1084),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1148),
.A2(n_1151),
.B(n_1144),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1107),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1139),
.B(n_1106),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1037),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1151),
.A2(n_1113),
.B(n_1099),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1120),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1138),
.B(n_1042),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1019),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1010),
.B(n_1053),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1072),
.A2(n_1083),
.B(n_1100),
.C(n_1098),
.Y(n_1228)
);

AO32x2_ASAP7_75t_L g1229 ( 
.A1(n_1119),
.A2(n_1027),
.A3(n_1112),
.B1(n_1149),
.B2(n_1140),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1019),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1098),
.A2(n_1100),
.B1(n_1059),
.B2(n_1045),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1092),
.A2(n_1097),
.B(n_1157),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1147),
.A2(n_1128),
.B(n_1118),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1127),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1071),
.A2(n_1029),
.B(n_1152),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1037),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1142),
.A2(n_1041),
.B(n_1123),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1063),
.B(n_1080),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1067),
.B(n_1121),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1093),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1155),
.B(n_1076),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1150),
.A2(n_1054),
.B(n_1055),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1060),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1150),
.A2(n_1088),
.B(n_1061),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1009),
.B(n_1081),
.Y(n_1247)
);

O2A1O1Ixp5_ASAP7_75t_L g1248 ( 
.A1(n_1063),
.A2(n_1080),
.B(n_1022),
.C(n_1112),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1004),
.A2(n_1058),
.B1(n_1085),
.B2(n_1103),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1155),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1022),
.A2(n_1103),
.B(n_1145),
.C(n_1014),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1020),
.A2(n_1046),
.B(n_1066),
.C(n_1079),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1046),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1014),
.A2(n_1104),
.B(n_1066),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1104),
.A2(n_1046),
.B(n_1066),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1079),
.A2(n_1129),
.B(n_1110),
.Y(n_1257)
);

NOR2x1_ASAP7_75t_SL g1258 ( 
.A(n_1079),
.B(n_1108),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1108),
.A2(n_982),
.A3(n_1130),
.B(n_1021),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1006),
.A2(n_754),
.B1(n_510),
.B2(n_381),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1015),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1011),
.A2(n_712),
.B(n_665),
.C(n_719),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1011),
.A2(n_820),
.B(n_819),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1013),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1011),
.A2(n_823),
.B(n_820),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1043),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1122),
.A2(n_1110),
.B(n_982),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1011),
.A2(n_712),
.B(n_665),
.C(n_719),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1043),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1011),
.B(n_826),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1011),
.B(n_826),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1130),
.A2(n_982),
.A3(n_1021),
.B(n_953),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1064),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1011),
.B(n_815),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1057),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1013),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1043),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1011),
.A2(n_823),
.B(n_820),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1283)
);

CKINVDCx12_ASAP7_75t_R g1284 ( 
.A(n_1027),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1015),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1015),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1013),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1122),
.A2(n_1043),
.B(n_1129),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1043),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1011),
.B(n_826),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1043),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1116),
.B(n_712),
.C(n_1117),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1015),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1115),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1064),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1095),
.A2(n_719),
.B(n_562),
.C(n_558),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1011),
.B(n_826),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1011),
.A2(n_823),
.B(n_820),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1130),
.A2(n_982),
.A3(n_1021),
.B(n_953),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1043),
.A2(n_899),
.B(n_823),
.Y(n_1304)
);

O2A1O1Ixp5_ASAP7_75t_SL g1305 ( 
.A1(n_1154),
.A2(n_473),
.B(n_1075),
.C(n_1130),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1011),
.A2(n_823),
.B(n_820),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1011),
.A2(n_826),
.B(n_712),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1011),
.B(n_826),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1208),
.Y(n_1309)
);

CKINVDCx6p67_ASAP7_75t_R g1310 ( 
.A(n_1202),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1292),
.A2(n_1231),
.B1(n_1159),
.B2(n_1162),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1245),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1234),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1214),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1227),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1220),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1239),
.B(n_1189),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1292),
.A2(n_1260),
.B1(n_1307),
.B2(n_1201),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1265),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1211),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1231),
.A2(n_1159),
.B1(n_1162),
.B2(n_1247),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1210),
.A2(n_1284),
.B1(n_1216),
.B2(n_1183),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1280),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1307),
.A2(n_1169),
.B1(n_1278),
.B2(n_1160),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1287),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1213),
.A2(n_1217),
.B1(n_1209),
.B2(n_1275),
.Y(n_1326)
);

INVx6_ASAP7_75t_L g1327 ( 
.A(n_1294),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1212),
.A2(n_1158),
.B1(n_1308),
.B2(n_1273),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1166),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1279),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1212),
.A2(n_1158),
.B1(n_1308),
.B2(n_1275),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1294),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1273),
.A2(n_1290),
.B1(n_1301),
.B2(n_1249),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1209),
.A2(n_1217),
.B1(n_1301),
.B2(n_1290),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1222),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1173),
.A2(n_1184),
.B1(n_1176),
.B2(n_1306),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1193),
.A2(n_1176),
.B1(n_1263),
.B2(n_1269),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1173),
.A2(n_1184),
.B1(n_1176),
.B2(n_1306),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1242),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1266),
.A2(n_1302),
.B1(n_1282),
.B2(n_1221),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1194),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1194),
.A2(n_1232),
.B1(n_1221),
.B2(n_1233),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1266),
.A2(n_1282),
.B1(n_1302),
.B2(n_1233),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1168),
.A2(n_1224),
.B1(n_1296),
.B2(n_1215),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1277),
.Y(n_1345)
);

OAI22x1_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_1236),
.B1(n_1224),
.B2(n_1250),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1207),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1294),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1298),
.A2(n_1228),
.B1(n_1170),
.B2(n_1204),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1170),
.A2(n_1261),
.B1(n_1293),
.B2(n_1286),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1174),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1252),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1241),
.A2(n_1285),
.B1(n_1198),
.B2(n_1161),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1226),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1240),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1161),
.A2(n_1246),
.B1(n_1171),
.B2(n_1186),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1264),
.A2(n_1203),
.B(n_1305),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1226),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1254),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1248),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1226),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1230),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1179),
.A2(n_1244),
.B1(n_1187),
.B2(n_1205),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1230),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1230),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1197),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1196),
.A2(n_1195),
.B1(n_1164),
.B2(n_1205),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1258),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1218),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1163),
.A2(n_1218),
.B1(n_1271),
.B2(n_1274),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1253),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1262),
.A2(n_1304),
.B1(n_1300),
.B2(n_1299),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1180),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1178),
.A2(n_1272),
.B1(n_1297),
.B2(n_1283),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1229),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1256),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1256),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1295),
.A2(n_1200),
.B1(n_1255),
.B2(n_1235),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1238),
.B(n_1172),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1251),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1237),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1276),
.B(n_1303),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1259),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1259),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1223),
.A2(n_1219),
.B1(n_1268),
.B2(n_1181),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1288),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1276),
.B(n_1303),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1172),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1172),
.B(n_1191),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1185),
.B(n_1191),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1288),
.A2(n_1185),
.B1(n_1165),
.B2(n_1177),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1191),
.B(n_1185),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1199),
.A2(n_1167),
.B1(n_1192),
.B2(n_1206),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1188),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1188),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1190),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1190),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1257),
.Y(n_1398)
);

CKINVDCx8_ASAP7_75t_R g1399 ( 
.A(n_1175),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1182),
.A2(n_1267),
.B1(n_1270),
.B2(n_1281),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1289),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1291),
.A2(n_1263),
.B1(n_1269),
.B2(n_815),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1263),
.A2(n_1269),
.B1(n_815),
.B2(n_1292),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1214),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1263),
.A2(n_1269),
.B1(n_815),
.B2(n_1292),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1202),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1214),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1225),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1294),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1245),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1202),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1214),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1292),
.A2(n_508),
.B1(n_815),
.B2(n_716),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1210),
.A2(n_508),
.B1(n_1292),
.B2(n_719),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1166),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1166),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1214),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1292),
.A2(n_716),
.B1(n_754),
.B2(n_359),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1292),
.A2(n_716),
.B1(n_754),
.B2(n_359),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1292),
.A2(n_716),
.B1(n_754),
.B2(n_359),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1292),
.A2(n_1136),
.B1(n_1260),
.B2(n_754),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1225),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1226),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1222),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1292),
.A2(n_716),
.B1(n_754),
.B2(n_359),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1357),
.A2(n_1389),
.B(n_1356),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1313),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1372),
.A2(n_1393),
.B(n_1400),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1398),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1329),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1349),
.A2(n_1405),
.B(n_1403),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1382),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1387),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1314),
.B(n_1319),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1408),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1393),
.A2(n_1400),
.B(n_1374),
.Y(n_1442)
);

AO31x2_ASAP7_75t_L g1443 ( 
.A1(n_1367),
.A2(n_1370),
.A3(n_1392),
.B(n_1309),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1379),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1383),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1383),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1398),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1404),
.B(n_1407),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1427),
.B(n_1320),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1384),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1384),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1380),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1334),
.B(n_1311),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1390),
.B(n_1375),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1413),
.Y(n_1456)
);

CKINVDCx6p67_ASAP7_75t_R g1457 ( 
.A(n_1406),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1388),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1360),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1374),
.A2(n_1385),
.B(n_1391),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1352),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1380),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1388),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1353),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1366),
.A2(n_1333),
.B(n_1337),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1356),
.A2(n_1378),
.B(n_1402),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1359),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1418),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1334),
.B1(n_1324),
.B2(n_1326),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1380),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1414),
.A2(n_1318),
.B(n_1344),
.C(n_1421),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1391),
.A2(n_1396),
.B(n_1378),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1339),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1352),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1396),
.A2(n_1363),
.B(n_1343),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1381),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1401),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1341),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1340),
.B(n_1321),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1343),
.B(n_1340),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1401),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1341),
.A2(n_1415),
.B(n_1346),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1328),
.A2(n_1331),
.B(n_1324),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1381),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1386),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1369),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1363),
.A2(n_1350),
.B(n_1326),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1317),
.B(n_1394),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1350),
.A2(n_1355),
.B(n_1377),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1394),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1395),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1395),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1397),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1347),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1354),
.A2(n_1371),
.B(n_1351),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1397),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1406),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1361),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1376),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1342),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1341),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1322),
.B(n_1358),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1409),
.A2(n_1417),
.B1(n_1416),
.B2(n_1421),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1315),
.B(n_1358),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1361),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1428),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1428),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1409),
.A2(n_1416),
.B(n_1417),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1315),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1498),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1437),
.A2(n_1426),
.B(n_1422),
.C(n_1429),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1467),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1469),
.A2(n_1426),
.B1(n_1422),
.B2(n_1423),
.C(n_1425),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1437),
.A2(n_1430),
.B(n_1424),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1459),
.B(n_1345),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1521)
);

OAI211xp5_ASAP7_75t_L g1522 ( 
.A1(n_1486),
.A2(n_1412),
.B(n_1316),
.C(n_1410),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1469),
.A2(n_1330),
.B1(n_1335),
.B2(n_1348),
.C(n_1373),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1507),
.A2(n_1486),
.B1(n_1513),
.B2(n_1454),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1459),
.B(n_1348),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1433),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1513),
.A2(n_1369),
.B1(n_1412),
.B2(n_1327),
.Y(n_1527)
);

AND2x4_ASAP7_75t_SL g1528 ( 
.A(n_1457),
.B(n_1411),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1435),
.B(n_1312),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1472),
.A2(n_1454),
.B(n_1466),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1513),
.A2(n_1327),
.B1(n_1332),
.B2(n_1310),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1457),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1475),
.B(n_1365),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1503),
.B(n_1365),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1503),
.B(n_1365),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1482),
.A2(n_1327),
.B(n_1332),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_SL g1539 ( 
.A1(n_1482),
.A2(n_1368),
.B(n_1436),
.C(n_1468),
.Y(n_1539)
);

AND2x6_ASAP7_75t_L g1540 ( 
.A(n_1478),
.B(n_1368),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1483),
.A2(n_1368),
.B1(n_1513),
.B2(n_1481),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1435),
.B(n_1448),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1441),
.B(n_1450),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1443),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1485),
.B(n_1494),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_R g1547 ( 
.A(n_1501),
.B(n_1489),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1448),
.B(n_1494),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1440),
.B(n_1447),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_R g1550 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1456),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1447),
.B(n_1449),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1449),
.B(n_1508),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1483),
.A2(n_1481),
.B1(n_1476),
.B2(n_1462),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_SL g1557 ( 
.A(n_1489),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1493),
.B(n_1500),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1502),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1493),
.B(n_1500),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1502),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1497),
.B(n_1478),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1476),
.A2(n_1504),
.B1(n_1464),
.B2(n_1470),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1453),
.A2(n_1462),
.B1(n_1471),
.B2(n_1506),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1431),
.B(n_1487),
.Y(n_1566)
);

OAI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1453),
.A2(n_1471),
.B(n_1460),
.C(n_1504),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1490),
.A2(n_1431),
.B(n_1460),
.C(n_1477),
.Y(n_1568)
);

INVx3_ASAP7_75t_SL g1569 ( 
.A(n_1510),
.Y(n_1569)
);

AOI211xp5_ASAP7_75t_L g1570 ( 
.A1(n_1506),
.A2(n_1490),
.B(n_1434),
.C(n_1442),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1458),
.B(n_1474),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1478),
.B(n_1444),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1442),
.A2(n_1434),
.B(n_1473),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1473),
.A2(n_1477),
.B(n_1499),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1465),
.B(n_1505),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_SL g1576 ( 
.A(n_1465),
.B(n_1480),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1552),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1554),
.B(n_1479),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1515),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1549),
.B(n_1432),
.Y(n_1581)
);

NAND2x1_ASAP7_75t_L g1582 ( 
.A(n_1566),
.B(n_1479),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1554),
.B(n_1479),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1455),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1544),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1526),
.B(n_1465),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1542),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1555),
.B(n_1432),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1518),
.A2(n_1464),
.B1(n_1470),
.B2(n_1465),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1544),
.Y(n_1590)
);

INVxp33_ASAP7_75t_L g1591 ( 
.A(n_1547),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1518),
.A2(n_1446),
.B1(n_1452),
.B2(n_1451),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1529),
.B(n_1509),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1559),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1559),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1577),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1558),
.B(n_1432),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1577),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1528),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1530),
.A2(n_1432),
.B1(n_1492),
.B2(n_1451),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.B(n_1484),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1543),
.B(n_1443),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1517),
.B(n_1443),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1571),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1575),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1538),
.B(n_1443),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1530),
.B(n_1546),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1520),
.B(n_1443),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1556),
.B(n_1488),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1525),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1574),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1524),
.A2(n_1512),
.B1(n_1511),
.B2(n_1509),
.C(n_1463),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1525),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1519),
.A2(n_1452),
.B1(n_1446),
.B2(n_1445),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1521),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1578),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1576),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1589),
.A2(n_1519),
.B1(n_1541),
.B2(n_1564),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1579),
.B(n_1566),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1541),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1579),
.B(n_1583),
.Y(n_1624)
);

AOI33xp33_ASAP7_75t_L g1625 ( 
.A1(n_1592),
.A2(n_1516),
.A3(n_1523),
.B1(n_1514),
.B2(n_1529),
.B3(n_1539),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1581),
.B(n_1568),
.Y(n_1628)
);

OAI211xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1608),
.A2(n_1516),
.B(n_1523),
.C(n_1522),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1613),
.A2(n_1522),
.B1(n_1567),
.B2(n_1527),
.C(n_1531),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1548),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1581),
.B(n_1597),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1567),
.C(n_1512),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1578),
.Y(n_1634)
);

AOI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1607),
.A2(n_1565),
.B(n_1537),
.C(n_1569),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1591),
.B(n_1560),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1585),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1582),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

AOI33xp33_ASAP7_75t_L g1640 ( 
.A1(n_1600),
.A2(n_1542),
.A3(n_1536),
.B1(n_1535),
.B2(n_1572),
.B3(n_1511),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1582),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1609),
.B(n_1488),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1615),
.A2(n_1534),
.B1(n_1566),
.B2(n_1545),
.C(n_1533),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1612),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1551),
.B1(n_1545),
.B2(n_1492),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1580),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1606),
.A2(n_1537),
.B1(n_1540),
.B2(n_1551),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1579),
.B(n_1572),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

AND2x2_ASAP7_75t_SL g1650 ( 
.A(n_1625),
.B(n_1610),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1616),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1644),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1618),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1617),
.B(n_1587),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1638),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.B(n_1587),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1634),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1623),
.B(n_1584),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1627),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1584),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1617),
.B(n_1601),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1646),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1623),
.B(n_1611),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1646),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1614),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1590),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1632),
.B(n_1624),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1627),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1583),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1635),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_R g1676 ( 
.A(n_1628),
.B(n_1545),
.Y(n_1676)
);

NAND2x1_ASAP7_75t_SL g1677 ( 
.A(n_1628),
.B(n_1583),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1632),
.B(n_1601),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1614),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1640),
.B(n_1596),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1635),
.B(n_1640),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1621),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1684),
.B(n_1534),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1653),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1661),
.B(n_1639),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1653),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1651),
.B(n_1625),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1675),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_SL g1695 ( 
.A(n_1656),
.B(n_1633),
.Y(n_1695)
);

NAND2xp33_ASAP7_75t_SL g1696 ( 
.A(n_1677),
.B(n_1532),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1658),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1624),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1636),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1661),
.B(n_1639),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1655),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1650),
.A2(n_1629),
.B1(n_1620),
.B2(n_1630),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1672),
.B(n_1648),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1650),
.A2(n_1620),
.B1(n_1630),
.B2(n_1643),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1648),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1663),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1660),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1663),
.B(n_1598),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1670),
.B(n_1636),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1664),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1664),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1648),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1666),
.Y(n_1717)
);

NAND2xp67_ASAP7_75t_L g1718 ( 
.A(n_1681),
.B(n_1637),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1666),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1656),
.B(n_1641),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1682),
.B(n_1648),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1598),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1668),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1674),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1674),
.B(n_1619),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1667),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1674),
.B(n_1619),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1685),
.B(n_1631),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1688),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1698),
.B(n_1674),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1718),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1698),
.B(n_1682),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1688),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.B(n_1680),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1693),
.B(n_1667),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1718),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1696),
.B(n_1622),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1709),
.B(n_1716),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.B(n_1680),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1695),
.B(n_1686),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1697),
.B(n_1669),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1710),
.B(n_1669),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1690),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1691),
.B(n_1686),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1709),
.B(n_1654),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1716),
.B(n_1654),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1659),
.Y(n_1752)
);

NAND4xp25_ASAP7_75t_L g1753 ( 
.A(n_1699),
.B(n_1629),
.C(n_1599),
.D(n_1633),
.Y(n_1753)
);

NAND2x1_ASAP7_75t_L g1754 ( 
.A(n_1725),
.B(n_1657),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1690),
.Y(n_1755)
);

INVxp33_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1702),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1707),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1725),
.B(n_1659),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1702),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1657),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1706),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1705),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1720),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

OAI32xp33_ASAP7_75t_L g1767 ( 
.A1(n_1763),
.A2(n_1700),
.A3(n_1689),
.B1(n_1723),
.B2(n_1717),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1732),
.B(n_1720),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1723),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1763),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1737),
.A2(n_1687),
.B1(n_1719),
.B2(n_1717),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1753),
.A2(n_1687),
.B(n_1720),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1737),
.A2(n_1687),
.B1(n_1676),
.B2(n_1645),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1730),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1743),
.B(n_1721),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1753),
.A2(n_1687),
.B(n_1720),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1765),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1741),
.A2(n_1687),
.B1(n_1719),
.B2(n_1726),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

AOI22x1_ASAP7_75t_L g1780 ( 
.A1(n_1738),
.A2(n_1745),
.B1(n_1765),
.B2(n_1761),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1738),
.A2(n_1724),
.B(n_1708),
.Y(n_1781)
);

XOR2x2_ASAP7_75t_L g1782 ( 
.A(n_1749),
.B(n_1677),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1738),
.A2(n_1689),
.B1(n_1700),
.B2(n_1692),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1749),
.B(n_1712),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1743),
.B(n_1752),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1733),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1745),
.A2(n_1728),
.B(n_1726),
.Y(n_1788)
);

AOI322xp5_ASAP7_75t_L g1789 ( 
.A1(n_1733),
.A2(n_1694),
.A3(n_1692),
.B1(n_1701),
.B2(n_1645),
.C1(n_1679),
.C2(n_1728),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1733),
.A2(n_1728),
.B1(n_1726),
.B2(n_1603),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1744),
.B(n_1712),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1777),
.B(n_1758),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1770),
.B(n_1761),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_SL g1794 ( 
.A(n_1770),
.B(n_1758),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1784),
.B(n_1745),
.C(n_1739),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1746),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1766),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1780),
.A2(n_1740),
.B(n_1739),
.Y(n_1799)
);

XNOR2x2_ASAP7_75t_L g1800 ( 
.A(n_1782),
.B(n_1746),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1784),
.B(n_1740),
.C(n_1744),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1786),
.B(n_1750),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1779),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1768),
.B(n_1754),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1782),
.A2(n_1740),
.B1(n_1762),
.B2(n_1760),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1767),
.A2(n_1754),
.B(n_1747),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1771),
.A2(n_1764),
.B1(n_1762),
.B2(n_1755),
.C(n_1760),
.Y(n_1808)
);

OAI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1788),
.A2(n_1789),
.B(n_1776),
.Y(n_1809)
);

OAI21xp33_ASAP7_75t_L g1810 ( 
.A1(n_1772),
.A2(n_1759),
.B(n_1747),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1768),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1792),
.Y(n_1812)
);

AOI31xp33_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1769),
.A3(n_1778),
.B(n_1783),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1807),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_SL g1815 ( 
.A(n_1794),
.B(n_1791),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1802),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1797),
.Y(n_1817)
);

NAND3x1_ASAP7_75t_L g1818 ( 
.A(n_1805),
.B(n_1781),
.C(n_1790),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1798),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1803),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1796),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1808),
.B(n_1750),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1795),
.B(n_1751),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1823),
.B(n_1793),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1815),
.B(n_1799),
.C(n_1801),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1814),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1815),
.B(n_1805),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1812),
.Y(n_1828)
);

OAI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1813),
.A2(n_1809),
.B(n_1810),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1821),
.B(n_1751),
.Y(n_1830)
);

NAND4xp25_ASAP7_75t_SL g1831 ( 
.A(n_1822),
.B(n_1806),
.C(n_1804),
.D(n_1800),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1817),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1816),
.B(n_1799),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1819),
.Y(n_1834)
);

NAND4xp25_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1761),
.C(n_1759),
.D(n_1787),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1825),
.A2(n_1818),
.B(n_1773),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1830),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1827),
.A2(n_1787),
.B1(n_1764),
.B2(n_1757),
.C(n_1755),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1831),
.A2(n_1757),
.B(n_1748),
.Y(n_1839)
);

OAI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1829),
.A2(n_1748),
.B(n_1731),
.C(n_1694),
.Y(n_1840)
);

AOI322xp5_ASAP7_75t_L g1841 ( 
.A1(n_1833),
.A2(n_1701),
.A3(n_1761),
.B1(n_1752),
.B2(n_1751),
.C1(n_1708),
.C2(n_1711),
.Y(n_1841)
);

OAI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1836),
.A2(n_1828),
.B(n_1826),
.C(n_1824),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_SL g1843 ( 
.A1(n_1838),
.A2(n_1834),
.B1(n_1832),
.B2(n_1731),
.Y(n_1843)
);

AOI32xp33_ASAP7_75t_L g1844 ( 
.A1(n_1837),
.A2(n_1835),
.A3(n_1752),
.B1(n_1742),
.B2(n_1735),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1839),
.A2(n_1835),
.B(n_1727),
.Y(n_1845)
);

OA22x2_ASAP7_75t_L g1846 ( 
.A1(n_1840),
.A2(n_1728),
.B1(n_1726),
.B2(n_1742),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1841),
.Y(n_1847)
);

NAND4xp75_ASAP7_75t_L g1848 ( 
.A(n_1847),
.B(n_1735),
.C(n_1734),
.D(n_1626),
.Y(n_1848)
);

AO22x2_ASAP7_75t_L g1849 ( 
.A1(n_1842),
.A2(n_1845),
.B1(n_1843),
.B2(n_1846),
.Y(n_1849)
);

NAND4xp75_ASAP7_75t_L g1850 ( 
.A(n_1844),
.B(n_1734),
.C(n_1626),
.D(n_1727),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1847),
.A2(n_1722),
.B1(n_1715),
.B2(n_1714),
.Y(n_1851)
);

NOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1842),
.B(n_1711),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1848),
.B(n_1851),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1852),
.B(n_1715),
.C(n_1714),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1849),
.B(n_1722),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1853),
.B(n_1850),
.C(n_1657),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1856),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1855),
.B1(n_1854),
.B2(n_1665),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1857),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1859),
.B(n_1657),
.Y(n_1860)
);

AOI22x1_ASAP7_75t_L g1861 ( 
.A1(n_1858),
.A2(n_1729),
.B1(n_1679),
.B2(n_1562),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1860),
.A2(n_1665),
.B1(n_1671),
.B2(n_1729),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1861),
.A2(n_1665),
.B(n_1671),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1863),
.A2(n_1557),
.B1(n_1649),
.B2(n_1644),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1864),
.A2(n_1862),
.B(n_1644),
.Y(n_1865)
);

XNOR2xp5_ASAP7_75t_L g1866 ( 
.A(n_1865),
.B(n_1563),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_R g1867 ( 
.A1(n_1866),
.A2(n_1557),
.B1(n_1647),
.B2(n_1671),
.C(n_1665),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1569),
.B(n_1593),
.C(n_1671),
.Y(n_1868)
);


endmodule