module fake_jpeg_28853_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

BUFx12f_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_31),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_26),
.B1(n_28),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_68),
.B1(n_42),
.B2(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_57),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_66),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_70),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_23),
.B1(n_33),
.B2(n_22),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_74),
.B(n_2),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_30),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_64),
.C(n_48),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_87),
.B1(n_106),
.B2(n_82),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_102),
.B1(n_103),
.B2(n_1),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_20),
.B(n_24),
.C(n_29),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_10),
.B(n_4),
.C(n_5),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_36),
.B1(n_21),
.B2(n_38),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_21),
.B1(n_38),
.B2(n_30),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_104),
.B1(n_108),
.B2(n_72),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_97),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_21),
.B1(n_19),
.B2(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_47),
.A2(n_23),
.B1(n_32),
.B2(n_27),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_59),
.B1(n_57),
.B2(n_56),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_27),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_0),
.Y(n_121)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_53),
.B1(n_58),
.B2(n_61),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_119),
.B1(n_106),
.B2(n_101),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_116),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_118),
.B1(n_107),
.B2(n_75),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_58),
.B1(n_64),
.B2(n_48),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_72),
.B1(n_27),
.B2(n_64),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_138),
.B(n_100),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_74),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_9),
.A3(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_75),
.B1(n_109),
.B2(n_80),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_6),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_6),
.C(n_15),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_87),
.C(n_80),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_103),
.B(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_155),
.B1(n_139),
.B2(n_126),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_156),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_162),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_158),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_76),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_129),
.B1(n_136),
.B2(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_76),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_95),
.B1(n_86),
.B2(n_94),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_93),
.B(n_105),
.C(n_110),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_168),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_109),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_140),
.B1(n_134),
.B2(n_138),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_185),
.B1(n_187),
.B2(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_197),
.B1(n_199),
.B2(n_145),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_134),
.B(n_139),
.C(n_136),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_195),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_99),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_142),
.A2(n_84),
.B1(n_96),
.B2(n_88),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_121),
.C(n_133),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_146),
.C(n_167),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_83),
.B1(n_110),
.B2(n_105),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_83),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_161),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_218),
.B(n_220),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_196),
.B(n_191),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_162),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_215),
.C(n_217),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_169),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_177),
.B1(n_197),
.B2(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_149),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_152),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_164),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_144),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_151),
.C(n_154),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_158),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_144),
.C(n_168),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_188),
.C(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_177),
.B(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_194),
.B1(n_191),
.B2(n_174),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_210),
.B1(n_203),
.B2(n_202),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_194),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_203),
.B1(n_204),
.B2(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_189),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_237),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_141),
.B(n_195),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_141),
.B(n_193),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_238),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_170),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_160),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_208),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_195),
.B1(n_199),
.B2(n_227),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_248),
.B1(n_233),
.B2(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_222),
.B1(n_212),
.B2(n_211),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_195),
.C(n_198),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_207),
.C(n_176),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_226),
.C(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_241),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_236),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_263),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_232),
.B1(n_237),
.B2(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_230),
.B1(n_223),
.B2(n_241),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_265),
.B1(n_246),
.B2(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_195),
.B1(n_206),
.B2(n_159),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_165),
.B1(n_206),
.B2(n_147),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_250),
.B(n_245),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_272),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_260),
.B1(n_249),
.B2(n_258),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_265),
.B1(n_263),
.B2(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

NAND2x1p5_ASAP7_75t_R g277 ( 
.A(n_267),
.B(n_249),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_277),
.A2(n_259),
.B1(n_256),
.B2(n_251),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_282),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_11),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_271),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_279),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_274),
.C(n_275),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_278),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_284),
.B(n_11),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_13),
.B(n_16),
.Y(n_294)
);

OAI21x1_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_293),
.B(n_16),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_2),
.B(n_294),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_296),
.Y(n_297)
);


endmodule