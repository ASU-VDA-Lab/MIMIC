module real_jpeg_1566_n_27 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_147, n_24, n_146, n_6, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_26, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_155, n_27);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_147;
input n_24;
input n_146;
input n_6;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_26;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_66),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_4),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_5),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_6),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_75),
.B1(n_77),
.B2(n_88),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_11),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_13),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_40),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_16),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_17),
.B(n_53),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_74),
.C(n_89),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_20),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_72),
.C(n_97),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_23),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_26),
.A2(n_70),
.B1(n_104),
.B2(n_107),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.C(n_141),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_48),
.Y(n_47)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_36),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_36),
.Y(n_96)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_144),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_140),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_46),
.B(n_49),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_56),
.C(n_139),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_135),
.C(n_136),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_134),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_138),
.Y(n_137)
);

OAI221xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_109),
.C(n_124),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_100),
.C(n_101),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_92),
.C(n_93),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_86),
.C(n_87),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_125),
.A3(n_126),
.B1(n_129),
.B2(n_130),
.C1(n_133),
.C2(n_156),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.C(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_146),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_147),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_148),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_149),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_150),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_151),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_152),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_153),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_154),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_155),
.Y(n_123)
);


endmodule