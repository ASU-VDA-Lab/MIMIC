module fake_jpeg_23633_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_33),
.CON(n_45),
.SN(n_45)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_28),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_7),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_40),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_60),
.B1(n_18),
.B2(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_61),
.B1(n_29),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_20),
.B1(n_18),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_63),
.B1(n_23),
.B2(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_22),
.B1(n_18),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_62),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_38),
.C(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_82),
.C(n_57),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_71),
.B1(n_21),
.B2(n_26),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_84),
.B1(n_48),
.B2(n_53),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_38),
.B1(n_33),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_56),
.B1(n_48),
.B2(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_24),
.B1(n_39),
.B2(n_21),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_50),
.B1(n_16),
.B2(n_27),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_38),
.C(n_33),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_33),
.B1(n_39),
.B2(n_37),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_33),
.A3(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_56),
.B(n_16),
.C(n_44),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_106),
.B1(n_107),
.B2(n_86),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_98),
.B1(n_70),
.B2(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_84),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_82),
.B1(n_84),
.B2(n_65),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_100),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_47),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_0),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_84),
.B1(n_79),
.B2(n_62),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_81),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_111),
.B(n_9),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_123),
.B1(n_130),
.B2(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_105),
.B1(n_102),
.B2(n_77),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_105),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_73),
.B(n_81),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_52),
.B1(n_49),
.B2(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_104),
.B1(n_75),
.B2(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_134),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_147),
.B1(n_153),
.B2(n_122),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_137),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_73),
.C(n_44),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_118),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_95),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_128),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_16),
.B1(n_27),
.B2(n_104),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_16),
.B(n_27),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_8),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_0),
.C(n_1),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_163),
.B1(n_165),
.B2(n_169),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_127),
.B(n_123),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_168),
.B(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_147),
.B1(n_154),
.B2(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_128),
.B1(n_123),
.B2(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_118),
.B1(n_115),
.B2(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_192),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_190),
.B1(n_177),
.B2(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_142),
.C(n_116),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.C(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_116),
.C(n_120),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_121),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_193),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_168),
.B1(n_163),
.B2(n_158),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_188),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_112),
.B1(n_131),
.B2(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_131),
.B1(n_112),
.B2(n_120),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_112),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_160),
.B1(n_167),
.B2(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_120),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_156),
.B(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_156),
.B(n_174),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_177),
.B1(n_193),
.B2(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_171),
.C(n_131),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_1),
.C(n_2),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_182),
.C(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_219),
.C(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_196),
.A2(n_188),
.B1(n_185),
.B2(n_11),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_219),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_7),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_207),
.B1(n_202),
.B2(n_194),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_3),
.C(n_4),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_226),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_227),
.B1(n_224),
.B2(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_204),
.B(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_230),
.B(n_221),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.C(n_212),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_198),
.B(n_6),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_198),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_211),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_6),
.B(n_8),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_12),
.B(n_13),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_246),
.B(n_248),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_232),
.B1(n_231),
.B2(n_13),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_247),
.A2(n_241),
.B(n_242),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_12),
.B(n_14),
.Y(n_253)
);

AOI221xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_4),
.B1(n_12),
.B2(n_14),
.C(n_248),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_254),
.Y(n_255)
);


endmodule