module fake_jpeg_13605_n_40 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_13),
.B(n_11),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_22),
.B1(n_17),
.B2(n_14),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_19),
.B(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_16),
.B(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_27),
.B1(n_25),
.B2(n_4),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.C(n_2),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_36),
.B(n_4),
.Y(n_39)
);

NAND4xp25_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_1),
.C(n_5),
.D(n_6),
.Y(n_40)
);


endmodule