module fake_netlist_1_4880_n_583 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_583);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_583;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_48), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_18), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_8), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_62), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_15), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_13), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_7), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_7), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_56), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_59), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_60), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_32), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_14), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_20), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_47), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_52), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_18), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_50), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_28), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_75), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_65), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_51), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_13), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_17), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_46), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_81), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_76), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_70), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_39), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_25), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_102), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_86), .B(n_0), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_115), .B(n_0), .Y(n_123) );
BUFx8_ASAP7_75t_L g124 ( .A(n_102), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_99), .Y(n_128) );
OAI22x1_ASAP7_75t_R g129 ( .A1(n_82), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_86), .B(n_1), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_99), .B(n_3), .Y(n_132) );
NOR2xp33_ASAP7_75t_SL g133 ( .A(n_113), .B(n_41), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_100), .B(n_4), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_88), .B(n_4), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_84), .A2(n_42), .B(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
OAI22x1_ASAP7_75t_L g142 ( .A1(n_88), .A2(n_5), .B1(n_6), .B2(n_9), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_105), .B(n_113), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_105), .B(n_5), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_143), .B(n_119), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_143), .B(n_98), .Y(n_146) );
NAND3xp33_ASAP7_75t_L g147 ( .A(n_134), .B(n_104), .C(n_93), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_123), .A2(n_115), .B1(n_83), .B2(n_91), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_138), .B(n_119), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_133), .A2(n_117), .B1(n_89), .B2(n_111), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_138), .B(n_87), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_133), .B(n_96), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_123), .B(n_94), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_132), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_124), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_127), .B(n_108), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_127), .B(n_114), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_127), .B(n_110), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_124), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_141), .B(n_112), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_146), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_146), .B(n_122), .Y(n_175) );
AO22x1_ASAP7_75t_L g176 ( .A1(n_148), .A2(n_129), .B1(n_85), .B2(n_134), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_145), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NAND2x1_ASAP7_75t_L g180 ( .A(n_152), .B(n_141), .Y(n_180) );
OR2x6_ASAP7_75t_L g181 ( .A(n_148), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_169), .B(n_130), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_163), .B(n_92), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_169), .B(n_130), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_169), .B(n_135), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_153), .B(n_135), .Y(n_186) );
NOR3x1_ASAP7_75t_L g187 ( .A(n_147), .B(n_129), .C(n_144), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_160), .B(n_144), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_169), .B(n_116), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_157), .B(n_142), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_157), .B(n_124), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_149), .A2(n_141), .B1(n_91), .B2(n_92), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_155), .A2(n_142), .B1(n_91), .B2(n_110), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_155), .B(n_137), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_172), .B(n_124), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_155), .B(n_124), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_161), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_170), .B(n_103), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_156), .B(n_95), .Y(n_205) );
OAI221xp5_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_95), .B1(n_97), .B2(n_101), .C(n_107), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_167), .B(n_97), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_154), .A2(n_101), .B1(n_107), .B2(n_109), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_175), .B(n_158), .Y(n_210) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_183), .A2(n_168), .B(n_171), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_191), .Y(n_212) );
NOR3xp33_ASAP7_75t_L g213 ( .A(n_176), .B(n_109), .C(n_165), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_183), .A2(n_166), .B(n_165), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_173), .B(n_166), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_191), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_166), .B1(n_165), .B2(n_164), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_200), .B(n_166), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_206), .A2(n_106), .B(n_118), .C(n_120), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_208), .A2(n_165), .B1(n_164), .B2(n_118), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_177), .B(n_182), .Y(n_222) );
NOR2x1_ASAP7_75t_L g223 ( .A(n_192), .B(n_164), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_194), .A2(n_120), .B(n_139), .C(n_136), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_184), .B(n_164), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_185), .A2(n_139), .B(n_136), .C(n_159), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_203), .B(n_6), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_200), .B(n_159), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_137), .B(n_151), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_186), .B(n_9), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_186), .B(n_139), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
AO21x1_ASAP7_75t_L g236 ( .A1(n_198), .A2(n_126), .B(n_151), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_200), .B(n_131), .Y(n_237) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_192), .B(n_139), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_188), .B(n_10), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_199), .A2(n_151), .B(n_126), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_192), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_193), .A2(n_126), .B(n_131), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_136), .B(n_131), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_174), .B(n_10), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_214), .A2(n_180), .B(n_197), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_205), .B(n_181), .C(n_188), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_218), .A2(n_202), .B(n_204), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_243), .A2(n_190), .B(n_207), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_245), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_222), .A2(n_209), .B1(n_207), .B2(n_195), .C(n_187), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_222), .B(n_181), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_233), .A2(n_195), .B(n_131), .C(n_125), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_212), .Y(n_255) );
BUFx12f_ASAP7_75t_L g256 ( .A(n_241), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
AOI221x1_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_131), .B1(n_125), .B2(n_121), .C(n_16), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_244), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_210), .B(n_11), .Y(n_260) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_236), .A2(n_131), .A3(n_125), .B(n_121), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_219), .A2(n_131), .B(n_125), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_244), .Y(n_264) );
NAND3xp33_ASAP7_75t_SL g265 ( .A(n_213), .B(n_11), .C(n_12), .Y(n_265) );
AOI21xp5_ASAP7_75t_SL g266 ( .A1(n_235), .A2(n_125), .B(n_121), .Y(n_266) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_236), .A2(n_125), .A3(n_121), .B(n_17), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_239), .B(n_12), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_125), .B1(n_121), .B2(n_14), .Y(n_269) );
O2A1O1Ixp5_ASAP7_75t_L g270 ( .A1(n_219), .A2(n_121), .B(n_23), .C(n_24), .Y(n_270) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_216), .B(n_21), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_27), .B(n_29), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_227), .A2(n_30), .B(n_31), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_237), .A2(n_33), .B(n_34), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_247), .A2(n_229), .B(n_228), .C(n_234), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_258), .A2(n_240), .B(n_237), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_252), .A2(n_225), .B(n_223), .C(n_238), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_253), .B(n_245), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_259), .B(n_230), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_248), .B(n_224), .Y(n_281) );
OAI21x1_ASAP7_75t_SL g282 ( .A1(n_249), .A2(n_221), .B(n_211), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_257), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_274), .Y(n_284) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_231), .B(n_226), .Y(n_285) );
OAI21x1_ASAP7_75t_SL g286 ( .A1(n_275), .A2(n_226), .B(n_235), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_264), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_231), .B(n_235), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_235), .B(n_36), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_261), .Y(n_290) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_250), .A2(n_35), .B(n_37), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_255), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_273), .A2(n_38), .A3(n_40), .B(n_43), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_274), .B(n_44), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_256), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_255), .B(n_80), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_263), .Y(n_297) );
OAI21x1_ASAP7_75t_SL g298 ( .A1(n_271), .A2(n_45), .B(n_49), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_256), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_263), .B(n_53), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
AOI21xp5_ASAP7_75t_SL g302 ( .A1(n_300), .A2(n_271), .B(n_265), .Y(n_302) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_276), .A2(n_268), .B(n_269), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_283), .B(n_267), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_290), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_267), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_282), .A2(n_272), .B(n_260), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_298), .A2(n_251), .B1(n_246), .B2(n_272), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_287), .B(n_267), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_292), .B(n_251), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_281), .B(n_251), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_292), .B(n_267), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_288), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_297), .B(n_261), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_300), .Y(n_321) );
OAI221xp5_ASAP7_75t_SL g322 ( .A1(n_295), .A2(n_266), .B1(n_261), .B2(n_270), .C(n_61), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_277), .A2(n_261), .B(n_266), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_298), .B(n_54), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_320), .B(n_310), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_304), .B(n_297), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_320), .B(n_284), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_304), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_307), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_320), .B(n_284), .Y(n_333) );
NOR2xp67_ASAP7_75t_L g334 ( .A(n_316), .B(n_319), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_309), .B(n_281), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_318), .B(n_289), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_305), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_281), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_306), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_306), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_317), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_314), .B(n_289), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_317), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_318), .B(n_289), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_318), .B(n_293), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_312), .B(n_289), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_293), .Y(n_355) );
AND2x4_ASAP7_75t_SL g356 ( .A(n_350), .B(n_301), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_350), .B(n_312), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_330), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_327), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_329), .B(n_319), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_327), .B(n_316), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_329), .B(n_313), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_331), .B(n_313), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_350), .B(n_313), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_326), .B(n_301), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_331), .B(n_301), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_350), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_333), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_332), .B(n_337), .Y(n_376) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_334), .B(n_324), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_326), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_332), .B(n_301), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_342), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_337), .B(n_324), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_335), .B(n_299), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_328), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_343), .B(n_321), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_343), .B(n_353), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_349), .B(n_321), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_349), .B(n_324), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_335), .A2(n_324), .B1(n_321), .B2(n_303), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_353), .B(n_315), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_339), .B(n_315), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_341), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_344), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_342), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_338), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_352), .Y(n_404) );
NAND2x1_ASAP7_75t_L g405 ( .A(n_377), .B(n_324), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_378), .B(n_339), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_359), .B(n_325), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_398), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_385), .B(n_352), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_366), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_362), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_378), .B(n_284), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_363), .B(n_352), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_363), .B(n_352), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_364), .B(n_351), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_364), .B(n_351), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_382), .B(n_284), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_375), .B(n_346), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_360), .B(n_351), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_365), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_373), .B(n_336), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_373), .B(n_336), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_377), .B(n_334), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_361), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_386), .B(n_336), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_386), .B(n_347), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_361), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_362), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_389), .B(n_346), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_372), .B(n_294), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_374), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_358), .B(n_325), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_390), .B(n_348), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_374), .B(n_348), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_381), .B(n_347), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_399), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_374), .B(n_355), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_379), .B(n_355), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_381), .B(n_355), .Y(n_444) );
AND2x4_ASAP7_75t_SL g445 ( .A(n_381), .B(n_338), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_358), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_396), .B(n_338), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_365), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_396), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_381), .B(n_354), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_383), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_383), .B(n_338), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_391), .B(n_345), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_391), .B(n_354), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_392), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_392), .B(n_354), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_421), .B(n_401), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_426), .B(n_388), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_444), .B(n_387), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_405), .A2(n_413), .B(n_418), .C(n_426), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_402), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_405), .A2(n_388), .B(n_387), .C(n_356), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_403), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_403), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_433), .A2(n_303), .B(n_278), .C(n_280), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_406), .A2(n_387), .B1(n_397), .B2(n_367), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_446), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_427), .B(n_387), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_411), .B(n_302), .C(n_311), .D(n_279), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_407), .B(n_397), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_426), .A2(n_356), .B(n_367), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_407), .B(n_368), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_421), .B(n_401), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_431), .B(n_357), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_404), .B(n_357), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_412), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_404), .B(n_357), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_449), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_368), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_444), .B(n_369), .Y(n_484) );
NAND2x1_ASAP7_75t_SL g485 ( .A(n_434), .B(n_369), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_416), .B(n_380), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_435), .B(n_357), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_434), .B(n_322), .C(n_296), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_434), .B(n_380), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_422), .B(n_400), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_444), .B(n_369), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_437), .B(n_369), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_409), .B(n_371), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_436), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_423), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_422), .B(n_400), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_423), .Y(n_498) );
INVx3_ASAP7_75t_SL g499 ( .A(n_445), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_445), .A2(n_371), .B(n_370), .C(n_322), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_420), .Y(n_501) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_409), .A2(n_370), .B(n_394), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_448), .B(n_395), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_490), .B(n_416), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_462), .B(n_417), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_464), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_460), .A2(n_447), .B1(n_438), .B2(n_432), .C(n_448), .Y(n_508) );
AOI21xp33_ASAP7_75t_SL g509 ( .A1(n_499), .A2(n_447), .B(n_442), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_482), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_465), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_478), .B(n_440), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_501), .B(n_425), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_459), .B(n_450), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_490), .B(n_417), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_481), .B(n_484), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_497), .B(n_424), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_496), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_470), .A2(n_456), .B1(n_454), .B2(n_415), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_479), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_484), .B(n_440), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_491), .Y(n_523) );
AOI32xp33_ASAP7_75t_L g524 ( .A1(n_467), .A2(n_414), .A3(n_415), .B1(n_428), .B2(n_429), .Y(n_524) );
NAND2xp33_ASAP7_75t_L g525 ( .A(n_463), .B(n_414), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_493), .B(n_428), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_498), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_495), .B(n_455), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_500), .A2(n_455), .B(n_451), .C(n_452), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_470), .A2(n_429), .B(n_450), .C(n_424), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_458), .A2(n_439), .B(n_442), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_468), .Y(n_532) );
O2A1O1Ixp5_ASAP7_75t_L g533 ( .A1(n_477), .A2(n_442), .B(n_439), .C(n_451), .Y(n_533) );
AOI321xp33_ASAP7_75t_SL g534 ( .A1(n_487), .A2(n_425), .A3(n_439), .B1(n_293), .B2(n_453), .C(n_419), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_457), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_505), .B(n_497), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_535), .B(n_472), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_519), .A2(n_466), .B(n_473), .C(n_488), .Y(n_538) );
XNOR2x2_ASAP7_75t_L g539 ( .A(n_508), .B(n_474), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_530), .A2(n_491), .B1(n_459), .B2(n_469), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_525), .A2(n_502), .B1(n_492), .B2(n_494), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_510), .B(n_476), .Y(n_542) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_508), .A2(n_483), .A3(n_475), .B1(n_486), .B2(n_457), .C1(n_476), .C2(n_503), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g544 ( .A1(n_530), .A2(n_489), .B(n_503), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_529), .A2(n_480), .B(n_410), .C(n_441), .Y(n_545) );
OAI321xp33_ASAP7_75t_L g546 ( .A1(n_534), .A2(n_408), .A3(n_441), .B1(n_419), .B2(n_410), .C(n_394), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_528), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_524), .A2(n_485), .B1(n_395), .B2(n_393), .C(n_323), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_531), .A2(n_393), .B1(n_308), .B2(n_323), .Y(n_549) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_521), .Y(n_550) );
AOI21xp33_ASAP7_75t_L g551 ( .A1(n_533), .A2(n_308), .B(n_323), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_528), .Y(n_552) );
AO22x1_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_323), .B1(n_293), .B2(n_308), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_513), .B(n_308), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g555 ( .A1(n_509), .A2(n_277), .B(n_293), .C(n_291), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_506), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_532), .A2(n_323), .B1(n_291), .B2(n_285), .C(n_293), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_523), .A2(n_282), .B1(n_286), .B2(n_285), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_506), .A2(n_286), .B1(n_57), .B2(n_63), .C(n_66), .Y(n_559) );
NAND3xp33_ASAP7_75t_SL g560 ( .A(n_515), .B(n_55), .C(n_67), .Y(n_560) );
AOI21xp33_ASAP7_75t_SL g561 ( .A1(n_514), .A2(n_68), .B(n_69), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_504), .B(n_71), .Y(n_562) );
AOI322xp5_ASAP7_75t_L g563 ( .A1(n_526), .A2(n_72), .A3(n_73), .B1(n_74), .B2(n_77), .C1(n_78), .C2(n_522), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_517), .B(n_526), .C(n_516), .Y(n_564) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_560), .B(n_562), .Y(n_565) );
NAND4xp25_ASAP7_75t_L g566 ( .A(n_538), .B(n_540), .C(n_563), .D(n_548), .Y(n_566) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_541), .B(n_539), .C(n_544), .D(n_559), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_550), .A2(n_561), .B(n_549), .C(n_564), .Y(n_568) );
OAI211xp5_ASAP7_75t_SL g569 ( .A1(n_545), .A2(n_554), .B(n_546), .C(n_555), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_552), .B(n_547), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_567), .B(n_551), .C(n_558), .D(n_546), .Y(n_571) );
NOR4xp25_ASAP7_75t_L g572 ( .A(n_568), .B(n_543), .C(n_542), .D(n_556), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_570), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_573), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_571), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_574), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_575), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_566), .B1(n_572), .B2(n_565), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_578), .A2(n_576), .B1(n_536), .B2(n_537), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_579), .A2(n_569), .B(n_553), .Y(n_580) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_520), .B(n_511), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_581), .A2(n_507), .B(n_518), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_512), .B1(n_527), .B2(n_557), .Y(n_583) );
endmodule