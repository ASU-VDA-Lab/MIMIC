module fake_jpeg_1507_n_650 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_553;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g202 ( 
.A(n_58),
.Y(n_202)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_60),
.B(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_68),
.B(n_72),
.Y(n_165)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_74),
.Y(n_214)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_77),
.B(n_83),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_87),
.B(n_94),
.Y(n_178)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_36),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_100),
.B(n_107),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_102),
.Y(n_137)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_37),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_36),
.A2(n_16),
.B1(n_15),
.B2(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_109),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_28),
.B(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_32),
.Y(n_155)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_37),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_115),
.B(n_118),
.Y(n_225)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_27),
.B(n_16),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_39),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_121),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_48),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_53),
.Y(n_170)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_126),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_55),
.B(n_53),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_131),
.B(n_170),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_132),
.B(n_135),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_67),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_138),
.B(n_145),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_84),
.B(n_31),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_92),
.B(n_32),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_148),
.B(n_152),
.Y(n_244)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_78),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_153),
.B(n_201),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_174),
.Y(n_228)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_55),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_89),
.B(n_52),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_175),
.B(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_52),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_66),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_177),
.B(n_182),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_102),
.Y(n_182)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_187),
.A2(n_10),
.B1(n_12),
.B2(n_225),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_50),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_215),
.Y(n_252)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_119),
.A2(n_120),
.B1(n_90),
.B2(n_105),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_199),
.A2(n_47),
.B1(n_41),
.B2(n_44),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_126),
.A2(n_58),
.B(n_122),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_90),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_205),
.B(n_217),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_58),
.Y(n_212)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_65),
.B(n_50),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_80),
.B(n_30),
.Y(n_217)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_79),
.Y(n_218)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g222 ( 
.A(n_74),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_82),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_3),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_44),
.B1(n_39),
.B2(n_49),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_231),
.A2(n_237),
.B1(n_238),
.B2(n_253),
.Y(n_320)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_236),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_130),
.A2(n_81),
.B1(n_103),
.B2(n_47),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_130),
.A2(n_47),
.B1(n_41),
.B2(n_30),
.Y(n_238)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_139),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_246),
.B(n_258),
.Y(n_331)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_133),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_247),
.Y(n_330)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_184),
.A2(n_47),
.B1(n_41),
.B2(n_44),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_249),
.A2(n_264),
.B1(n_277),
.B2(n_281),
.Y(n_315)
);

CKINVDCx12_ASAP7_75t_R g250 ( 
.A(n_140),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_163),
.Y(n_254)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_254),
.Y(n_353)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_202),
.A2(n_34),
.B1(n_42),
.B2(n_49),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_266),
.Y(n_327)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_168),
.B(n_34),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_197),
.A2(n_49),
.B1(n_44),
.B2(n_127),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_167),
.A2(n_49),
.B1(n_74),
.B2(n_85),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_178),
.Y(n_262)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_124),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_168),
.B(n_2),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_268),
.B(n_280),
.Y(n_346)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_143),
.Y(n_270)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_272),
.Y(n_369)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_143),
.Y(n_273)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_276),
.A2(n_284),
.B1(n_285),
.B2(n_200),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_183),
.Y(n_279)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_180),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_154),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_199),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_212),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_157),
.A2(n_191),
.B1(n_170),
.B2(n_190),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_164),
.Y(n_286)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_140),
.B(n_7),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_290),
.Y(n_355)
);

CKINVDCx12_ASAP7_75t_R g288 ( 
.A(n_165),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_134),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_179),
.Y(n_291)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_188),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_293),
.A2(n_298),
.B1(n_301),
.B2(n_149),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_165),
.B(n_208),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_299),
.Y(n_363)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_146),
.Y(n_296)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_159),
.Y(n_297)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_134),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_144),
.Y(n_300)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_196),
.A2(n_12),
.B1(n_206),
.B2(n_136),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_141),
.B(n_142),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_302),
.B(n_307),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_204),
.Y(n_321)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_129),
.Y(n_304)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_154),
.Y(n_305)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_137),
.Y(n_306)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_306),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_150),
.B(n_147),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_181),
.Y(n_308)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_158),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_309),
.B(n_207),
.Y(n_352)
);

AO22x2_ASAP7_75t_SL g310 ( 
.A1(n_241),
.A2(n_193),
.B1(n_160),
.B2(n_161),
.Y(n_310)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_240),
.B(n_211),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_335),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_321),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_322),
.A2(n_341),
.B1(n_366),
.B2(n_229),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_241),
.B(n_173),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_340),
.C(n_308),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_203),
.Y(n_329)
);

NAND2x1_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_344),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_252),
.B(n_181),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_230),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_337),
.B(n_273),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_195),
.C(n_219),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_228),
.A2(n_244),
.B1(n_249),
.B2(n_238),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_274),
.A2(n_214),
.B(n_200),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_343),
.A2(n_350),
.B(n_266),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_185),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_345),
.A2(n_361),
.B1(n_260),
.B2(n_209),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_162),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_362),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_285),
.A2(n_223),
.B(n_210),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_283),
.A2(n_169),
.B1(n_186),
.B2(n_193),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_239),
.B(n_169),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_256),
.A2(n_186),
.B1(n_209),
.B2(n_166),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_370),
.B(n_410),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_320),
.A2(n_237),
.B1(n_264),
.B2(n_301),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_371),
.A2(n_405),
.B1(n_407),
.B2(n_408),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_316),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_372),
.B(n_381),
.Y(n_426)
);

INVx11_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_373),
.A2(n_382),
.B1(n_393),
.B2(n_400),
.Y(n_439)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_281),
.B(n_293),
.C(n_276),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_375),
.B(n_383),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_377),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_358),
.Y(n_381)
);

INVx13_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_236),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_384),
.Y(n_420)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_321),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_386),
.B(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_388),
.A2(n_330),
.B1(n_367),
.B2(n_328),
.Y(n_428)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_321),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_395),
.A2(n_403),
.B(n_379),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_251),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_406),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_371),
.B1(n_392),
.B2(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

INVx11_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_325),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_325),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_412),
.Y(n_443)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_327),
.A2(n_226),
.B1(n_235),
.B2(n_282),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_312),
.B(n_289),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_L g407 ( 
.A1(n_310),
.A2(n_232),
.B1(n_242),
.B2(n_227),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_324),
.A2(n_359),
.B1(n_310),
.B2(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_323),
.B(n_275),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_346),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_356),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_363),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_360),
.B(n_369),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_413),
.B(n_414),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_270),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_368),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_315),
.B1(n_350),
.B2(n_343),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_421),
.A2(n_428),
.B1(n_448),
.B2(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_397),
.C(n_402),
.Y(n_478)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_354),
.B(n_326),
.C(n_333),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_425),
.A2(n_431),
.B(n_436),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_380),
.A2(n_329),
.B(n_331),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_429),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_330),
.B(n_326),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_378),
.B(n_329),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_433),
.B(n_415),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_344),
.B1(n_328),
.B2(n_311),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_447),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_378),
.A2(n_344),
.B(n_354),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_403),
.A2(n_375),
.B(n_408),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_437),
.B(n_440),
.Y(n_485)
);

AND2x2_ASAP7_75t_SL g440 ( 
.A(n_396),
.B(n_365),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_384),
.A2(n_311),
.B1(n_357),
.B2(n_226),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_407),
.A2(n_357),
.B1(n_367),
.B2(n_333),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_455),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_406),
.Y(n_450)
);

INVx13_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_454),
.B(n_411),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_391),
.A2(n_235),
.B1(n_305),
.B2(n_243),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_451),
.B(n_412),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_457),
.B(n_463),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_391),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_458),
.B(n_478),
.C(n_483),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_445),
.Y(n_459)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

AND2x2_ASAP7_75t_SL g462 ( 
.A(n_444),
.B(n_456),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_462),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_397),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_464),
.B(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_422),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_467),
.B(n_469),
.Y(n_509)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_451),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_484),
.Y(n_505)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_471),
.B(n_474),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_437),
.A2(n_383),
.B1(n_405),
.B2(n_385),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_419),
.B1(n_435),
.B2(n_429),
.Y(n_500)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_374),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_475),
.B(n_477),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_401),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_454),
.B(n_365),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_479),
.B(n_420),
.Y(n_506)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_482),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_440),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_433),
.B(n_397),
.C(n_381),
.Y(n_483)
);

AOI322xp5_ASAP7_75t_L g484 ( 
.A1(n_446),
.A2(n_372),
.A3(n_376),
.B1(n_387),
.B2(n_390),
.C1(n_409),
.C2(n_389),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_488),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_399),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_441),
.Y(n_518)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_493),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_434),
.Y(n_503)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_476),
.A2(n_418),
.B(n_446),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_502),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_489),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_504),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_498),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_421),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_499),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_500),
.A2(n_506),
.B1(n_520),
.B2(n_524),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_491),
.Y(n_501)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_476),
.A2(n_485),
.B(n_487),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_503),
.B(n_490),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_485),
.A2(n_425),
.B(n_434),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_462),
.A2(n_419),
.B1(n_420),
.B2(n_444),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_525),
.B1(n_465),
.B2(n_488),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_478),
.B(n_436),
.C(n_440),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_483),
.C(n_458),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_460),
.B(n_461),
.Y(n_516)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_487),
.B(n_453),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_517),
.B(n_516),
.Y(n_543)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_518),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_470),
.A2(n_448),
.B1(n_455),
.B2(n_425),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_485),
.A2(n_431),
.B(n_439),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_465),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_464),
.Y(n_523)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_523),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_472),
.A2(n_447),
.B1(n_432),
.B2(n_441),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_462),
.A2(n_453),
.B1(n_438),
.B2(n_445),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_482),
.A2(n_438),
.B1(n_452),
.B2(n_449),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_526),
.A2(n_400),
.B1(n_373),
.B2(n_271),
.Y(n_555)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_533),
.B(n_556),
.Y(n_577)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_534),
.Y(n_572)
);

HB1xp67_ASAP7_75t_SL g536 ( 
.A(n_499),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g565 ( 
.A(n_536),
.Y(n_565)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_514),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_500),
.A2(n_473),
.B1(n_480),
.B2(n_471),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_545),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_543),
.A2(n_550),
.B1(n_552),
.B2(n_553),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_473),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_544),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_508),
.A2(n_480),
.B1(n_467),
.B2(n_481),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_492),
.C(n_493),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_551),
.C(n_502),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_547),
.B(n_549),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_503),
.B(n_486),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_508),
.A2(n_474),
.B1(n_469),
.B2(n_466),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_496),
.B(n_314),
.C(n_416),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_499),
.A2(n_442),
.B1(n_284),
.B2(n_404),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_507),
.A2(n_442),
.B1(n_376),
.B2(n_314),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_555),
.A2(n_557),
.B1(n_520),
.B2(n_538),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_512),
.B(n_513),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_524),
.A2(n_227),
.B1(n_242),
.B2(n_351),
.Y(n_557)
);

XNOR2x1_ASAP7_75t_L g590 ( 
.A(n_558),
.B(n_547),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_549),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_526),
.C(n_501),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_560),
.B(n_568),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_537),
.A2(n_494),
.B(n_504),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_561),
.A2(n_564),
.B(n_540),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_540),
.A2(n_498),
.B(n_523),
.Y(n_564)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_567),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_512),
.C(n_513),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_495),
.B1(n_527),
.B2(n_506),
.Y(n_569)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_569),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_535),
.A2(n_495),
.B1(n_527),
.B2(n_522),
.Y(n_570)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_570),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_548),
.A2(n_522),
.B1(n_519),
.B2(n_505),
.Y(n_571)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_571),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_533),
.B(n_525),
.C(n_519),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_579),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_529),
.A2(n_518),
.B1(n_517),
.B2(n_515),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_578),
.A2(n_556),
.B1(n_542),
.B2(n_544),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_521),
.C(n_511),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_530),
.B(n_511),
.C(n_515),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_532),
.C(n_545),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_577),
.B(n_534),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_581),
.B(n_585),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_541),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_SL g604 ( 
.A(n_584),
.B(n_591),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_572),
.A2(n_529),
.B1(n_554),
.B2(n_531),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_574),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_586),
.B(n_594),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_590),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_592),
.A2(n_563),
.B1(n_572),
.B2(n_573),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_561),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_577),
.B(n_510),
.Y(n_594)
);

AOI321xp33_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_510),
.A3(n_528),
.B1(n_550),
.B2(n_552),
.C(n_377),
.Y(n_595)
);

INVx11_ASAP7_75t_L g605 ( 
.A(n_595),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_559),
.B(n_553),
.C(n_557),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_596),
.B(n_597),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_528),
.C(n_364),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_598),
.B(n_560),
.C(n_580),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_601),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_597),
.B(n_599),
.C(n_596),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_602),
.A2(n_603),
.B1(n_336),
.B2(n_313),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_583),
.A2(n_573),
.B1(n_563),
.B2(n_566),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_558),
.C(n_566),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_607),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_579),
.C(n_574),
.Y(n_607)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

OA21x2_ASAP7_75t_L g612 ( 
.A1(n_588),
.A2(n_562),
.B(n_578),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_233),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_576),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_613),
.B(n_356),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_565),
.C(n_576),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_317),
.Y(n_626)
);

AOI21xp33_ASAP7_75t_L g616 ( 
.A1(n_610),
.A2(n_587),
.B(n_589),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_617),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_586),
.C(n_590),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_592),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_619),
.B(n_621),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_615),
.A2(n_382),
.B1(n_368),
.B2(n_351),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_620),
.A2(n_605),
.B1(n_614),
.B2(n_609),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_313),
.C(n_317),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_606),
.C(n_607),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_623),
.A2(n_624),
.B1(n_612),
.B2(n_608),
.Y(n_628)
);

INVx11_ASAP7_75t_L g630 ( 
.A(n_626),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_628),
.A2(n_633),
.B1(n_629),
.B2(n_634),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_629),
.B(n_632),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_612),
.C(n_604),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_627),
.A2(n_605),
.B(n_609),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_635),
.A2(n_622),
.B(n_620),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_631),
.A2(n_623),
.B(n_625),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_637),
.B(n_639),
.Y(n_643)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_617),
.Y(n_638)
);

OAI21x1_ASAP7_75t_SL g642 ( 
.A1(n_638),
.A2(n_640),
.B(n_630),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_628),
.C(n_630),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_641),
.B(n_642),
.C(n_279),
.Y(n_644)
);

A2O1A1O1Ixp25_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_645),
.B(n_292),
.C(n_303),
.D(n_348),
.Y(n_646)
);

AOI322xp5_ASAP7_75t_L g645 ( 
.A1(n_643),
.A2(n_393),
.A3(n_303),
.B1(n_292),
.B2(n_233),
.C1(n_263),
.C2(n_348),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_263),
.C(n_292),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_647),
.B(n_353),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_353),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_SL g650 ( 
.A(n_649),
.B(n_172),
.Y(n_650)
);


endmodule