module fake_jpeg_27159_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_46),
.CON(n_51),
.SN(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_26),
.B1(n_27),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_62),
.B1(n_74),
.B2(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_27),
.B1(n_17),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_75),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_22),
.B1(n_21),
.B2(n_16),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_32),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_22),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_93),
.C(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_97),
.B1(n_47),
.B2(n_58),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_53),
.B1(n_7),
.B2(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_33),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_0),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_106),
.B1(n_107),
.B2(n_8),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_0),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_104),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_32),
.C(n_2),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_3),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_4),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_53),
.B(n_49),
.C(n_48),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_122),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_120),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_136),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_85),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_47),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_13),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_96),
.Y(n_126)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_14),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_138),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_7),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_133),
.B(n_109),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_139),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_66),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_66),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_144),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_15),
.C(n_109),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_91),
.C(n_83),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_164),
.C(n_133),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_160),
.B1(n_159),
.B2(n_121),
.C(n_158),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_98),
.B(n_97),
.C(n_82),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_160),
.B(n_132),
.Y(n_179)
);

OR2x4_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_83),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_91),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_15),
.C(n_82),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_79),
.C(n_94),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_81),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_170),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_134),
.B1(n_110),
.B2(n_121),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_174),
.B1(n_133),
.B2(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_173),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_110),
.B(n_138),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_158),
.B(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_136),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_116),
.B1(n_94),
.B2(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_127),
.B1(n_81),
.B2(n_131),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_180),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_184),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_119),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_164),
.C(n_141),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_151),
.A3(n_147),
.B1(n_140),
.B2(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_196),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_145),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_154),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_187),
.B1(n_172),
.B2(n_184),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_146),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_174),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_185),
.B1(n_175),
.B2(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_210),
.B1(n_213),
.B2(n_207),
.Y(n_222)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_168),
.B1(n_171),
.B2(n_182),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_189),
.C(n_192),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_182),
.B1(n_177),
.B2(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_197),
.B1(n_186),
.B2(n_200),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_202),
.Y(n_219)
);

OA21x2_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_201),
.B(n_192),
.Y(n_220)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_220),
.A2(n_204),
.B(n_205),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_223),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_215),
.B(n_203),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_225),
.B(n_224),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_217),
.Y(n_234)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_228),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_224),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_229),
.B(n_227),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_242),
.A3(n_235),
.B1(n_238),
.B2(n_243),
.C1(n_231),
.C2(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_210),
.Y(n_248)
);


endmodule