module fake_jpeg_1263_n_54 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_13),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_25),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_16),
.B(n_17),
.C(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_29),
.C(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_11),
.C(n_10),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_24),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_43),
.B(n_44),
.C(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_0),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_17),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_38),
.C(n_12),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_48),
.C(n_5),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_43),
.A3(n_6),
.B1(n_7),
.B2(n_5),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.C(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_9),
.C(n_6),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_7),
.Y(n_54)
);


endmodule