module fake_ibex_1385_n_578 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_578);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_578;

wire n_151;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_86;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_545;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_88;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_89;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_543;
wire n_483;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_98;
wire n_267;
wire n_245;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_553;
wire n_554;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_365;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_444;
wire n_546;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_238;
wire n_214;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_202;
wire n_159;
wire n_298;
wire n_231;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

BUFx8_ASAP7_75t_SL g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_36),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_12),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_51),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_17),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_56),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_21),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_41),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_54),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_40),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_42),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_18),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_0),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_10),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_25),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

OAI22x1_ASAP7_75t_R g158 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_39),
.B(n_82),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_6),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_87),
.A2(n_47),
.B(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_27),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_28),
.B(n_29),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_30),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_97),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_127),
.A2(n_38),
.B(n_49),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_126),
.A2(n_149),
.B(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_115),
.B(n_52),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_112),
.C(n_129),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

CKINVDCx6p67_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_98),
.B1(n_97),
.B2(n_148),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_165),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_204),
.Y(n_223)
);

OR2x6_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_155),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_191),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_98),
.B1(n_148),
.B2(n_93),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

CKINVDCx11_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_153),
.B(n_90),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_193),
.B(n_90),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_170),
.B(n_124),
.Y(n_239)
);

CKINVDCx6p67_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_166),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx6p67_ASAP7_75t_R g253 ( 
.A(n_166),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_201),
.B(n_138),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

OR2x6_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_136),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_173),
.B(n_135),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_162),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_188),
.B(n_184),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_162),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_188),
.B(n_128),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_201),
.B(n_118),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_181),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_263),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_206),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_230),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_257),
.B(n_111),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_176),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

OAI22x1_ASAP7_75t_R g287 ( 
.A1(n_224),
.A2(n_174),
.B1(n_158),
.B2(n_163),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_176),
.B(n_175),
.C(n_192),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_180),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_180),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_210),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_238),
.B(n_208),
.Y(n_294)
);

BUFx6f_ASAP7_75t_SL g295 ( 
.A(n_224),
.Y(n_295)
);

BUFx6f_ASAP7_75t_SL g296 ( 
.A(n_224),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_192),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_215),
.B(n_225),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_213),
.Y(n_299)
);

OR2x2_ASAP7_75t_SL g300 ( 
.A(n_210),
.B(n_158),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_246),
.B(n_101),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_211),
.A2(n_161),
.B(n_198),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

OR2x6_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_168),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_L g305 ( 
.A(n_209),
.B(n_175),
.C(n_192),
.Y(n_305)
);

NAND2x1_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_190),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_219),
.B(n_179),
.Y(n_307)
);

O2A1O1Ixp5_ASAP7_75t_L g308 ( 
.A1(n_214),
.A2(n_185),
.B(n_179),
.C(n_196),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_239),
.B(n_185),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_234),
.Y(n_311)
);

NOR2x1p5_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_163),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_167),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_214),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_228),
.B(n_167),
.C(n_169),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_260),
.A2(n_217),
.B(n_218),
.C(n_276),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_171),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_221),
.B(n_169),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_217),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_223),
.B(n_151),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_212),
.B(n_151),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_240),
.B(n_154),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_218),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_235),
.B(n_202),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_245),
.A2(n_157),
.B1(n_159),
.B2(n_199),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_161),
.B(n_183),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_198),
.B(n_168),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_200),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_316),
.B(n_308),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_200),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_200),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_313),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_198),
.B(n_183),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_199),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_203),
.B1(n_199),
.B2(n_272),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_203),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_289),
.A2(n_232),
.B(n_233),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_254),
.B1(n_262),
.B2(n_272),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_280),
.A2(n_254),
.B(n_262),
.C(n_266),
.Y(n_344)
);

CKINVDCx10_ASAP7_75t_R g345 ( 
.A(n_281),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_247),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_256),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_259),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_259),
.B(n_222),
.C(n_227),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_264),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_294),
.A2(n_271),
.B(n_274),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_231),
.B(n_269),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g356 ( 
.A1(n_287),
.A2(n_229),
.B1(n_265),
.B2(n_261),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_229),
.B(n_265),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_60),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_61),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_309),
.B(n_64),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_320),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_288),
.A2(n_237),
.B(n_251),
.C(n_250),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_305),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_295),
.A2(n_241),
.B1(n_251),
.B2(n_250),
.Y(n_365)
);

AO21x1_ASAP7_75t_L g366 ( 
.A1(n_315),
.A2(n_216),
.B(n_248),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_296),
.A2(n_226),
.B1(n_244),
.B2(n_243),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_300),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_68),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_284),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_R g376 ( 
.A(n_342),
.B(n_71),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_324),
.Y(n_377)
);

CKINVDCx11_ASAP7_75t_R g378 ( 
.A(n_370),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_348),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_292),
.Y(n_383)
);

NAND2x1p5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_249),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_368),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_355),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_340),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_354),
.Y(n_390)
);

AND3x1_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_358),
.C(n_359),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_349),
.A2(n_360),
.B(n_343),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_338),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

AO31x2_ASAP7_75t_L g396 ( 
.A1(n_366),
.A2(n_344),
.A3(n_350),
.B(n_362),
.Y(n_396)
);

AO31x2_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_341),
.A3(n_372),
.B(n_352),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_367),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_242),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_334),
.B(n_242),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_342),
.Y(n_403)
);

AO31x2_ASAP7_75t_L g404 ( 
.A1(n_366),
.A2(n_330),
.A3(n_337),
.B(n_328),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_347),
.B(n_242),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_326),
.A2(n_357),
.B(n_353),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_326),
.A2(n_357),
.B(n_353),
.Y(n_408)
);

AO31x2_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_330),
.A3(n_337),
.B(n_328),
.Y(n_409)
);

INVx3_ASAP7_75t_SL g410 ( 
.A(n_369),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_326),
.A2(n_357),
.B(n_353),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_334),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_242),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_334),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

NAND2x1p5_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_291),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_345),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_334),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_334),
.B(n_291),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

AO21x2_ASAP7_75t_L g427 ( 
.A1(n_337),
.A2(n_330),
.B(n_328),
.Y(n_427)
);

NOR2x1_ASAP7_75t_SL g428 ( 
.A(n_347),
.B(n_291),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_422),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_403),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_379),
.B(n_423),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_407),
.A2(n_408),
.B(n_411),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_416),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_378),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_376),
.Y(n_440)
);

OR2x6_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_389),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_386),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_391),
.B(n_384),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_414),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_392),
.A2(n_393),
.B(n_394),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_386),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_380),
.A2(n_375),
.B(n_387),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_429),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_381),
.A2(n_390),
.B(n_400),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_381),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_SL g463 ( 
.A1(n_412),
.A2(n_417),
.B(n_418),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_398),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_427),
.A2(n_409),
.B(n_404),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_409),
.A2(n_382),
.B(n_395),
.Y(n_468)
);

CKINVDCx6p67_ASAP7_75t_R g469 ( 
.A(n_410),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_396),
.A2(n_397),
.B(n_377),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_401),
.B(n_406),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_458),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_436),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_460),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_461),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_450),
.B(n_453),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_468),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_438),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_472),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_470),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_459),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_438),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_496),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_475),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_467),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_494),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_481),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_481),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_467),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_467),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_475),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_440),
.C(n_463),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_478),
.A2(n_459),
.B1(n_440),
.B2(n_458),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_499),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_500),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_510),
.A2(n_493),
.B1(n_482),
.B2(n_495),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_511),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_494),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_479),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_488),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_488),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_501),
.Y(n_522)
);

NAND4xp25_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_508),
.C(n_432),
.D(n_510),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_502),
.Y(n_524)
);

NOR3xp33_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_508),
.C(n_430),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_512),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_502),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_513),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_506),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_509),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_528),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_521),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_519),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_519),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_525),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_523),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_533),
.A2(n_503),
.B1(n_504),
.B2(n_509),
.Y(n_541)
);

OAI322xp33_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_531),
.A3(n_529),
.B1(n_524),
.B2(n_505),
.C1(n_484),
.C2(n_474),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_533),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_538),
.A2(n_529),
.B1(n_521),
.B2(n_504),
.Y(n_544)
);

AOI221xp5_ASAP7_75t_L g545 ( 
.A1(n_534),
.A2(n_537),
.B1(n_536),
.B2(n_535),
.C(n_532),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_514),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_506),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_437),
.Y(n_548)
);

AOI221xp5_ASAP7_75t_L g549 ( 
.A1(n_542),
.A2(n_532),
.B1(n_446),
.B2(n_431),
.C(n_493),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_543),
.A2(n_509),
.B1(n_511),
.B2(n_458),
.Y(n_550)
);

OAI211xp5_ASAP7_75t_L g551 ( 
.A1(n_544),
.A2(n_509),
.B(n_511),
.C(n_483),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_545),
.C(n_546),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_541),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_550),
.B(n_469),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_552),
.B(n_469),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_SL g556 ( 
.A(n_553),
.B(n_551),
.C(n_547),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_555),
.B(n_490),
.Y(n_557)
);

NAND4xp25_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_554),
.C(n_442),
.D(n_449),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_558),
.B(n_505),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_557),
.A2(n_490),
.B(n_497),
.Y(n_560)
);

AND3x2_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_471),
.C(n_433),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_497),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_561),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_562),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_564),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_452),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_564),
.Y(n_567)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_563),
.A2(n_441),
.B(n_486),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_566),
.A2(n_441),
.B(n_444),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_486),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_567),
.A2(n_509),
.B1(n_485),
.B2(n_483),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_568),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_570),
.B1(n_571),
.B2(n_569),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_441),
.B(n_487),
.Y(n_574)
);

AO22x1_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_509),
.B1(n_487),
.B2(n_462),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_468),
.B(n_444),
.Y(n_576)
);

OA22x2_ASAP7_75t_L g577 ( 
.A1(n_575),
.A2(n_477),
.B1(n_482),
.B2(n_492),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_576),
.B1(n_509),
.B2(n_477),
.Y(n_578)
);


endmodule