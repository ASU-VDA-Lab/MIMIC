module fake_jpeg_19838_n_205 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_27),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_10),
.Y(n_30)
);

NAND2xp67_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_21),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_52),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_31),
.B(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_54),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_37),
.B1(n_18),
.B2(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_34),
.B1(n_35),
.B2(n_11),
.Y(n_67)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_38),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_34),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_44),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_31),
.A3(n_34),
.B1(n_22),
.B2(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_61),
.B1(n_56),
.B2(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_53),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_43),
.B(n_48),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_45),
.B1(n_47),
.B2(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_59),
.B1(n_67),
.B2(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_47),
.B1(n_46),
.B2(n_49),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_67),
.B1(n_58),
.B2(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_81),
.B1(n_73),
.B2(n_74),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_79),
.C(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_21),
.Y(n_116)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_65),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_77),
.C(n_62),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_113),
.C(n_105),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_110),
.B1(n_95),
.B2(n_89),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_72),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_114),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_74),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_9),
.B(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_57),
.B1(n_63),
.B2(n_83),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_63),
.B(n_83),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_11),
.B(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_66),
.C(n_49),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_49),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_51),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_92),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_51),
.B(n_46),
.C(n_11),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_95),
.B1(n_96),
.B2(n_89),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_124),
.B1(n_135),
.B2(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_21),
.C(n_15),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_113),
.C(n_106),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_21),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_9),
.C(n_18),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_138),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_38),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_86),
.B1(n_9),
.B2(n_12),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_119),
.B(n_106),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_132),
.B(n_137),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_120),
.B1(n_122),
.B2(n_138),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_114),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_153),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_127),
.B1(n_130),
.B2(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_149),
.C(n_151),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_111),
.C(n_21),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_17),
.C(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_131),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_17),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_129),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_134),
.B(n_38),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_3),
.B(n_4),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_17),
.C(n_15),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_149),
.C(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_144),
.C(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_174),
.C(n_163),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_141),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_157),
.C(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_166),
.C(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_155),
.B1(n_165),
.B2(n_5),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_180),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_181),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_179),
.B(n_4),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_17),
.C(n_15),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_190),
.Y(n_193)
);

AOI321xp33_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_186),
.A3(n_15),
.B1(n_12),
.B2(n_7),
.C(n_4),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_5),
.B(n_6),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.C(n_8),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_3),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_6),
.B(n_8),
.C(n_26),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_192),
.C(n_26),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_201),
.B(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_8),
.Y(n_205)
);


endmodule