module fake_jpeg_10167_n_311 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_26),
.B(n_17),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_62),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_49),
.B1(n_31),
.B2(n_33),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_17),
.B2(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_58),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_60),
.B2(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_19),
.B1(n_35),
.B2(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_29),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_18),
.B1(n_35),
.B2(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_29),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_38),
.B(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_35),
.B2(n_20),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_66),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR4xp25_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_9),
.C(n_16),
.D(n_15),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_87),
.C(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_84),
.Y(n_126)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_45),
.B(n_33),
.C(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_49),
.B1(n_67),
.B2(n_106),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_44),
.B1(n_25),
.B2(n_24),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_103),
.B1(n_90),
.B2(n_104),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_28),
.B1(n_20),
.B2(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_18),
.B1(n_20),
.B2(n_32),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_32),
.B1(n_30),
.B2(n_21),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_36),
.CI(n_34),
.CON(n_100),
.SN(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_63),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_106),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_44),
.B1(n_21),
.B2(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_22),
.Y(n_133)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_102),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_136),
.B1(n_81),
.B2(n_77),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_134),
.B1(n_89),
.B2(n_82),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_78),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_66),
.C(n_36),
.Y(n_163)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_34),
.A3(n_25),
.B1(n_36),
.B2(n_24),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_73),
.B(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_25),
.B1(n_22),
.B2(n_34),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_160),
.B1(n_92),
.B2(n_85),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_139),
.B(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_144),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_80),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_157),
.B(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_151),
.B1(n_158),
.B2(n_127),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_78),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_84),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_164),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_162),
.B1(n_167),
.B2(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_161),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_105),
.B(n_70),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_88),
.B1(n_96),
.B2(n_100),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_68),
.B(n_100),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_75),
.B1(n_76),
.B2(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_107),
.C(n_114),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_83),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_83),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_66),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_1),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_120),
.B(n_107),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_174),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_188),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_116),
.B1(n_137),
.B2(n_109),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_189),
.B1(n_191),
.B2(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_182),
.C(n_187),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_126),
.C(n_130),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_126),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_120),
.B(n_114),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_109),
.B1(n_113),
.B2(n_119),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_113),
.C(n_119),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_194),
.C(n_196),
.Y(n_225)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_149),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_91),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_36),
.B(n_95),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_197),
.B(n_1),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_95),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_1),
.B(n_2),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_209),
.C(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_204),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_140),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_142),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_206),
.B(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_152),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_162),
.B(n_168),
.C(n_166),
.D(n_138),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_214),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_146),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_168),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_168),
.Y(n_214)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx11_ASAP7_75t_R g216 ( 
.A(n_193),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_226),
.C(n_14),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_224),
.B1(n_197),
.B2(n_173),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_155),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_223),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_161),
.C(n_147),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_175),
.Y(n_232)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_10),
.B(n_9),
.C(n_16),
.D(n_15),
.Y(n_223)
);

AOI31xp33_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_85),
.A3(n_10),
.B(n_15),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_186),
.B1(n_179),
.B2(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_188),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_242),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_243),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_181),
.C(n_190),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_236),
.C(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_212),
.C(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_174),
.B1(n_192),
.B2(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_173),
.B1(n_195),
.B2(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_222),
.B1(n_201),
.B2(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_2),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_172),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_178),
.C(n_129),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_129),
.C(n_3),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_254),
.Y(n_274)
);

OA21x2_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_205),
.B(n_208),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_257),
.B(n_228),
.Y(n_272)
);

OAI22x1_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_211),
.B1(n_224),
.B2(n_223),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_250),
.A2(n_230),
.B(n_246),
.Y(n_266)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_247),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_201),
.B1(n_219),
.B2(n_214),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_213),
.B1(n_207),
.B2(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_265),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_247),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_14),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_10),
.C2(n_7),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_2),
.B(n_3),
.Y(n_260)
);

FAx1_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_250),
.CI(n_257),
.CON(n_270),
.SN(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_228),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_286)
);

XOR2x2_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_232),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_278),
.B(n_279),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_234),
.C(n_245),
.Y(n_269)
);

AOI31xp67_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_260),
.A3(n_265),
.B(n_251),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_273),
.Y(n_285)
);

AOI321xp33_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_260),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_8),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_236),
.C(n_231),
.Y(n_273)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_242),
.C(n_4),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_3),
.C(n_4),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_258),
.B1(n_253),
.B2(n_248),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_270),
.B1(n_278),
.B2(n_279),
.Y(n_292)
);

OAI221xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_255),
.B1(n_269),
.B2(n_254),
.C(n_270),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_258),
.B(n_253),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_288),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_289),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_293),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_271),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_285),
.C(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_292),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_289),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_290),
.B1(n_291),
.B2(n_11),
.C(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_303),
.C(n_7),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_304),
.B(n_303),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_302),
.B(n_308),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_298),
.Y(n_311)
);


endmodule