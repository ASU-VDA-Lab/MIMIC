module fake_jpeg_18131_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_17),
.Y(n_82)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_19),
.B1(n_30),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_35),
.B1(n_40),
.B2(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_37),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_47),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_35),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_38),
.B(n_16),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_34),
.B(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_42),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_38),
.B(n_29),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_56),
.B(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_55),
.B1(n_53),
.B2(n_48),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_66),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_55),
.B1(n_53),
.B2(n_19),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_19),
.B1(n_39),
.B2(n_29),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_96),
.B(n_106),
.Y(n_138)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_95),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_34),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_42),
.B1(n_35),
.B2(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_27),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_65),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AND2x4_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_34),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_32),
.Y(n_135)
);

AOI22x1_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_38),
.B1(n_36),
.B2(n_32),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_69),
.B1(n_83),
.B2(n_61),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_38),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_79),
.B1(n_72),
.B2(n_80),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_68),
.B(n_78),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_135),
.B(n_139),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_66),
.B1(n_78),
.B2(n_65),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_77),
.C(n_39),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_96),
.C(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_92),
.B1(n_108),
.B2(n_88),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_85),
.B1(n_107),
.B2(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_38),
.C(n_62),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_86),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_16),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_18),
.B1(n_26),
.B2(n_20),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_141),
.B1(n_85),
.B2(n_15),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_18),
.B1(n_26),
.B2(n_15),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_155),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_138),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_159),
.B1(n_125),
.B2(n_128),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_135),
.B(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_166),
.B(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_129),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_91),
.B1(n_87),
.B2(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_99),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_167),
.B1(n_169),
.B2(n_139),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_96),
.B(n_97),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_106),
.B1(n_98),
.B2(n_100),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_86),
.B1(n_101),
.B2(n_105),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_173),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_103),
.B1(n_104),
.B2(n_87),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_141),
.B1(n_116),
.B2(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_91),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_205),
.B(n_143),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_181),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_183),
.B1(n_194),
.B2(n_196),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_182),
.B1(n_191),
.B2(n_204),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_163),
.B1(n_164),
.B2(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_121),
.B1(n_122),
.B2(n_134),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_145),
.B1(n_161),
.B2(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_91),
.B1(n_73),
.B2(n_38),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_28),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_62),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_166),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_145),
.A2(n_31),
.A3(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_171),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_157),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_202),
.B1(n_160),
.B2(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_28),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_149),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_153),
.C(n_147),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_228),
.C(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_216),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_214),
.B1(n_192),
.B2(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_188),
.B1(n_198),
.B2(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_143),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_195),
.B1(n_188),
.B2(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_219),
.B1(n_226),
.B2(n_201),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_22),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_223),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_24),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_9),
.C(n_12),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_179),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_220),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_232),
.C(n_244),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_196),
.C(n_179),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_200),
.B(n_189),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_225),
.B(n_7),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_203),
.B1(n_206),
.B2(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_206),
.B1(n_224),
.B2(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_203),
.B1(n_176),
.B2(n_199),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_209),
.B1(n_226),
.B2(n_212),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

FAx1_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_223),
.CI(n_215),
.CON(n_249),
.SN(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_237),
.B1(n_238),
.B2(n_246),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_220),
.C(n_176),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_264),
.C(n_233),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_260),
.B(n_10),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_7),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_10),
.C(n_11),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_252),
.Y(n_287)
);

XOR2x2_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_241),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_249),
.B(n_11),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_229),
.C(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_269),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_243),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_234),
.C(n_237),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_243),
.C(n_238),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_10),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_256),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_277),
.A2(n_262),
.B1(n_257),
.B2(n_252),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_11),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_278),
.B(n_251),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_289),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_249),
.B1(n_263),
.B2(n_5),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_2),
.B(n_4),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_265),
.C(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_267),
.C(n_273),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_274),
.B(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_295),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_266),
.C(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_298),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_297),
.A2(n_288),
.B(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_301),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_13),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_296),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_290),
.B(n_294),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_305),
.B(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_303),
.C(n_13),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_4),
.B1(n_6),
.B2(n_308),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_4),
.B(n_6),
.Y(n_313)
);


endmodule