module fake_ariane_528_n_1677 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1677);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1677;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_36),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_24),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_30),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_95),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_27),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_94),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_107),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_31),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_21),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_40),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_49),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_52),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_40),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_26),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_13),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_73),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_1),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_47),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_9),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_11),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_0),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_28),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_70),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_106),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_8),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_114),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_88),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_53),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_46),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_86),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_120),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_58),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_67),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_118),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_138),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_75),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_81),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_17),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_12),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_21),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_59),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_125),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_48),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_84),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_99),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_111),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_65),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_92),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_103),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_79),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_143),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_82),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_83),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_128),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_105),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_135),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_98),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_7),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_76),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_31),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_121),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_43),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_100),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_131),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_93),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_32),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_22),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_60),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_20),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_61),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_35),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_101),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_87),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_150),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_26),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_174),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_174),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_174),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_153),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_166),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_166),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_186),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_156),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_189),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_187),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_223),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_223),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_194),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_188),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_153),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_187),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_213),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_178),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_183),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_191),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_208),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_203),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_233),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_162),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_167),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_157),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_262),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_207),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_214),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_167),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_226),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_232),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_272),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_158),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_239),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_161),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_170),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_168),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_158),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_169),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_157),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_190),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_221),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_192),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_195),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_240),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_294),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_228),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_367),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_311),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_320),
.B(n_257),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_R g384 ( 
.A(n_376),
.B(n_152),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_310),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_277),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_318),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_279),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_197),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_307),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_307),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_321),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_331),
.A2(n_202),
.B(n_201),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_294),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_219),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

OA22x2_ASAP7_75t_L g410 ( 
.A1(n_334),
.A2(n_273),
.B1(n_185),
.B2(n_253),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_327),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_219),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_302),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_316),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_204),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_302),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_332),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_312),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_219),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_312),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_302),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_313),
.A2(n_234),
.B(n_231),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_313),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_374),
.B(n_185),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_342),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_336),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_315),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_324),
.B(n_273),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_325),
.B(n_163),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_317),
.A2(n_229),
.B(n_227),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_317),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_363),
.B(n_163),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g438 ( 
.A(n_319),
.B(n_175),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_338),
.B(n_164),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_352),
.B(n_211),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_322),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_429),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_397),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_328),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_441),
.B(n_350),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_170),
.B1(n_172),
.B2(n_298),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_401),
.B(n_351),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_308),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_381),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_386),
.B(n_221),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_353),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_413),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_413),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_360),
.C(n_355),
.Y(n_463)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_375),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_416),
.A2(n_293),
.B1(n_303),
.B2(n_184),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_403),
.B(n_372),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_385),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_385),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_293),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_416),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_403),
.B(n_314),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_416),
.A2(n_303),
.B1(n_184),
.B2(n_180),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_403),
.B(n_164),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_381),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_338),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_433),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_418),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_433),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_339),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_420),
.B(n_335),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_386),
.B(n_165),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_433),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_394),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_339),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_378),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_422),
.A2(n_265),
.B1(n_264),
.B2(n_261),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_437),
.B(n_340),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_378),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_437),
.B(n_340),
.Y(n_508)
);

CKINVDCx6p67_ASAP7_75t_R g509 ( 
.A(n_418),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_388),
.B(n_171),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_409),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_409),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_439),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_418),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_341),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_380),
.B(n_341),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_379),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_410),
.A2(n_356),
.B1(n_362),
.B2(n_361),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_343),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_388),
.B(n_171),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_377),
.B(n_343),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_432),
.B(n_344),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_380),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_400),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_399),
.B(n_173),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_377),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_411),
.B(n_173),
.Y(n_534)
);

INVxp67_ASAP7_75t_R g535 ( 
.A(n_407),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_379),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_411),
.B(n_249),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_400),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_400),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_380),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_380),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_379),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_390),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_406),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_417),
.B(n_249),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_379),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_344),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_439),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_439),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_382),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_390),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_390),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_382),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_382),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_382),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_389),
.A2(n_172),
.B1(n_298),
.B2(n_368),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_440),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_391),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_395),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_430),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_395),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_395),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_377),
.A2(n_330),
.B1(n_358),
.B2(n_364),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_427),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_427),
.B(n_250),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_396),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_377),
.B(n_348),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_396),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_391),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_SL g579 ( 
.A1(n_439),
.A2(n_362),
.B(n_361),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_430),
.A2(n_280),
.B1(n_243),
.B2(n_245),
.Y(n_580)
);

CKINVDCx6p67_ASAP7_75t_R g581 ( 
.A(n_414),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_377),
.A2(n_269),
.B1(n_281),
.B2(n_241),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_400),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_377),
.B(n_349),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_400),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_392),
.B(n_349),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_410),
.A2(n_359),
.B1(n_357),
.B2(n_356),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_419),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_443),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_503),
.A2(n_387),
.B1(n_383),
.B2(n_252),
.C(n_256),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_392),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_500),
.B(n_392),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_508),
.B(n_392),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_480),
.B(n_392),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_524),
.A2(n_426),
.B1(n_392),
.B2(n_412),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_512),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_454),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_494),
.B(n_387),
.C(n_383),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_480),
.B(n_384),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_542),
.B(n_426),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_516),
.B(n_426),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_486),
.A2(n_496),
.B1(n_457),
.B2(n_473),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_542),
.B(n_426),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_482),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_512),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_426),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_562),
.B(n_426),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_472),
.B(n_406),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_465),
.B(n_406),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_457),
.B(n_406),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_461),
.B(n_473),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_484),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_515),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_524),
.A2(n_406),
.B1(n_412),
.B2(n_440),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_449),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_461),
.B(n_406),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_501),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_460),
.B(n_414),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_464),
.B(n_486),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_513),
.B(n_412),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_562),
.B(n_412),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_482),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_446),
.B(n_428),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_509),
.B(n_354),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_464),
.B(n_496),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_552),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_455),
.B(n_384),
.Y(n_634)
);

BUFx5_ASAP7_75t_L g635 ( 
.A(n_529),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_449),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_474),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_445),
.B(n_428),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_467),
.B(n_412),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_474),
.B(n_440),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_464),
.B(n_250),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_551),
.A2(n_410),
.B1(n_405),
.B2(n_402),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_552),
.B(n_436),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_450),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_509),
.B(n_230),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_524),
.A2(n_410),
.B1(n_423),
.B2(n_402),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_464),
.B(n_251),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_526),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_586),
.B(n_436),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_448),
.B(n_393),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_535),
.B(n_440),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_524),
.A2(n_410),
.B1(n_405),
.B2(n_423),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_517),
.A2(n_408),
.B(n_402),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_562),
.B(n_436),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_564),
.B(n_400),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_564),
.B(n_405),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_408),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_533),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_581),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_525),
.B(n_251),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_468),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_581),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_495),
.B(n_301),
.C(n_247),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_546),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_525),
.B(n_408),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_547),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_502),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_547),
.B(n_423),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_505),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_505),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_531),
.A2(n_393),
.B1(n_415),
.B2(n_260),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_507),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_545),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_554),
.B(n_424),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_573),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_531),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_527),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_555),
.B(n_424),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_463),
.B(n_415),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_535),
.B(n_354),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_565),
.B(n_424),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_568),
.B(n_424),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_578),
.B(n_424),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_582),
.B(n_267),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_569),
.B(n_295),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_479),
.B(n_424),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_531),
.A2(n_424),
.B1(n_434),
.B2(n_435),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_518),
.Y(n_690)
);

BUFx5_ASAP7_75t_L g691 ( 
.A(n_529),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_510),
.B(n_299),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_490),
.B(n_579),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_522),
.B(n_357),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_573),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_573),
.B(n_154),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_530),
.B(n_359),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_507),
.Y(n_698)
);

BUFx5_ASAP7_75t_L g699 ( 
.A(n_538),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_504),
.B(n_159),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_576),
.A2(n_322),
.B1(n_255),
.B2(n_274),
.Y(n_702)
);

AO221x1_ASAP7_75t_L g703 ( 
.A1(n_559),
.A2(n_179),
.B1(n_175),
.B2(n_209),
.C(n_296),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_516),
.B(n_160),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_453),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_518),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_476),
.A2(n_217),
.B1(n_300),
.B2(n_290),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_519),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_528),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_536),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_536),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_534),
.B(n_268),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_475),
.A2(n_434),
.B1(n_435),
.B2(n_396),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_444),
.B(n_434),
.Y(n_715)
);

AO221x1_ASAP7_75t_L g716 ( 
.A1(n_580),
.A2(n_175),
.B1(n_179),
.B2(n_209),
.C(n_224),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_543),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_545),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_447),
.B(n_396),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_444),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_495),
.B(n_287),
.C(n_435),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_584),
.B(n_176),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_521),
.B(n_177),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_544),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_452),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_550),
.A2(n_434),
.B1(n_435),
.B2(n_398),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_470),
.B(n_434),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_471),
.B(n_434),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_453),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_456),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_398),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_548),
.B(n_181),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_574),
.B(n_182),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_498),
.B(n_434),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_456),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_563),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_563),
.B(n_193),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_538),
.A2(n_425),
.B1(n_421),
.B2(n_404),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_539),
.A2(n_425),
.B1(n_421),
.B2(n_404),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_458),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_458),
.B(n_398),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_572),
.B(n_198),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_520),
.B(n_199),
.Y(n_743)
);

BUFx8_ASAP7_75t_L g744 ( 
.A(n_539),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_469),
.B(n_398),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_540),
.B(n_404),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_523),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_451),
.B(n_404),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_593),
.B(n_587),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_639),
.A2(n_540),
.B1(n_585),
.B2(n_583),
.Y(n_750)
);

CKINVDCx8_ASAP7_75t_R g751 ( 
.A(n_606),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_611),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_636),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_675),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_593),
.A2(n_583),
.B1(n_585),
.B2(n_553),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_620),
.B(n_469),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_549),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_592),
.B(n_466),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_682),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_611),
.B(n_668),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_644),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_592),
.A2(n_553),
.B1(n_577),
.B2(n_575),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_596),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_638),
.B(n_483),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_589),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_663),
.B(n_487),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_597),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_629),
.Y(n_768)
);

NOR2x2_ASAP7_75t_L g769 ( 
.A(n_623),
.B(n_483),
.Y(n_769)
);

AO22x1_ASAP7_75t_L g770 ( 
.A1(n_742),
.A2(n_514),
.B1(n_288),
.B2(n_286),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_631),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_605),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_637),
.B(n_549),
.Y(n_773)
);

OAI21xp33_ASAP7_75t_L g774 ( 
.A1(n_687),
.A2(n_506),
.B(n_488),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_659),
.B(n_556),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_635),
.B(n_523),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_603),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_612),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_591),
.B(n_489),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_640),
.B(n_651),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_675),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_598),
.B(n_511),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_607),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_613),
.B(n_459),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_617),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_556),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_590),
.B(n_459),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_622),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_649),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_625),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_666),
.B(n_557),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_595),
.B(n_588),
.Y(n_793)
);

BUFx4f_ASAP7_75t_L g794 ( 
.A(n_660),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_619),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_666),
.B(n_557),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_695),
.B(n_462),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_619),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_SL g799 ( 
.A1(n_630),
.A2(n_222),
.B1(n_236),
.B2(n_235),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_645),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_594),
.B(n_462),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_677),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_633),
.B(n_558),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_661),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_558),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_595),
.B(n_523),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_601),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_601),
.B(n_523),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_693),
.A2(n_561),
.B(n_577),
.C(n_575),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_729),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_669),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_667),
.B(n_561),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_736),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_671),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_705),
.B(n_462),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_679),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_693),
.A2(n_571),
.B(n_570),
.C(n_567),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_746),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_690),
.B(n_567),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_709),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_713),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_692),
.B(n_212),
.C(n_206),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_717),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_643),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_706),
.B(n_570),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_744),
.A2(n_571),
.B1(n_485),
.B2(n_491),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_635),
.B(n_523),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_610),
.A2(n_716),
.B1(n_703),
.B2(n_688),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_678),
.B(n_481),
.Y(n_831)
);

CKINVDCx6p67_ASAP7_75t_R g832 ( 
.A(n_729),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_656),
.A2(n_481),
.B(n_497),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_634),
.B(n_497),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_602),
.B(n_499),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_664),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_704),
.B(n_646),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_616),
.B(n_532),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_736),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_697),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_720),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_672),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_725),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_730),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_681),
.B(n_499),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_674),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_688),
.A2(n_491),
.B1(n_493),
.B2(n_492),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_714),
.A2(n_492),
.B1(n_493),
.B2(n_485),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_615),
.B(n_532),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_599),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_746),
.B(n_514),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_735),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_621),
.B(n_532),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_656),
.A2(n_588),
.B(n_560),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_731),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_626),
.B(n_532),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_655),
.Y(n_857)
);

OR2x2_ASAP7_75t_SL g858 ( 
.A(n_665),
.B(n_421),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_662),
.B(n_712),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_698),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_736),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_746),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_702),
.A2(n_743),
.B1(n_731),
.B2(n_642),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_628),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_650),
.A2(n_421),
.B(n_425),
.C(n_5),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_657),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_732),
.A2(n_588),
.B1(n_560),
.B2(n_259),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_676),
.A2(n_685),
.B(n_684),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_635),
.B(n_560),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_696),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_700),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_715),
.A2(n_425),
.B(n_438),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_628),
.B(n_560),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_657),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_600),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_658),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_686),
.B(n_618),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_702),
.A2(n_438),
.B1(n_419),
.B2(n_514),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_707),
.B(n_0),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_708),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_658),
.Y(n_882)
);

BUFx10_ASAP7_75t_L g883 ( 
.A(n_740),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_710),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_670),
.B(n_588),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_711),
.Y(n_886)
);

AO22x1_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_514),
.B1(n_254),
.B2(n_244),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_718),
.B(n_514),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_724),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_747),
.B(n_419),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_747),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_733),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_741),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_741),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_635),
.B(n_283),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_745),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_745),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_701),
.B(n_4),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_748),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_635),
.B(n_419),
.Y(n_900)
);

AO22x2_ASAP7_75t_L g901 ( 
.A1(n_727),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_600),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_719),
.B(n_210),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_673),
.B(n_419),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_604),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_604),
.B(n_608),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_723),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_608),
.B(n_215),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_641),
.B(n_289),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_737),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_722),
.B(n_6),
.Y(n_911)
);

BUFx5_ASAP7_75t_L g912 ( 
.A(n_691),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_648),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_R g914 ( 
.A(n_728),
.B(n_216),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_609),
.B(n_218),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_691),
.B(n_419),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_691),
.A2(n_438),
.B1(n_296),
.B2(n_179),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_647),
.B(n_9),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_840),
.B(n_609),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_868),
.A2(n_632),
.B(n_624),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_780),
.B(n_699),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_SL g922 ( 
.A1(n_795),
.A2(n_685),
.B(n_676),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_795),
.B(n_699),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_822),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_859),
.A2(n_654),
.B(n_726),
.C(n_684),
.Y(n_925)
);

OAI22x1_ASAP7_75t_L g926 ( 
.A1(n_859),
.A2(n_653),
.B1(n_680),
.B2(n_683),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_798),
.B(n_699),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_753),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_798),
.A2(n_680),
.B1(n_683),
.B2(n_715),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_898),
.A2(n_734),
.B(n_738),
.C(n_739),
.Y(n_930)
);

NOR2x1_ASAP7_75t_R g931 ( 
.A(n_768),
.B(n_810),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_866),
.B(n_699),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_689),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_862),
.B(n_296),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_864),
.B(n_10),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_823),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_918),
.A2(n_258),
.B1(n_220),
.B2(n_278),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_SL g938 ( 
.A1(n_776),
.A2(n_10),
.B(n_20),
.C(n_23),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_837),
.B(n_276),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_761),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_829),
.A2(n_242),
.B(n_225),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_751),
.B(n_237),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_789),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_829),
.A2(n_270),
.B(n_263),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_862),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_854),
.A2(n_438),
.B(n_119),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_800),
.B(n_23),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_805),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_869),
.A2(n_271),
.B(n_296),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_825),
.Y(n_950)
);

AND3x4_ASAP7_75t_L g951 ( 
.A(n_802),
.B(n_870),
.C(n_794),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_SL g952 ( 
.A(n_892),
.B(n_25),
.C(n_28),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_875),
.A2(n_179),
.B1(n_209),
.B2(n_224),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_765),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_837),
.B(n_794),
.Y(n_955)
);

OR2x4_ASAP7_75t_L g956 ( 
.A(n_898),
.B(n_25),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_808),
.B(n_438),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_862),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_862),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_911),
.A2(n_29),
.B(n_32),
.C(n_34),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_836),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_864),
.B(n_29),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_851),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_764),
.B(n_34),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_850),
.B(n_35),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_851),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_799),
.B(n_905),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_913),
.B(n_39),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_900),
.A2(n_224),
.B(n_275),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_812),
.B(n_132),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_775),
.B(n_39),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_769),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_911),
.A2(n_41),
.B(n_42),
.C(n_438),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_785),
.A2(n_438),
.B(n_275),
.C(n_224),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_877),
.B(n_438),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_757),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_916),
.A2(n_44),
.B(n_51),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_882),
.B(n_905),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_820),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_916),
.A2(n_55),
.B(n_68),
.Y(n_982)
);

BUFx12f_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_766),
.B(n_78),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_832),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_797),
.B(n_438),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_888),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_754),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_767),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_758),
.A2(n_779),
.B1(n_749),
.B2(n_906),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_766),
.B(n_89),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_797),
.B(n_438),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_438),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_876),
.B(n_116),
.Y(n_994)
);

AOI22x1_ASAP7_75t_L g995 ( 
.A1(n_857),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_813),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_756),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_816),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_855),
.B(n_147),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_880),
.B(n_772),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_SL g1001 ( 
.A(n_820),
.B(n_148),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_757),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_788),
.A2(n_779),
.B(n_878),
.C(n_785),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_902),
.B(n_893),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_902),
.B(n_894),
.Y(n_1005)
);

INVx3_ASAP7_75t_SL g1006 ( 
.A(n_910),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_833),
.A2(n_819),
.B(n_811),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_896),
.B(n_897),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_888),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_874),
.A2(n_849),
.B(n_853),
.Y(n_1010)
);

CKINVDCx11_ASAP7_75t_R g1011 ( 
.A(n_883),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_754),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_806),
.A2(n_814),
.B(n_856),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_835),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_842),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_788),
.A2(n_878),
.B(n_774),
.C(n_824),
.Y(n_1016)
);

CKINVDCx6p67_ASAP7_75t_R g1017 ( 
.A(n_757),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_778),
.A2(n_818),
.B1(n_790),
.B2(n_786),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_871),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_883),
.B(n_773),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_899),
.B(n_826),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_847),
.A2(n_755),
.B(n_787),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_824),
.A2(n_835),
.B1(n_914),
.B2(n_809),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_781),
.Y(n_1024)
);

NAND2x2_ASAP7_75t_L g1025 ( 
.A(n_907),
.B(n_817),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_752),
.B(n_783),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_838),
.A2(n_895),
.B(n_807),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_750),
.B(n_863),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_863),
.A2(n_750),
.B1(n_884),
.B2(n_889),
.Y(n_1029)
);

AND2x2_ASAP7_75t_SL g1030 ( 
.A(n_828),
.B(n_830),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_SL g1031 ( 
.A(n_865),
.B(n_828),
.C(n_909),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_792),
.B(n_796),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_803),
.A2(n_793),
.B(n_845),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_870),
.B(n_831),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_914),
.A2(n_801),
.B1(n_831),
.B2(n_760),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_821),
.B(n_827),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_841),
.B(n_843),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_815),
.B(n_763),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_846),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_SL g1040 ( 
.A(n_834),
.B(n_908),
.C(n_915),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_754),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_865),
.A2(n_801),
.B(n_903),
.C(n_784),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_860),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_901),
.B(n_844),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_777),
.A2(n_852),
.B(n_885),
.C(n_891),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_872),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_885),
.A2(n_830),
.B(n_867),
.C(n_762),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_891),
.A2(n_848),
.B(n_873),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_963),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_984),
.A2(n_770),
.B(n_887),
.C(n_904),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1000),
.B(n_901),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_997),
.B(n_886),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_919),
.B(n_881),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_945),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_1007),
.A2(n_890),
.B(n_917),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_990),
.A2(n_912),
.B(n_901),
.Y(n_1057)
);

AOI221x1_ASAP7_75t_L g1058 ( 
.A1(n_1016),
.A2(n_754),
.B1(n_782),
.B2(n_839),
.C(n_861),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_963),
.B(n_782),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_917),
.B(n_879),
.Y(n_1060)
);

OA22x2_ASAP7_75t_L g1061 ( 
.A1(n_951),
.A2(n_858),
.B1(n_879),
.B2(n_782),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_936),
.Y(n_1062)
);

AOI211x1_ASAP7_75t_L g1063 ( 
.A1(n_1018),
.A2(n_782),
.B(n_839),
.C(n_861),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_922),
.A2(n_912),
.B(n_839),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_991),
.A2(n_839),
.B(n_861),
.C(n_912),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_990),
.A2(n_912),
.B(n_861),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_1034),
.B(n_912),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_920),
.A2(n_912),
.B(n_1027),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_932),
.A2(n_927),
.B(n_923),
.Y(n_1069)
);

OAI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_1040),
.A2(n_962),
.B(n_935),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_967),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1048),
.A2(n_925),
.B(n_929),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_960),
.B(n_975),
.C(n_1047),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_929),
.A2(n_926),
.A3(n_953),
.B(n_1010),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_950),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_980),
.B(n_1021),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_937),
.A2(n_1008),
.B1(n_1028),
.B2(n_932),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_930),
.A2(n_1042),
.B(n_1023),
.C(n_1026),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_921),
.A2(n_1013),
.B(n_1032),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_954),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_968),
.A2(n_1031),
.B(n_966),
.C(n_969),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_SL g1083 ( 
.A1(n_1036),
.A2(n_953),
.B(n_994),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_940),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_1022),
.A2(n_970),
.B(n_1044),
.Y(n_1085)
);

OAI22x1_ASAP7_75t_L g1086 ( 
.A1(n_974),
.A2(n_1035),
.B1(n_956),
.B2(n_981),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_989),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1045),
.A2(n_982),
.B(n_979),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_977),
.A2(n_965),
.B(n_993),
.Y(n_1089)
);

NAND3x1_ASAP7_75t_L g1090 ( 
.A(n_956),
.B(n_1020),
.C(n_972),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_995),
.A2(n_934),
.B(n_949),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_934),
.A2(n_1018),
.B(n_1012),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1001),
.A2(n_1037),
.B(n_976),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_928),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1030),
.A2(n_1025),
.B1(n_1014),
.B2(n_1034),
.Y(n_1095)
);

AOI31xp67_ASAP7_75t_L g1096 ( 
.A1(n_986),
.A2(n_992),
.A3(n_1039),
.B(n_998),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_974),
.B(n_981),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_967),
.B(n_1034),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_941),
.A2(n_944),
.B(n_933),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1038),
.A2(n_952),
.B(n_1009),
.C(n_987),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1046),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1041),
.B(n_987),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_961),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_943),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_948),
.B(n_955),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1019),
.B(n_1009),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_985),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_947),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_945),
.Y(n_1110)
);

AOI31xp67_ASAP7_75t_L g1111 ( 
.A1(n_964),
.A2(n_1043),
.A3(n_1015),
.B(n_996),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_978),
.A2(n_1002),
.B(n_1029),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1006),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_938),
.A2(n_1012),
.B(n_988),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_999),
.A2(n_939),
.B(n_973),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_942),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_957),
.A2(n_1024),
.B(n_978),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_983),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1002),
.A2(n_1017),
.B(n_988),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_957),
.A2(n_958),
.B(n_959),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

NAND3x1_ASAP7_75t_L g1122 ( 
.A(n_931),
.B(n_971),
.C(n_945),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_945),
.B(n_958),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_959),
.A2(n_990),
.B(n_920),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1003),
.A2(n_922),
.B(n_990),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_919),
.B(n_620),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1007),
.A2(n_920),
.B(n_946),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_929),
.A2(n_926),
.A3(n_1016),
.B(n_990),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_SL g1130 ( 
.A(n_961),
.B(n_751),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_943),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_920),
.B(n_946),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_990),
.A2(n_1003),
.B(n_991),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_1012),
.B(n_980),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_928),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_943),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_1011),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_1011),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1000),
.B(n_636),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_924),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_L g1142 ( 
.A(n_1003),
.B(n_795),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_924),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_920),
.A2(n_1027),
.B(n_1033),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_859),
.B1(n_795),
.B2(n_798),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1007),
.A2(n_920),
.B(n_946),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_963),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1003),
.A2(n_922),
.B(n_990),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_990),
.B(n_984),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_963),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_919),
.B(n_620),
.Y(n_1155)
);

O2A1O1Ixp5_ASAP7_75t_L g1156 ( 
.A1(n_984),
.A2(n_991),
.B(n_1003),
.C(n_1016),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_968),
.B(n_372),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_924),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_963),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1030),
.A2(n_859),
.B1(n_795),
.B2(n_798),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1007),
.A2(n_920),
.B(n_946),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_943),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1003),
.A2(n_798),
.B1(n_795),
.B2(n_840),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1007),
.A2(n_1003),
.B(n_1016),
.Y(n_1164)
);

AOI21x1_ASAP7_75t_L g1165 ( 
.A1(n_920),
.A2(n_1027),
.B(n_1033),
.Y(n_1165)
);

O2A1O1Ixp5_ASAP7_75t_L g1166 ( 
.A1(n_984),
.A2(n_991),
.B(n_1003),
.C(n_1016),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_968),
.B(n_372),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_924),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_940),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_919),
.B(n_620),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_SL g1172 ( 
.A1(n_960),
.A2(n_1003),
.B1(n_975),
.B2(n_990),
.C(n_898),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_984),
.A2(n_991),
.B(n_990),
.Y(n_1173)
);

AND2x6_ASAP7_75t_L g1174 ( 
.A(n_958),
.B(n_862),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1000),
.B(n_636),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_943),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1003),
.A2(n_446),
.B(n_465),
.C(n_859),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_990),
.A2(n_920),
.B(n_1003),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_963),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1161),
.A2(n_1165),
.B(n_1144),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1152),
.A2(n_1082),
.B1(n_1133),
.B2(n_1156),
.C(n_1166),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1173),
.A2(n_1160),
.B1(n_1146),
.B2(n_1060),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1177),
.A2(n_1163),
.B(n_1149),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1068),
.A2(n_1124),
.B(n_1093),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1054),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1054),
.B(n_1110),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1091),
.A2(n_1066),
.B(n_1088),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1062),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1136),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1174),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1129),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1174),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1072),
.A2(n_1125),
.B(n_1149),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1146),
.A2(n_1160),
.B1(n_1060),
.B2(n_1061),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1094),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1075),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1076),
.B(n_1126),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1064),
.A2(n_1178),
.B(n_1134),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1083),
.A2(n_1073),
.B(n_1155),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1140),
.B(n_1175),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1138),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1073),
.A2(n_1157),
.B1(n_1167),
.B2(n_1051),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1128),
.A2(n_1145),
.B(n_1168),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1058),
.A2(n_1153),
.B(n_1151),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1171),
.B(n_1070),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1070),
.A2(n_1170),
.B1(n_1150),
.B2(n_1101),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1142),
.A2(n_1078),
.B(n_1077),
.C(n_1084),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1164),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1170),
.A2(n_1090),
.B1(n_1109),
.B2(n_1053),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_1116),
.B(n_1104),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1055),
.A2(n_1092),
.B(n_1100),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1067),
.B(n_1098),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1172),
.A2(n_1050),
.B(n_1081),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1099),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1114),
.A2(n_1112),
.B(n_1095),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1089),
.A2(n_1102),
.B(n_1143),
.Y(n_1217)
);

CKINVDCx11_ASAP7_75t_R g1218 ( 
.A(n_1139),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1080),
.A2(n_1158),
.B(n_1141),
.Y(n_1219)
);

NOR4xp25_ASAP7_75t_L g1220 ( 
.A(n_1122),
.B(n_1106),
.C(n_1087),
.D(n_1169),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1115),
.A2(n_1085),
.B(n_1119),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1135),
.A2(n_1096),
.B(n_1103),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1129),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1097),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1110),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1067),
.B(n_1098),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1059),
.B(n_1049),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1129),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1074),
.Y(n_1229)
);

AO32x2_ASAP7_75t_L g1230 ( 
.A1(n_1063),
.A2(n_1074),
.A3(n_1086),
.B1(n_1108),
.B2(n_1052),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1105),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1117),
.A2(n_1123),
.B(n_1121),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1067),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1131),
.A2(n_1137),
.A3(n_1162),
.B(n_1176),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1049),
.A2(n_1179),
.B(n_1071),
.Y(n_1235)
);

BUFx8_ASAP7_75t_L g1236 ( 
.A(n_1113),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1107),
.A2(n_1071),
.B1(n_1159),
.B2(n_1154),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1148),
.A2(n_1179),
.B(n_1154),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1148),
.A2(n_1120),
.B(n_1059),
.C(n_1130),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1118),
.A2(n_1174),
.B1(n_639),
.B2(n_1152),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1118),
.A2(n_1057),
.B(n_1058),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1111),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1057),
.A2(n_1058),
.B(n_1128),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1111),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1056),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1056),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1056),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1067),
.B(n_1098),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1067),
.B(n_1098),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1140),
.B(n_1175),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1057),
.A2(n_1058),
.B(n_1128),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1111),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1111),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1152),
.B(n_1133),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1136),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1111),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1111),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1067),
.B(n_1061),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1067),
.B(n_1061),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1152),
.A2(n_639),
.B1(n_1028),
.B2(n_1173),
.Y(n_1260)
);

CKINVDCx11_ASAP7_75t_R g1261 ( 
.A(n_1138),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1056),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1056),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1140),
.B(n_1175),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1067),
.B(n_1098),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1152),
.A2(n_1133),
.B1(n_1160),
.B2(n_1146),
.Y(n_1268)
);

AO21x1_ASAP7_75t_L g1269 ( 
.A1(n_1152),
.A2(n_1082),
.B(n_1125),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1054),
.B(n_945),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1067),
.B(n_1061),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1152),
.A2(n_639),
.B1(n_1028),
.B2(n_1173),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1111),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_SL g1275 ( 
.A(n_1104),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1140),
.B(n_1175),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1136),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1111),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1173),
.A2(n_1058),
.A3(n_1057),
.B(n_1079),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1152),
.A2(n_639),
.B1(n_1028),
.B2(n_1173),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1056),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1156),
.A2(n_1166),
.B(n_1152),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1156),
.A2(n_1166),
.B(n_1152),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1056),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1084),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1111),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1140),
.B(n_1175),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1076),
.B(n_1126),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1173),
.B(n_1152),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1132),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1173),
.A2(n_1058),
.A3(n_1057),
.B(n_1079),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1056),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1152),
.A2(n_1166),
.B(n_1156),
.C(n_1177),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_1166),
.B(n_1152),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1116),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1152),
.B(n_1133),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1056),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1111),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1163),
.A2(n_1077),
.A3(n_1095),
.B1(n_990),
.B2(n_929),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1219),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1194),
.A2(n_1289),
.B(n_1254),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1254),
.B(n_1297),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1202),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1198),
.B(n_1288),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1224),
.B(n_1201),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1250),
.B(n_1265),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1213),
.B(n_1226),
.Y(n_1308)
);

AOI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1206),
.A2(n_1203),
.B1(n_1183),
.B2(n_1268),
.C(n_1182),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1297),
.A2(n_1183),
.B1(n_1206),
.B2(n_1195),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1192),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1195),
.A2(n_1184),
.B1(n_1260),
.B2(n_1280),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1218),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1285),
.B(n_1196),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1285),
.B(n_1276),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1287),
.B(n_1190),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1203),
.A2(n_1275),
.B1(n_1215),
.B2(n_1200),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1294),
.A2(n_1208),
.B(n_1207),
.C(n_1283),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1204),
.A2(n_1188),
.B(n_1209),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1282),
.A2(n_1295),
.B(n_1269),
.C(n_1214),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1260),
.A2(n_1273),
.B1(n_1280),
.B2(n_1240),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1189),
.B(n_1197),
.Y(n_1322)
);

O2A1O1Ixp5_ASAP7_75t_L g1323 ( 
.A1(n_1222),
.A2(n_1237),
.B(n_1228),
.C(n_1223),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1273),
.A2(n_1240),
.B1(n_1210),
.B2(n_1255),
.Y(n_1325)
);

O2A1O1Ixp5_ASAP7_75t_L g1326 ( 
.A1(n_1237),
.A2(n_1223),
.B(n_1228),
.C(n_1185),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1247),
.B(n_1262),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1191),
.A2(n_1193),
.B(n_1239),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1236),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1264),
.B(n_1281),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1277),
.A2(n_1259),
.B1(n_1271),
.B2(n_1258),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1236),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1284),
.B(n_1293),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1298),
.B(n_1213),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1191),
.A2(n_1193),
.B(n_1258),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1217),
.B(n_1220),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1181),
.A2(n_1199),
.B(n_1212),
.Y(n_1337)
);

CKINVDCx9p33_ASAP7_75t_R g1338 ( 
.A(n_1300),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1231),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1248),
.B(n_1249),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1216),
.A2(n_1211),
.B(n_1229),
.C(n_1205),
.Y(n_1341)
);

INVx8_ASAP7_75t_L g1342 ( 
.A(n_1296),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_SL g1343 ( 
.A1(n_1266),
.A2(n_1300),
.B(n_1292),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1227),
.A2(n_1251),
.B(n_1243),
.C(n_1225),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1227),
.A2(n_1296),
.B1(n_1275),
.B2(n_1251),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1300),
.A2(n_1292),
.B(n_1279),
.Y(n_1347)
);

AND2x2_ASAP7_75t_SL g1348 ( 
.A(n_1241),
.B(n_1233),
.Y(n_1348)
);

INVx8_ASAP7_75t_L g1349 ( 
.A(n_1186),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1243),
.A2(n_1251),
.B(n_1241),
.C(n_1253),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1202),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1186),
.B(n_1234),
.Y(n_1352)
);

AOI221x1_ASAP7_75t_SL g1353 ( 
.A1(n_1300),
.A2(n_1261),
.B1(n_1218),
.B2(n_1215),
.C(n_1256),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1241),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1233),
.B(n_1279),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1230),
.B(n_1232),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1230),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1187),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1235),
.B(n_1238),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1292),
.B(n_1270),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1242),
.A2(n_1299),
.B(n_1274),
.C(n_1278),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1261),
.B(n_1221),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.B(n_1252),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1180),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1257),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1263),
.A2(n_1267),
.B(n_1272),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1291),
.A2(n_1152),
.B(n_1082),
.C(n_1177),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1208),
.A2(n_1156),
.B(n_1166),
.C(n_1152),
.Y(n_1369)
);

NOR2xp67_ASAP7_75t_L g1370 ( 
.A(n_1254),
.B(n_1297),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1206),
.A2(n_956),
.B1(n_1297),
.B2(n_1254),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1255),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1268),
.A2(n_1152),
.B(n_1082),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1202),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1254),
.B(n_1297),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1301),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1363),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1336),
.A2(n_1302),
.B(n_1350),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1311),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1311),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1330),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1339),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1362),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1359),
.B(n_1364),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1353),
.B(n_1322),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1364),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1312),
.A2(n_1310),
.B1(n_1321),
.B2(n_1371),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1324),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1327),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1367),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1367),
.B(n_1356),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1333),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1354),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1357),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1303),
.B(n_1375),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1397)
);

CKINVDCx16_ASAP7_75t_R g1398 ( 
.A(n_1332),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1319),
.B(n_1337),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1319),
.B(n_1337),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1370),
.B(n_1305),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1361),
.A2(n_1360),
.B(n_1369),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1355),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1366),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1314),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1315),
.B(n_1334),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1338),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1306),
.B(n_1348),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1326),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1323),
.A2(n_1369),
.B(n_1309),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1346),
.B(n_1307),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1348),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1349),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1365),
.B(n_1316),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1323),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1338),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1415),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1392),
.B(n_1341),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1394),
.Y(n_1421)
);

OAI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1388),
.A2(n_1368),
.B(n_1325),
.C(n_1351),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1387),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1391),
.B(n_1343),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1399),
.B(n_1347),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1385),
.B(n_1308),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1378),
.B(n_1403),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1379),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1381),
.B(n_1372),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1340),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1379),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1397),
.B(n_1332),
.Y(n_1432)
);

CKINVDCx8_ASAP7_75t_R g1433 ( 
.A(n_1411),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1378),
.B(n_1328),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1308),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1380),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1405),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1376),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1391),
.B(n_1329),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1377),
.B(n_1331),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1388),
.A2(n_1313),
.B1(n_1342),
.B2(n_1358),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1387),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1405),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1438),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1445)
);

AOI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1422),
.A2(n_1397),
.B(n_1412),
.C(n_1386),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1426),
.B(n_1424),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1428),
.B(n_1406),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1433),
.B(n_1412),
.C(n_1411),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1422),
.B(n_1411),
.C(n_1410),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1438),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1441),
.A2(n_1411),
.B1(n_1413),
.B2(n_1386),
.Y(n_1454)
);

OAI33xp33_ASAP7_75t_L g1455 ( 
.A1(n_1429),
.A2(n_1402),
.A3(n_1389),
.B1(n_1390),
.B2(n_1393),
.B3(n_1407),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1441),
.A2(n_1411),
.B1(n_1413),
.B2(n_1398),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1406),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1435),
.B(n_1384),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1433),
.A2(n_1411),
.B1(n_1417),
.B2(n_1410),
.C(n_1413),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1429),
.B(n_1402),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1438),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_R g1462 ( 
.A(n_1432),
.B(n_1304),
.Y(n_1462)
);

OAI33xp33_ASAP7_75t_L g1463 ( 
.A1(n_1440),
.A2(n_1393),
.A3(n_1407),
.B1(n_1396),
.B2(n_1382),
.B3(n_1395),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1425),
.A2(n_1409),
.B1(n_1395),
.B2(n_1418),
.C(n_1408),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1420),
.A2(n_1417),
.B1(n_1378),
.B2(n_1418),
.Y(n_1465)
);

AOI211xp5_ASAP7_75t_L g1466 ( 
.A1(n_1425),
.A2(n_1424),
.B(n_1432),
.C(n_1420),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1374),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_L g1468 ( 
.A(n_1425),
.B(n_1400),
.C(n_1405),
.D(n_1384),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1442),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1407),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1425),
.A2(n_1417),
.B1(n_1401),
.B2(n_1409),
.C(n_1396),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1420),
.A2(n_1414),
.B1(n_1378),
.B2(n_1404),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_SL g1473 ( 
.A(n_1419),
.B(n_1383),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1431),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1431),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1421),
.B(n_1409),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1427),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1435),
.B(n_1384),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1475),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1474),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1469),
.Y(n_1481)
);

CKINVDCx14_ASAP7_75t_R g1482 ( 
.A(n_1462),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1466),
.B(n_1424),
.Y(n_1483)
);

INVx4_ASAP7_75t_SL g1484 ( 
.A(n_1449),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1466),
.B(n_1435),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1444),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1453),
.B(n_1421),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_SL g1489 ( 
.A(n_1446),
.B(n_1433),
.C(n_1423),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1434),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1446),
.B(n_1427),
.C(n_1434),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1449),
.B(n_1435),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1449),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1452),
.A2(n_1434),
.B(n_1378),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1452),
.A2(n_1433),
.B(n_1439),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1453),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1477),
.A2(n_1443),
.B(n_1437),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1473),
.B(n_1442),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1464),
.A2(n_1443),
.B(n_1437),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1461),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1486),
.B(n_1445),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1485),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1485),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1487),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1487),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1502),
.B(n_1489),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1502),
.B(n_1450),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1445),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1497),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1486),
.B(n_1447),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1483),
.B(n_1454),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1484),
.B(n_1447),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1502),
.B(n_1470),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1497),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1484),
.B(n_1448),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1484),
.B(n_1448),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1482),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1500),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1483),
.B(n_1465),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1484),
.B(n_1478),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1495),
.A2(n_1459),
.B(n_1456),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1503),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1498),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1499),
.B(n_1398),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1491),
.B(n_1475),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1482),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1503),
.Y(n_1536)
);

AND2x2_ASAP7_75t_SL g1537 ( 
.A(n_1491),
.B(n_1419),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1479),
.Y(n_1538)
);

AND2x2_ASAP7_75t_SL g1539 ( 
.A(n_1501),
.B(n_1419),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1540)
);

NAND4xp25_ASAP7_75t_L g1541 ( 
.A(n_1489),
.B(n_1468),
.C(n_1471),
.D(n_1467),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1498),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1480),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1543),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1543),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1506),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1541),
.B(n_1494),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1538),
.B(n_1501),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1535),
.B(n_1522),
.Y(n_1551)
);

AO21x1_ASAP7_75t_L g1552 ( 
.A1(n_1516),
.A2(n_1496),
.B(n_1495),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1506),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1518),
.B(n_1470),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1507),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1518),
.B(n_1501),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1557)
);

NOR4xp25_ASAP7_75t_L g1558 ( 
.A(n_1526),
.B(n_1496),
.C(n_1488),
.D(n_1472),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1539),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1522),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1539),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1504),
.B(n_1494),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1565)
);

AOI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1512),
.A2(n_1490),
.B(n_1501),
.Y(n_1566)
);

NOR2x1_ASAP7_75t_L g1567 ( 
.A(n_1541),
.B(n_1479),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1537),
.Y(n_1568)
);

OR2x6_ASAP7_75t_L g1569 ( 
.A(n_1524),
.B(n_1342),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1504),
.B(n_1479),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1513),
.B(n_1494),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1513),
.B(n_1479),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1530),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1515),
.B(n_1481),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1515),
.B(n_1499),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1510),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1552),
.B(n_1537),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1577),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1508),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1547),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1567),
.A2(n_1549),
.B1(n_1537),
.B2(n_1569),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1569),
.A2(n_1534),
.B1(n_1533),
.B2(n_1525),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1548),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1574),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1551),
.B(n_1455),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1551),
.Y(n_1590)
);

INVxp33_ASAP7_75t_SL g1591 ( 
.A(n_1570),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1517),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1553),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1463),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1532),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1574),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1517),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1572),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1520),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1555),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1563),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1545),
.B(n_1532),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1593),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1593),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1590),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1582),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1582),
.A2(n_1556),
.B1(n_1557),
.B2(n_1566),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1600),
.Y(n_1609)
);

AOI32xp33_ASAP7_75t_L g1610 ( 
.A1(n_1589),
.A2(n_1552),
.A3(n_1550),
.B1(n_1559),
.B2(n_1560),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1585),
.A2(n_1568),
.B(n_1560),
.Y(n_1612)
);

AOI31xp33_ASAP7_75t_L g1613 ( 
.A1(n_1581),
.A2(n_1575),
.A3(n_1573),
.B(n_1548),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1591),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1600),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1592),
.B(n_1597),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1594),
.A2(n_1525),
.B1(n_1556),
.B2(n_1557),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1342),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1598),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_SL g1621 ( 
.A(n_1587),
.B(n_1559),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1624)
);

CKINVDCx16_ASAP7_75t_R g1625 ( 
.A(n_1606),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1619),
.B(n_1587),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1617),
.B(n_1599),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1599),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1620),
.B(n_1603),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1616),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1607),
.B(n_1602),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1554),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1616),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1625),
.B(n_1611),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1633),
.Y(n_1636)
);

AOI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1630),
.A2(n_1608),
.B(n_1612),
.C(n_1621),
.Y(n_1637)
);

OA22x2_ASAP7_75t_L g1638 ( 
.A1(n_1627),
.A2(n_1586),
.B1(n_1618),
.B2(n_1604),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1632),
.A2(n_1610),
.B(n_1613),
.Y(n_1639)
);

OAI31xp33_ASAP7_75t_L g1640 ( 
.A1(n_1631),
.A2(n_1596),
.A3(n_1622),
.B(n_1562),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1634),
.A2(n_1562),
.B1(n_1596),
.B2(n_1622),
.Y(n_1641)
);

AOI311xp33_ASAP7_75t_L g1642 ( 
.A1(n_1629),
.A2(n_1615),
.A3(n_1609),
.B(n_1605),
.C(n_1583),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1626),
.B(n_1627),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1636),
.B(n_1635),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1643),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1638),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1639),
.B(n_1624),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1637),
.A2(n_1623),
.B1(n_1565),
.B2(n_1592),
.Y(n_1648)
);

CKINVDCx16_ASAP7_75t_R g1649 ( 
.A(n_1645),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1646),
.A2(n_1641),
.B(n_1640),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1644),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1647),
.A2(n_1621),
.B1(n_1642),
.B2(n_1578),
.C(n_1601),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1648),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1649),
.A2(n_1628),
.B1(n_1578),
.B2(n_1601),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1651),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1654),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_R g1658 ( 
.A(n_1653),
.B(n_1652),
.Y(n_1658)
);

XNOR2xp5_ASAP7_75t_L g1659 ( 
.A(n_1650),
.B(n_1597),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1656),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1655),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1659),
.B(n_1564),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1660),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1657),
.B1(n_1661),
.B2(n_1662),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1658),
.B1(n_1542),
.B2(n_1530),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1665),
.A2(n_1525),
.B1(n_1542),
.B2(n_1508),
.Y(n_1666)
);

AOI22x1_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1571),
.B1(n_1564),
.B2(n_1540),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1667),
.Y(n_1668)
);

AOI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1667),
.A2(n_1542),
.B(n_1571),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1668),
.A2(n_1540),
.B1(n_1536),
.B2(n_1514),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1536),
.B(n_1519),
.Y(n_1671)
);

NOR2xp67_ASAP7_75t_L g1672 ( 
.A(n_1671),
.B(n_1509),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1670),
.A2(n_1509),
.B(n_1514),
.Y(n_1673)
);

AOI322xp5_ASAP7_75t_L g1674 ( 
.A1(n_1672),
.A2(n_1673),
.A3(n_1520),
.B1(n_1521),
.B2(n_1529),
.C1(n_1527),
.C2(n_1523),
.Y(n_1674)
);

AOI22x1_ASAP7_75t_L g1675 ( 
.A1(n_1672),
.A2(n_1493),
.B1(n_1481),
.B2(n_1528),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1523),
.B1(n_1519),
.B2(n_1528),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1676),
.A2(n_1674),
.B1(n_1521),
.B2(n_1529),
.Y(n_1677)
);


endmodule