module real_aes_7599_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_112;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_0), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_1), .A2(n_226), .B(n_230), .C(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_2), .A2(n_221), .B(n_317), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_3), .A2(n_49), .B1(n_111), .B2(n_116), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_4), .B(n_258), .Y(n_324) );
INVx1_ASAP7_75t_L g206 ( .A(n_5), .Y(n_206) );
AND2x6_ASAP7_75t_L g226 ( .A(n_5), .B(n_204), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_5), .B(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g187 ( .A1(n_6), .A2(n_188), .B1(n_191), .B2(n_192), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_6), .Y(n_191) );
INVx1_ASAP7_75t_L g237 ( .A(n_7), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_8), .B(n_235), .Y(n_272) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_9), .A2(n_29), .B1(n_96), .B2(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g219 ( .A(n_10), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g82 ( .A1(n_11), .A2(n_33), .B1(n_83), .B2(n_84), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_11), .A2(n_238), .B(n_252), .C(n_256), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_12), .B(n_258), .Y(n_257) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_13), .A2(n_32), .B1(n_96), .B2(n_100), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_14), .B(n_364), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_15), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_16), .A2(n_282), .B(n_283), .C(n_285), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_17), .B(n_235), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_18), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_19), .B(n_235), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_20), .Y(n_306) );
INVx1_ASAP7_75t_L g294 ( .A(n_21), .Y(n_294) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_22), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_23), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_24), .A2(n_48), .B1(n_123), .B2(n_127), .Y(n_122) );
INVx1_ASAP7_75t_L g360 ( .A(n_25), .Y(n_360) );
AOI22xp5_ASAP7_75t_SL g522 ( .A1(n_25), .A2(n_85), .B1(n_181), .B2(n_360), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_26), .A2(n_46), .B1(n_132), .B2(n_136), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_27), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_28), .A2(n_57), .B1(n_184), .B2(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_28), .Y(n_185) );
INVx2_ASAP7_75t_L g224 ( .A(n_30), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_31), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g197 ( .A1(n_32), .A2(n_43), .B1(n_55), .B2(n_198), .C(n_199), .Y(n_197) );
INVxp67_ASAP7_75t_L g200 ( .A(n_32), .Y(n_200) );
INVx1_ASAP7_75t_L g84 ( .A(n_33), .Y(n_84) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_33), .A2(n_282), .B(n_320), .C(n_322), .Y(n_319) );
INVxp67_ASAP7_75t_L g361 ( .A(n_34), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_35), .A2(n_230), .B(n_293), .C(n_299), .Y(n_292) );
CKINVDCx14_ASAP7_75t_R g318 ( .A(n_36), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_37), .A2(n_234), .B(n_236), .C(n_239), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_38), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_39), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_40), .Y(n_146) );
INVx1_ASAP7_75t_L g280 ( .A(n_41), .Y(n_280) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_42), .A2(n_65), .B1(n_189), .B2(n_190), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_42), .Y(n_190) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_43), .A2(n_68), .B1(n_96), .B2(n_100), .Y(n_103) );
INVxp67_ASAP7_75t_L g201 ( .A(n_43), .Y(n_201) );
CKINVDCx14_ASAP7_75t_R g228 ( .A(n_44), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_45), .A2(n_85), .B1(n_181), .B2(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_45), .Y(n_534) );
INVx1_ASAP7_75t_L g204 ( .A(n_47), .Y(n_204) );
INVx1_ASAP7_75t_L g218 ( .A(n_50), .Y(n_218) );
INVx1_ASAP7_75t_SL g321 ( .A(n_51), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_52), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_53), .B(n_258), .Y(n_287) );
INVx1_ASAP7_75t_L g309 ( .A(n_54), .Y(n_309) );
AO22x2_ASAP7_75t_L g105 ( .A1(n_55), .A2(n_73), .B1(n_96), .B2(n_97), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_56), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_57), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_58), .A2(n_221), .B(n_227), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g88 ( .A1(n_59), .A2(n_72), .B1(n_89), .B2(n_106), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_60), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_61), .A2(n_221), .B(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_62), .A2(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g250 ( .A(n_63), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_64), .Y(n_291) );
INVx1_ASAP7_75t_L g189 ( .A(n_65), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_66), .A2(n_221), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g253 ( .A(n_67), .Y(n_253) );
INVx2_ASAP7_75t_L g216 ( .A(n_69), .Y(n_216) );
INVx1_ASAP7_75t_L g269 ( .A(n_70), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_71), .A2(n_230), .B(n_308), .C(n_311), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_74), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_75), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g96 ( .A(n_76), .Y(n_96) );
INVx1_ASAP7_75t_L g98 ( .A(n_76), .Y(n_98) );
INVx2_ASAP7_75t_L g284 ( .A(n_77), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_194), .B1(n_207), .B2(n_520), .C(n_521), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_182), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_85), .B2(n_181), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_SL g181 ( .A(n_85), .Y(n_181) );
AND2x2_ASAP7_75t_SL g85 ( .A(n_86), .B(n_140), .Y(n_85) );
NOR2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_121), .Y(n_86) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_110), .Y(n_87) );
INVx2_ASAP7_75t_SL g89 ( .A(n_90), .Y(n_89) );
INVx11_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x6_ASAP7_75t_L g91 ( .A(n_92), .B(n_101), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
OR2x2_ASAP7_75t_L g144 ( .A(n_93), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_99), .Y(n_93) );
AND2x2_ASAP7_75t_L g109 ( .A(n_94), .B(n_99), .Y(n_109) );
AND2x2_ASAP7_75t_L g114 ( .A(n_94), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x2_ASAP7_75t_L g154 ( .A(n_95), .B(n_99), .Y(n_154) );
AND2x2_ASAP7_75t_L g161 ( .A(n_95), .B(n_103), .Y(n_161) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g100 ( .A(n_98), .Y(n_100) );
INVx2_ASAP7_75t_L g115 ( .A(n_99), .Y(n_115) );
INVx1_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
AND2x4_ASAP7_75t_L g108 ( .A(n_101), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g113 ( .A(n_101), .B(n_114), .Y(n_113) );
AND2x6_ASAP7_75t_L g153 ( .A(n_101), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
AND2x2_ASAP7_75t_L g126 ( .A(n_102), .B(n_105), .Y(n_126) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g119 ( .A(n_103), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_103), .B(n_105), .Y(n_130) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
INVx1_ASAP7_75t_L g160 ( .A(n_105), .Y(n_160) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx6_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g135 ( .A(n_109), .B(n_119), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g149 ( .A(n_109), .B(n_126), .Y(n_149) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g118 ( .A(n_114), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g125 ( .A(n_114), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g128 ( .A(n_114), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g159 ( .A(n_115), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g180 ( .A(n_120), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_131), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g145 ( .A(n_126), .Y(n_145) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x6_ASAP7_75t_L g138 ( .A(n_130), .B(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx8_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx4f_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx6_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
NOR3xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_150), .C(n_168), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_146), .B2(n_147), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI221xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B1(n_156), .B2(n_162), .C(n_163), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AND2x4_ASAP7_75t_L g166 ( .A(n_161), .B(n_167), .Y(n_166) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_161), .B(n_173), .Y(n_172) );
BUFx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B1(n_174), .B2(n_175), .Y(n_168) );
INVx3_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B1(n_187), .B2(n_193), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_183), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g192 ( .A(n_188), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
AND3x1_ASAP7_75t_SL g196 ( .A(n_197), .B(n_202), .C(n_205), .Y(n_196) );
INVxp67_ASAP7_75t_L g526 ( .A(n_197), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_SL g528 ( .A(n_202), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_202), .A2(n_230), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g538 ( .A(n_202), .Y(n_538) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_203), .B(n_206), .Y(n_531) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_SL g537 ( .A(n_205), .B(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_450), .Y(n_209) );
NAND5xp2_ASAP7_75t_L g210 ( .A(n_211), .B(n_365), .C(n_397), .D(n_414), .E(n_437), .Y(n_210) );
AOI221xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_288), .B1(n_325), .B2(n_329), .C(n_333), .Y(n_211) );
INVx1_ASAP7_75t_L g477 ( .A(n_212), .Y(n_477) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_260), .Y(n_212) );
AND3x2_ASAP7_75t_L g452 ( .A(n_213), .B(n_262), .C(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_245), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_214), .B(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g340 ( .A(n_214), .Y(n_340) );
AND2x2_ASAP7_75t_L g344 ( .A(n_214), .B(n_276), .Y(n_344) );
INVx2_ASAP7_75t_L g374 ( .A(n_214), .Y(n_374) );
OR2x2_ASAP7_75t_L g385 ( .A(n_214), .B(n_277), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_214), .B(n_261), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_214), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g464 ( .A(n_214), .B(n_277), .Y(n_464) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_220), .B(n_242), .Y(n_214) );
INVx1_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_215), .A2(n_266), .B(n_291), .C(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g314 ( .A(n_215), .Y(n_314) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g244 ( .A(n_216), .B(n_217), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
BUFx2_ASAP7_75t_L g355 ( .A(n_221), .Y(n_355) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_222), .B(n_226), .Y(n_266) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g231 ( .A(n_224), .Y(n_231) );
INVx1_ASAP7_75t_L g286 ( .A(n_224), .Y(n_286) );
INVx1_ASAP7_75t_L g232 ( .A(n_225), .Y(n_232) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_225), .Y(n_235) );
INVx3_ASAP7_75t_L g238 ( .A(n_225), .Y(n_238) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_225), .Y(n_255) );
INVx4_ASAP7_75t_SL g241 ( .A(n_226), .Y(n_241) );
BUFx3_ASAP7_75t_L g299 ( .A(n_226), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_SL g227 ( .A1(n_228), .A2(n_229), .B(n_233), .C(n_241), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_229), .A2(n_241), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_229), .A2(n_241), .B(n_280), .C(n_281), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_229), .A2(n_241), .B(n_318), .C(n_319), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_SL g356 ( .A1(n_229), .A2(n_241), .B(n_357), .C(n_358), .Y(n_356) );
INVx5_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g520 ( .A(n_230), .B(n_299), .Y(n_520) );
AND2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
BUFx3_ASAP7_75t_L g240 ( .A(n_231), .Y(n_240) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_231), .Y(n_323) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g282 ( .A(n_235), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx5_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
INVx2_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g256 ( .A(n_240), .Y(n_256) );
INVx1_ASAP7_75t_L g311 ( .A(n_241), .Y(n_311) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_243), .Y(n_247) );
INVx4_ASAP7_75t_L g259 ( .A(n_243), .Y(n_259) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g352 ( .A(n_244), .Y(n_352) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_245), .Y(n_343) );
AND2x2_ASAP7_75t_L g405 ( .A(n_245), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_245), .B(n_261), .Y(n_424) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g332 ( .A(n_246), .B(n_261), .Y(n_332) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_246), .Y(n_339) );
AND2x2_ASAP7_75t_L g391 ( .A(n_246), .B(n_277), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_246), .B(n_260), .C(n_374), .Y(n_416) );
AND2x2_ASAP7_75t_L g481 ( .A(n_246), .B(n_262), .Y(n_481) );
AND2x2_ASAP7_75t_L g515 ( .A(n_246), .B(n_261), .Y(n_515) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_257), .Y(n_246) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_247), .A2(n_278), .B(n_287), .Y(n_277) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_247), .A2(n_316), .B(n_324), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_254), .B(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_254), .A2(n_295), .B1(n_360), .B2(n_361), .Y(n_359) );
INVx4_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_259), .B(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_259), .B(n_301), .Y(n_300) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_259), .A2(n_305), .B(n_312), .Y(n_304) );
INVxp67_ASAP7_75t_L g341 ( .A(n_260), .Y(n_341) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_276), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_261), .B(n_374), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_261), .B(n_405), .Y(n_413) );
AND2x2_ASAP7_75t_L g463 ( .A(n_261), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g491 ( .A(n_261), .Y(n_491) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g398 ( .A(n_262), .B(n_391), .Y(n_398) );
BUFx3_ASAP7_75t_L g430 ( .A(n_262), .Y(n_430) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_274), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_267), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_266), .A2(n_306), .B(n_307), .Y(n_305) );
O2A1O1Ixp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_272), .C(n_273), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_273), .B(n_309), .C(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g406 ( .A(n_276), .Y(n_406) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_277), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_282), .B(n_321), .Y(n_320) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_288), .A2(n_466), .B1(n_468), .B2(n_469), .Y(n_465) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_302), .Y(n_288) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_326), .Y(n_325) );
INVx3_ASAP7_75t_SL g336 ( .A(n_289), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_289), .B(n_369), .Y(n_401) );
OR2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_303), .Y(n_420) );
AND2x2_ASAP7_75t_L g425 ( .A(n_289), .B(n_377), .Y(n_425) );
AND2x2_ASAP7_75t_L g428 ( .A(n_289), .B(n_370), .Y(n_428) );
AND2x2_ASAP7_75t_L g440 ( .A(n_289), .B(n_315), .Y(n_440) );
AND2x2_ASAP7_75t_L g456 ( .A(n_289), .B(n_304), .Y(n_456) );
AND2x4_ASAP7_75t_L g459 ( .A(n_289), .B(n_327), .Y(n_459) );
OR2x2_ASAP7_75t_L g476 ( .A(n_289), .B(n_412), .Y(n_476) );
OR2x2_ASAP7_75t_L g507 ( .A(n_289), .B(n_349), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_289), .B(n_435), .Y(n_509) );
OR2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_300), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_296), .C(n_297), .Y(n_293) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_298), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_302), .B(n_347), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_302), .B(n_370), .Y(n_502) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_315), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_303), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g369 ( .A(n_303), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g377 ( .A(n_303), .B(n_349), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_303), .B(n_327), .Y(n_395) );
OR2x2_ASAP7_75t_L g412 ( .A(n_303), .B(n_370), .Y(n_412) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
AND2x2_ASAP7_75t_L g435 ( .A(n_304), .B(n_315), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g364 ( .A(n_314), .Y(n_364) );
INVx2_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
INVx1_ASAP7_75t_L g447 ( .A(n_315), .Y(n_447) );
AND2x2_ASAP7_75t_L g497 ( .A(n_315), .B(n_336), .Y(n_497) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_326), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g381 ( .A(n_326), .B(n_336), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_326), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g368 ( .A(n_327), .B(n_336), .Y(n_368) );
OR2x2_ASAP7_75t_L g484 ( .A(n_328), .B(n_458), .Y(n_484) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_331), .B(n_464), .Y(n_470) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OAI32xp33_ASAP7_75t_L g426 ( .A1(n_332), .A2(n_427), .A3(n_429), .B1(n_431), .B2(n_432), .Y(n_426) );
OR2x2_ASAP7_75t_L g443 ( .A(n_332), .B(n_385), .Y(n_443) );
OAI21xp33_ASAP7_75t_SL g468 ( .A1(n_332), .A2(n_342), .B(n_373), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .B1(n_342), .B2(n_345), .Y(n_333) );
INVxp33_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_335), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_336), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g394 ( .A(n_336), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g494 ( .A(n_336), .B(n_435), .Y(n_494) );
OR2x2_ASAP7_75t_L g518 ( .A(n_336), .B(n_412), .Y(n_518) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_337), .A2(n_400), .B(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_339), .B(n_344), .Y(n_396) );
AND2x2_ASAP7_75t_L g418 ( .A(n_340), .B(n_391), .Y(n_418) );
INVx1_ASAP7_75t_L g431 ( .A(n_340), .Y(n_431) );
OR2x2_ASAP7_75t_L g436 ( .A(n_340), .B(n_370), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_343), .B(n_385), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_367), .B1(n_372), .B2(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_347), .A2(n_409), .B1(n_416), .B2(n_417), .Y(n_415) );
AND2x2_ASAP7_75t_L g493 ( .A(n_347), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_349), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g512 ( .A(n_349), .B(n_395), .Y(n_512) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B(n_362), .Y(n_349) );
INVx1_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_354), .A2(n_363), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_357), .Y(n_532) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_378), .B1(n_379), .B2(n_384), .C(n_386), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_368), .B(n_370), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_368), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_369), .A2(n_475), .B(n_476), .C(n_477), .Y(n_474) );
AND2x2_ASAP7_75t_L g479 ( .A(n_369), .B(n_459), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_369), .A2(n_458), .B(n_518), .C(n_519), .Y(n_517) );
BUFx3_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_373), .B(n_430), .Y(n_473) );
AOI211xp5_ASAP7_75t_L g492 ( .A1(n_373), .A2(n_493), .B(n_495), .C(n_501), .Y(n_492) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVxp67_ASAP7_75t_L g453 ( .A(n_375), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_377), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_381), .A2(n_398), .B(n_399), .C(n_407), .Y(n_397) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
OR2x2_ASAP7_75t_L g499 ( .A(n_385), .B(n_429), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_393), .B2(n_396), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_388), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g486 ( .A(n_390), .B(n_430), .Y(n_486) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g441 ( .A(n_391), .B(n_431), .Y(n_441) );
INVx1_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_395), .B(n_409), .Y(n_457) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_405), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g514 ( .A(n_406), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_413), .Y(n_407) );
INVx1_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_409), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_409), .B(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g460 ( .A(n_409), .B(n_435), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_409), .B(n_456), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_409), .A2(n_419), .B(n_459), .C(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_419), .B1(n_421), .B2(n_425), .C(n_426), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_423), .B(n_431), .Y(n_505) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_425), .A2(n_440), .B(n_442), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_428), .B(n_435), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_429), .B(n_482), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
INVxp33_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g445 ( .A1(n_434), .A2(n_446), .B(n_448), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_434), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_435), .B(n_489), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_444), .C(n_445), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_441), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g475 ( .A(n_447), .Y(n_475) );
NAND5xp2_ASAP7_75t_L g450 ( .A(n_451), .B(n_478), .C(n_492), .D(n_503), .E(n_516), .Y(n_450) );
AOI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B(n_461), .C(n_474), .Y(n_451) );
INVx2_ASAP7_75t_SL g498 ( .A(n_452), .Y(n_498) );
NAND4xp25_ASAP7_75t_SL g454 ( .A(n_455), .B(n_457), .C(n_458), .D(n_460), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g461 ( .A1(n_460), .A2(n_462), .B(n_465), .C(n_471), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_463), .A2(n_504), .B1(n_506), .B2(n_508), .C(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI221xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B1(n_483), .B2(n_485), .C(n_487), .Y(n_478) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_486), .A2(n_509), .B1(n_511), .B2(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_495) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI322xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .A3(n_527), .B1(n_529), .B2(n_532), .C1(n_533), .C2(n_535), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
endmodule