module fake_jpeg_4924_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_26),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_27),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_21),
.B1(n_16),
.B2(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_21),
.B1(n_11),
.B2(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_30),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_48),
.C(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_18),
.B1(n_11),
.B2(n_19),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_25),
.B(n_24),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_44),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_47),
.C(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_7),
.B1(n_3),
.B2(n_5),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_43),
.Y(n_60)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_61),
.C(n_62),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_38),
.B1(n_43),
.B2(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_54),
.B1(n_55),
.B2(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_25),
.C(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

HB1xp67_ASAP7_75t_SL g64 ( 
.A(n_57),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_67),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_50),
.C(n_51),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_54),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_49),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.C(n_73),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_17),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_68),
.B1(n_6),
.B2(n_8),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_8),
.B(n_9),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_74),
.Y(n_77)
);


endmodule