module fake_jpeg_15606_n_388 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_14),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_61),
.B(n_54),
.C(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_0),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_54),
.B(n_62),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_1),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_36),
.B1(n_15),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_29),
.B1(n_37),
.B2(n_24),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_36),
.B1(n_63),
.B2(n_15),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_75),
.A2(n_84),
.B(n_99),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_36),
.B1(n_15),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_76),
.A2(n_110),
.B1(n_111),
.B2(n_34),
.Y(n_151)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_15),
.B1(n_31),
.B2(n_27),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_45),
.B(n_28),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_2),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_49),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_26),
.B1(n_22),
.B2(n_39),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_24),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_117),
.Y(n_150)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_121),
.Y(n_147)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_124),
.Y(n_155)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_40),
.A2(n_39),
.B1(n_22),
.B2(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_26),
.B1(n_39),
.B2(n_22),
.Y(n_129)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_78),
.B1(n_105),
.B2(n_94),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_130),
.A2(n_158),
.B1(n_169),
.B2(n_149),
.Y(n_215)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_131),
.Y(n_178)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_23),
.B1(n_20),
.B2(n_55),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_134),
.A2(n_141),
.B1(n_162),
.B2(n_163),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_23),
.B1(n_59),
.B2(n_33),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_169),
.B(n_174),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_153),
.Y(n_177)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_166),
.Y(n_195)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_96),
.B1(n_12),
.B2(n_13),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_11),
.Y(n_192)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_107),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_167),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_34),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_171),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_82),
.A2(n_34),
.A3(n_33),
.B1(n_17),
.B2(n_8),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_11),
.A3(n_12),
.B1(n_79),
.B2(n_91),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_90),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_105),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_173),
.Y(n_199)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_99),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_9),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_93),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_170),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_10),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_88),
.B(n_33),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_95),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_75),
.A2(n_33),
.B1(n_34),
.B2(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_85),
.B(n_33),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_109),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_160),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_201),
.C(n_159),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_204),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_76),
.B(n_89),
.C(n_114),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_186),
.B(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_192),
.B1(n_151),
.B2(n_174),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_127),
.A2(n_11),
.B(n_12),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_83),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_202),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_147),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_215),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_205),
.B(n_172),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_91),
.C(n_100),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_100),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_137),
.B(n_11),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_120),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_120),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_209),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_145),
.B(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_217),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_159),
.B1(n_166),
.B2(n_170),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_211),
.A2(n_182),
.B1(n_200),
.B2(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_149),
.B(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_150),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_142),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_254),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_222),
.B1(n_235),
.B2(n_201),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_178),
.B1(n_190),
.B2(n_188),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_220),
.A2(n_176),
.B1(n_232),
.B2(n_253),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_252),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_143),
.B1(n_132),
.B2(n_157),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_155),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_199),
.C(n_216),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_143),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_135),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_236),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_253),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_132),
.B1(n_157),
.B2(n_135),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_133),
.B1(n_152),
.B2(n_138),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_251),
.B1(n_245),
.B2(n_221),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_131),
.A3(n_139),
.B1(n_138),
.B2(n_128),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_244),
.A3(n_230),
.B1(n_229),
.B2(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_250),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_185),
.B1(n_205),
.B2(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_193),
.B(n_172),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_182),
.B1(n_183),
.B2(n_205),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_176),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_256),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_233),
.B(n_235),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_265),
.C(n_276),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_273),
.B1(n_277),
.B2(n_248),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_178),
.B1(n_188),
.B2(n_214),
.Y(n_262)
);

OAI22x1_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_240),
.B1(n_232),
.B2(n_222),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_270),
.B1(n_279),
.B2(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_189),
.C(n_215),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_266),
.B(n_267),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_219),
.A2(n_195),
.B1(n_178),
.B2(n_217),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_195),
.B(n_209),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_272),
.A2(n_275),
.B(n_270),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_206),
.B1(n_179),
.B2(n_213),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_177),
.C(n_196),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_283),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_246),
.A2(n_181),
.B1(n_179),
.B2(n_177),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_280),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_252),
.B1(n_225),
.B2(n_226),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_287),
.A2(n_299),
.B1(n_305),
.B2(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_233),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_301),
.C(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_262),
.B1(n_264),
.B2(n_266),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_298),
.A2(n_279),
.B1(n_272),
.B2(n_262),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_243),
.B1(n_224),
.B2(n_227),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_224),
.Y(n_300)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_227),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_241),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_302),
.B(n_308),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_247),
.B(n_249),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_274),
.B(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_218),
.C(n_259),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_218),
.B1(n_275),
.B2(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_310),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_317),
.A2(n_319),
.B1(n_321),
.B2(n_323),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_271),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_325),
.C(n_330),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_264),
.B1(n_278),
.B2(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_284),
.B1(n_285),
.B2(n_269),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_285),
.C(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_293),
.B1(n_297),
.B2(n_307),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_327),
.A2(n_297),
.B1(n_298),
.B2(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_288),
.C(n_287),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_315),
.B1(n_324),
.B2(n_333),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_342),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_288),
.C(n_289),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_345),
.C(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_300),
.Y(n_341)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_341),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_291),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_331),
.B(n_324),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_346),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_304),
.B1(n_309),
.B2(n_311),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_313),
.B1(n_315),
.B2(n_342),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_299),
.C(n_310),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_312),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_325),
.C(n_318),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_319),
.B(n_327),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_357),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_335),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_360),
.C(n_338),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_317),
.B(n_322),
.Y(n_357)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_331),
.C(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_314),
.Y(n_360)
);

AOI21x1_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_321),
.B(n_347),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_344),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_355),
.A2(n_337),
.B1(n_346),
.B2(n_341),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_364),
.A2(n_356),
.B1(n_357),
.B2(n_362),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_363),
.B(n_339),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_365),
.B(n_370),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_355),
.B(n_348),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_354),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_375),
.B(n_360),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_364),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_352),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_377),
.B(n_378),
.Y(n_381)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_374),
.A2(n_367),
.B(n_368),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_371),
.C(n_372),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_380),
.B(n_358),
.Y(n_382)
);

NAND4xp25_ASAP7_75t_SL g383 ( 
.A(n_382),
.B(n_376),
.C(n_381),
.D(n_358),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_383),
.A2(n_373),
.B(n_369),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_384),
.A2(n_351),
.B(n_376),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_368),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_373),
.C(n_349),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_353),
.B1(n_313),
.B2(n_347),
.Y(n_388)
);


endmodule