module fake_jpeg_1442_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_0),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_0),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_53),
.B1(n_55),
.B2(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_43),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_1),
.Y(n_88)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_1),
.B(n_2),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_4),
.B(n_5),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_69),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_17),
.C(n_36),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_89),
.C(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_92),
.Y(n_106)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_2),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_97),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_27),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_84),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_89),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_87),
.B(n_25),
.C(n_26),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_23),
.B(n_29),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_8),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_40),
.B(n_31),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_22),
.C(n_32),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_112),
.C(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_122),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_116),
.B1(n_101),
.B2(n_113),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_12),
.B(n_14),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_110),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_118),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_132),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_129),
.C(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_142),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_138),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_126),
.B(n_137),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_127),
.B(n_123),
.Y(n_150)
);


endmodule