module real_aes_9979_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_0), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g15 ( .A(n_1), .B(n_8), .C(n_16), .Y(n_15) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_1), .B(n_7), .C(n_21), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_2), .B(n_5), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g21 ( .A(n_3), .B(n_17), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_4), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_6), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_9), .Y(n_23) );
NAND2xp33_ASAP7_75t_R g10 ( .A(n_11), .B(n_24), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
NAND2xp33_ASAP7_75t_R g12 ( .A(n_13), .B(n_23), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_14), .B(n_19), .Y(n_13) );
NAND2xp33_ASAP7_75t_R g14 ( .A(n_15), .B(n_18), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_22), .Y(n_19) );
endmodule