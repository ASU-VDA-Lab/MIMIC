module fake_aes_267_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
HB1xp67_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_7), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_14), .B(n_8), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx3_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_17), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_16), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_15), .B1(n_18), .B2(n_0), .C(n_6), .Y(n_24) );
AOI22x1_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_26) );
endmodule