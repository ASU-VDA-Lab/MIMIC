module fake_jpeg_8776_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_18),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_26),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_58),
.B1(n_59),
.B2(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_52),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_27),
.B1(n_29),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_16),
.B1(n_20),
.B2(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_74),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_72),
.B1(n_73),
.B2(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_66),
.Y(n_88)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_22),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_20),
.B(n_25),
.C(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_41),
.C(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_47),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_25),
.B(n_26),
.C(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_0),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_63),
.B(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_97),
.B1(n_50),
.B2(n_48),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_56),
.B1(n_43),
.B2(n_49),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_68),
.B1(n_62),
.B2(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_19),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_1),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_105),
.C(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_36),
.C(n_41),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_91),
.C(n_87),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_19),
.B1(n_15),
.B2(n_17),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_50),
.B1(n_17),
.B2(n_15),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_129),
.B1(n_130),
.B2(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_125),
.C(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_1),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_95),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_86),
.A3(n_96),
.B1(n_95),
.B2(n_94),
.C1(n_81),
.C2(n_93),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_101),
.C(n_107),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_84),
.B1(n_97),
.B2(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_94),
.B1(n_17),
.B2(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_99),
.B1(n_103),
.B2(n_109),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_128),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_108),
.B1(n_104),
.B2(n_105),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_133),
.A3(n_137),
.B1(n_121),
.B2(n_119),
.C1(n_140),
.C2(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.C(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_139),
.B(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_106),
.C(n_53),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_106),
.C(n_53),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_116),
.C(n_53),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_152),
.C(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_14),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_3),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_127),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_155),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_14),
.B(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_159),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_2),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_152),
.B1(n_143),
.B2(n_10),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_148),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_4),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_165),
.B1(n_154),
.B2(n_153),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_144),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_3),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_6),
.B(n_8),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_163),
.C(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_172),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_164),
.C(n_167),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_6),
.B(n_8),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);


endmodule