module fake_netlist_1_9688_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp33_ASAP7_75t_L g11 ( .A(n_2), .B(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_11), .B(n_0), .Y(n_17) );
OAI22xp5_ASAP7_75t_SL g18 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_19), .B(n_16), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
BUFx3_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI22xp33_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_22), .B1(n_12), .B2(n_15), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_22), .B(n_25), .Y(n_28) );
AOI211xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B(n_17), .C(n_21), .Y(n_29) );
AOI21xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_22), .B(n_23), .Y(n_30) );
NOR2xp33_ASAP7_75t_SL g31 ( .A(n_30), .B(n_22), .Y(n_31) );
OR5x1_ASAP7_75t_L g32 ( .A(n_29), .B(n_1), .C(n_3), .D(n_4), .E(n_5), .Y(n_32) );
NAND5xp2_ASAP7_75t_L g33 ( .A(n_28), .B(n_6), .C(n_7), .D(n_8), .E(n_9), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_21), .Y(n_34) );
XNOR2xp5_ASAP7_75t_L g35 ( .A(n_32), .B(n_7), .Y(n_35) );
NOR4xp75_ASAP7_75t_L g36 ( .A(n_34), .B(n_32), .C(n_33), .D(n_9), .Y(n_36) );
OAI221xp5_ASAP7_75t_R g37 ( .A1(n_36), .A2(n_14), .B1(n_23), .B2(n_35), .C(n_32), .Y(n_37) );
endmodule