module fake_jpeg_15465_n_271 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_271);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_13;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_7),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_19),
.B1(n_27),
.B2(n_15),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_27),
.B1(n_19),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_32),
.B1(n_31),
.B2(n_15),
.Y(n_64)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_28),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_69),
.B1(n_32),
.B2(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_32),
.B1(n_31),
.B2(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_28),
.Y(n_67)
);

NAND2xp67_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_52),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_42),
.C(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_72),
.B1(n_44),
.B2(n_91),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_42),
.C(n_32),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_28),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_91),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_100),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_72),
.B(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_76),
.B(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_73),
.B1(n_86),
.B2(n_77),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_109),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_55),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_64),
.B1(n_51),
.B2(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_63),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_34),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_58),
.B1(n_53),
.B2(n_57),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_19),
.B1(n_60),
.B2(n_27),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_108),
.B1(n_101),
.B2(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_114),
.B(n_110),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_93),
.B1(n_82),
.B2(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_134),
.B1(n_137),
.B2(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_63),
.C(n_29),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_133),
.C(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.Y(n_142)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_29),
.C(n_30),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_94),
.B1(n_107),
.B2(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_81),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_93),
.B1(n_82),
.B2(n_66),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_141),
.Y(n_178)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_98),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_160),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_97),
.C(n_112),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_129),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_110),
.C(n_99),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_128),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_114),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_124),
.B1(n_17),
.B2(n_22),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_121),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_117),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_82),
.B1(n_15),
.B2(n_89),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_37),
.B1(n_30),
.B2(n_17),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_144),
.B1(n_145),
.B2(n_158),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_124),
.Y(n_163)
);

XOR2x1_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_168),
.C(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_118),
.B1(n_132),
.B2(n_122),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_133),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_160),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_127),
.B1(n_17),
.B2(n_22),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_146),
.B1(n_36),
.B2(n_26),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_148),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_201),
.C(n_202),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_151),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_155),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_149),
.B1(n_141),
.B2(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_171),
.B1(n_163),
.B2(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_211),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_172),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_215),
.C(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_183),
.C(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_181),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_0),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_0),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_206),
.A2(n_203),
.B1(n_200),
.B2(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_229),
.B1(n_217),
.B2(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_201),
.C(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_198),
.C(n_37),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_207),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_37),
.C(n_29),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_214),
.C(n_212),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_24),
.B(n_21),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_218),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_235),
.Y(n_249)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_7),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_240),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_213),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.C(n_227),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.C(n_247),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_232),
.C(n_221),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_16),
.C(n_13),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_16),
.C(n_13),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_252),
.C(n_23),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_13),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_258),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_242),
.B(n_243),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_259),
.B(n_8),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_7),
.B(n_10),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_0),
.B(n_1),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_10),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_262),
.B(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_1),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_10),
.B(n_3),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_265),
.B(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_267),
.C(n_3),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_264),
.A2(n_253),
.B(n_16),
.Y(n_267)
);

AOI21x1_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_3),
.B(n_4),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_4),
.B(n_5),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_4),
.B(n_5),
.Y(n_271)
);


endmodule